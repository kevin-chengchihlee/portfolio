PK
     !M[������  ��     cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_0":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_1":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_2":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3":["pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1"],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_4":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_5":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_6":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_7":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_8":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_9":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_10":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_11":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_12":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_13":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14":["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_5"],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_15":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_16":["pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_7"],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_17":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_18":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_19":["pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_6"],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_20":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_21":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_22":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_23":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_24":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_25":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_26":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_27":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28":["pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0"],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_29":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_30":[],"pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0":["pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1"],"pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1":["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14"],"pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_4":["pin-type-component_b00b0f46-5dcc-4451-a676-221697210905_0"],"pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_5":["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14"],"pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_6":["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_19"],"pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_7":["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_16"],"pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0":["pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0"],"pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0":["pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0"],"pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1":["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3"],"pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0":["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28"],"pin-type-component_b00b0f46-5dcc-4451-a676-221697210905_0":["pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_4"]},"pin_to_color":{"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_0":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_1":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_2":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_4":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_5":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_6":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_7":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_8":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_9":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_10":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_11":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_12":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_13":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14":"#ff0000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_15":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_16":"#44ff00","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_17":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_18":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_19":"#0040ff","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_20":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_21":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_22":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_23":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_24":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_25":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_26":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_27":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_29":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_30":"#000000","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0":"#000000","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1":"#ff0000","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_4":"#000000","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_5":"#ff0000","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_6":"#0040ff","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_7":"#44ff00","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0":"#000000","pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0":"#000000","pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1":"#000000","pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0":"#000000","pin-type-component_b00b0f46-5dcc-4451-a676-221697210905_0":"#000000"},"pin_to_state":{"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_0":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_1":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_2":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_4":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_5":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_6":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_7":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_8":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_9":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_10":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_11":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_12":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_13":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_15":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_16":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_17":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_18":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_19":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_20":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_21":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_22":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_23":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_24":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_25":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_26":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_27":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_29":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_30":"neutral","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0":"neutral","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1":"neutral","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_4":"neutral","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_5":"neutral","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_6":"neutral","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_7":"neutral","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0":"neutral","pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0":"neutral","pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1":"neutral","pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0":"neutral","pin-type-component_b00b0f46-5dcc-4451-a676-221697210905_0":"neutral"},"next_color_idx":27,"wires_placed_in_order":[["pin-type-component_a3ae65d4-c858-4cbe-bb67-1538767c17f8_5","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_7"],["pin-type-component_a3ae65d4-c858-4cbe-bb67-1538767c17f8_7","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_8"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_29_polarity-pos"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_13","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_28_polarity-neg"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_29","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_29_polarity-pos"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_28_polarity-neg"],["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_1","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"],["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_0","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16"],["pin-type-fake_0","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16"],["pin-type-fake_1","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"],["pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_17","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16"],["pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_12","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"],["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_0","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_1"],["pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_0","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_1"],["pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_0","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_1"],["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_1"],["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_1","pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_1"],["pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_1","pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_1"],["pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_1","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1"],["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0"],["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_1"],["pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_1","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_1"],["pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_1","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_1"],["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_1","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_1"],["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0"],["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0","pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0"],["pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0","pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0"],["pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0"],["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_7","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_0"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_8","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_0"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_9","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_0"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_10","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_0"],["pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0"],["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3"],["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0","pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0"],["pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28"],["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0"],["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_5"],["pin-type-component_b00b0f46-5dcc-4451-a676-221697210905_0","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_4"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_19","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_6"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_16","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_7"],["pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0","pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0"],["pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3"]],"wires_removed_and_placed_in_order":[[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_a3ae65d4-c858-4cbe-bb67-1538767c17f8_5","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_7"]]],[[],[["pin-type-component_a3ae65d4-c858-4cbe-bb67-1538767c17f8_7","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_8"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[["pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_7","pin-type-component_a3ae65d4-c858-4cbe-bb67-1538767c17f8_5"]],[]],[[["pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_8","pin-type-component_a3ae65d4-c858-4cbe-bb67-1538767c17f8_7"]],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_29_polarity-pos"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_13","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_28_polarity-neg"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_29","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_29_polarity-pos"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_28_polarity-neg"]]],[[],[["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_1","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"]]],[[],[["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_0","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16"]]],[[["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_0","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16"]],[]],[[],[["pin-type-fake_0","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16"]]],[[],[]],[[["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_1","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"]],[]],[[],[["pin-type-fake_1","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"]]],[[],[]],[[["pin-type-fake_0","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16"]],[]],[[],[["pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_17","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16"]]],[[],[]],[[["pin-type-fake_1","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"]],[]],[[],[["pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_12","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"]]],[[],[]],[[["pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_12","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"]],[]],[[["pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_17"]],[]],[[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_13","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_28_polarity-neg"]],[]],[[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_28_polarity-neg"]],[]],[[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_29_polarity-pos"]],[]],[[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_29","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_29_polarity-pos"]],[]],[[],[["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_0","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_1"]]],[[],[["pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_0","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_1"]]],[[],[["pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_0","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_1"]]],[[],[["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_1"]]],[[],[["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_1","pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_1"]]],[[],[["pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_1","pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_1"]]],[[],[["pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_1","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1"]]],[[],[["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0"]]],[[["pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_1","pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_0"]],[]],[[["pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_1","pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_1"]],[]],[[["pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_0","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_1"]],[]],[[["pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_1","pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_1"]],[]],[[["pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_0","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_1"]],[]],[[["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1","pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_1"]],[]],[[["pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_1","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0"]],[]],[[["pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1"]],[]],[[],[["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_1"]]],[[],[["pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_1","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_1"]]],[[],[["pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_1","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_1"]]],[[],[["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_1","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_1"]]],[[],[["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0"]]],[[["pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0","pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0"]],[]],[[],[["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0","pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0"]]],[[],[["pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0","pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0"]]],[[],[["pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0"]]],[[],[["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_7","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_0"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_8","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_0"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_9","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_0"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_10","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_0"]]],[[],[["pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0"]]],[[],[["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3"]]],[[],[["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0","pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0"]]],[[],[["pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28"]]],[[],[["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0"]]],[[["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3"]],[]],[[["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1"]],[]],[[],[["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_5"]]],[[],[["pin-type-component_b00b0f46-5dcc-4451-a676-221697210905_0","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_4"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_19","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_6"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_16","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_7"]]],[[["pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_10"]],[]],[[["pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_1","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1"]],[]],[[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_9","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_0"]],[]],[[["pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_1","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_1"]],[]],[[["pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_8"]],[]],[[["pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_1","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_1"]],[]],[[["pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_7"]],[]],[[["pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_1","pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_1"]],[]],[[["pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0"],["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0","pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0"]],[["pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0","pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0"]]],[[["pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0","pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0"]],[]],[[["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0","pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0"]],[]],[[["pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0","pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0"]],[]],[[["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3"]],[]],[[],[["pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_0":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_1":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_2":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3":"0000000000000009","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_4":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_5":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_6":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_7":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_8":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_9":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_10":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_11":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_12":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_13":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14":"0000000000000010","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_15":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_16":"0000000000000014","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_17":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_18":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_19":"0000000000000013","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_20":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_21":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_22":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_23":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_24":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_25":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_26":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_27":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28":"0000000000000011","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_29":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_30":"_","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0":"0000000000000009","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1":"0000000000000010","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_4":"0000000000000012","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_5":"0000000000000010","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_6":"0000000000000013","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_7":"0000000000000014","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0":"0000000000000004","pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0":"0000000000000004","pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1":"0000000000000009","pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0":"0000000000000011","pin-type-component_b00b0f46-5dcc-4451-a676-221697210905_0":"0000000000000012"},"component_id_to_pins":{"f0fd6315-2925-41b3-9764-248681cdce0c":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30"],"636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35":["0","1"],"0232f75e-f080-4dd3-8137-8958c98da454":["4","5","6","7"],"2829c8e4-4312-47ed-a029-8eab57667ef2":["0"],"28debeb4-25ba-40b7-880d-a84ab194857a":["0","1"],"a21c1a89-038d-4d33-9463-f2151579a9e0":["0"],"e87dc4da-e2d8-41cc-bc12-69ed72c01d9e":[],"d710e40b-242b-4d55-aff1-d25d4416cf71":[],"b00b0f46-5dcc-4451-a676-221697210905":["0"],"2dd2b242-eb34-4791-b8ff-53525115782a":[],"208137c0-256c-4563-a200-a8fe7094349e":[],"b1be3c37-6458-4463-9c21-0cddf8035423":[]},"uid_to_net":{"_":[],"0000000000000004":["pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0","pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0"],"0000000000000009":["pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3"],"0000000000000011":["pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28"],"0000000000000010":["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_5"],"0000000000000012":["pin-type-component_b00b0f46-5dcc-4451-a676-221697210905_0","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_4"],"0000000000000013":["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_19","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_6"],"0000000000000014":["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_16","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_7"]},"uid_to_text_label":{"0000000000000004":"Net 4","0000000000000009":"Net 9","0000000000000011":"Net 11","0000000000000010":"Net 10","0000000000000012":"Net 12","0000000000000013":"Net 13","0000000000000014":"Net 14"},"all_breadboard_info_list":["bf214f1e-c792-43f5-846b-d34128e4e83a_30_2_True_955_100_up","bc941250-d2ab-4f36-99ca-60371a583e71_63_2_True_835_10_up","295e808d-80c9-46a1-9a2f-f0256ea548ee_30_2_True_940.5_145.49999999999955_right"],"breadboard_info_list":[],"componentsData":[{"compProperties":{},"position":[803.2100499999999,309.8848895],"typeId":"5dd9522a-ac85-4cae-b2c3-8ba3fec8b601","componentVersion":2,"instanceId":"f0fd6315-2925-41b3-9764-248681cdce0c","orientation":"left","circleData":[[752.5,230],[751.6624749999999,240.99967700000002],[752.7453145,250.29215899999986],[752.1075655,261.7580989999999],[752.3877774999999,271.7645255],[752.5665445,281.7735544999998],[752.5665445,291.86251249999987],[752.1075655,301.8715924999999],[753.0255249999998,311.49889699999983],[753.5859504999999,321.96691999999985],[752.5665445,332.78988649999985],[751.9287969999998,342.6227749999998],[752.8467579999997,353.5204279999999],[753.4845054999998,362.90210149999996],[753.4845054999998,373.2634804999999],[854.4709314999998,230.39584999999988],[854.4709314999998,240.90942199999995],[855.060628,251.10101299999997],[854.5456779999997,261.6919805],[855.135376,272.437451],[854.7284064999999,281.4854839999998],[854.3214354999998,292.41885049999996],[854.063962,302.0928889999999],[854.7284064999999,312.6888079999999],[854.8819884999998,322.9092259999999],[853.6610784999998,333.63743599999987],[854.4445854999999,343.0979329999999],[854.8819884999998,353.7271684999997],[854.0680494999999,364.2397129999998],[854.851555,374.5201729999998],[804.8739519999999,408.6976309999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"161","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"Adafruit Industries","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[625.654174,295.80002],"typeId":"84ae97c1-8e69-5e6b-4fa6-dfe46d477633","componentVersion":1,"instanceId":"636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35","orientation":"up","circleData":[[602.5,305],[648.8083479999996,305]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[453.1307005000001,383.442893],"typeId":"98d6e125-552a-4063-90e5-58c04872effd","componentVersion":1,"instanceId":"2829c8e4-4312-47ed-a029-8eab57667ef2","orientation":"up","circleData":[[452.5,365]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[654.5702454999994,1.0316959999999824],"typeId":"db03155d-4b7a-4e64-a4d7-f9e505c5d345","componentVersion":3,"instanceId":"0232f75e-f080-4dd3-8137-8958c98da454","orientation":"up","circleData":[[902.5,94.99999999999999],[902.7937105000001,113.74855700000005],[902.2139035,132.35993000000008],[902.0429485,150.4458965]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"10000","displayFormat":"input","showOnComp":true,"isVisibleToUser":true,"name":"Resistance","unit":"Ω","required":true,"validRange":[0,70000]},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.25%","value":"0.25%"},{"label":"0.1%","value":"0.1%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false,"isVisibleToUser":true,"name":"Tolerance","required":true},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"string","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false,"isVisibleToUser":true,"name":"Number Of Bands","required":true}},"position":[502.22504875383447,305.69373781154127],"typeId":"72c75556-baa3-04e7-55a5-e13f447c8c5a","componentVersion":1,"instanceId":"28debeb4-25ba-40b7-880d-a84ab194857a","orientation":"up","circleData":[[467.5,305],[542.5,305]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1008.1307005000001,383.4428929999999],"typeId":"98d6e125-552a-4063-90e5-58c04872effd","componentVersion":1,"instanceId":"a21c1a89-038d-4d33-9463-f2151579a9e0","orientation":"up","circleData":[[1007.5000000000001,365]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"5v dc","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[688.5146147612892,322.037732766394],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"e87dc4da-e2d8-41cc-bc12-69ed72c01d9e","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"5v dc","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[891.2520860259777,419.8110375396785],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"d710e40b-242b-4d55-aff1-d25d4416cf71","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1008.1307004999999,83.44289299999994],"typeId":"98d6e125-552a-4063-90e5-58c04872effd","componentVersion":1,"instanceId":"b00b0f46-5dcc-4451-a676-221697210905","orientation":"up","circleData":[[1007.5,65.00000000000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"GPIO21 SDA","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[910.120468903076,258.0396692910173],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"2dd2b242-eb34-4791-b8ff-53525115782a","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"GPIO22 SCL","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[909.54183626089,221.79194479635257],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"208137c0-256c-4563-a200-a8fe7094349e","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"GPIO34","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[693.7762858314251,242.75732919044282],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"b1be3c37-6458-4463-9c21-0cddf8035423","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"-247.74580","left":"304.15575","width":"731.79691","height":"696.05684","x":"304.15575","y":"-247.74580"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0\",\"endPinId\":\"pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0\",\"rawStartPinId\":\"pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0\",\"rawEndPinId\":\"pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"452.5000000000_365.0000000000\\\",\\\"452.5000000000_305.0000000000\\\",\\\"467.5000000000_305.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1\",\"endPinId\":\"pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0\",\"rawStartPinId\":\"pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1\",\"rawEndPinId\":\"pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"542.5000000000_305.0000000000\\\",\\\"602.5000000000_305.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1\",\"endPinId\":\"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3\",\"rawStartPinId\":\"pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1\",\"rawEndPinId\":\"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"542.5000000000_305.0000000000\\\",\\\"542.5000000000_261.7580990000\\\",\\\"752.1075655000_261.7580990000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0\",\"endPinId\":\"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28\",\"rawStartPinId\":\"pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0\",\"rawEndPinId\":\"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1007.5000000000_365.0000000000\\\",\\\"870.7840247500_365.0000000000\\\",\\\"870.7840247500_364.2397130000\\\",\\\"854.0680495000_364.2397130000\\\"]}\"}","{\"color\":\"#ff0000\",\"startPinId\":\"pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1\",\"endPinId\":\"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14\",\"rawStartPinId\":\"pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1\",\"rawEndPinId\":\"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"648.8083480000_305.0000000000\\\",\\\"730.0000000000_305.0000000000\\\",\\\"730.0000000000_372.5000000000\\\",\\\"753.4845055000_372.5000000000\\\",\\\"753.4845055000_373.2634805000\\\"]}\"}","{\"color\":\"#ff0000\",\"startPinId\":\"pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_5\",\"endPinId\":\"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14\",\"rawStartPinId\":\"pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_5\",\"rawEndPinId\":\"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"902.7937105000_113.7485570000\\\",\\\"1067.5000000000_113.7485570000\\\",\\\"1067.5000000000_440.0000000000\\\",\\\"767.5000000000_440.0000000000\\\",\\\"767.5000000000_373.2634805000\\\",\\\"753.4845055000_373.2634805000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_4\",\"endPinId\":\"pin-type-component_b00b0f46-5dcc-4451-a676-221697210905_0\",\"rawStartPinId\":\"pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_4\",\"rawEndPinId\":\"pin-type-component_b00b0f46-5dcc-4451-a676-221697210905_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"902.5000000000_95.0000000000\\\",\\\"902.5000000000_65.0000000000\\\",\\\"1007.5000000000_65.0000000000\\\"]}\"}","{\"color\":\"#0040ff\",\"startPinId\":\"pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_6\",\"endPinId\":\"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_19\",\"rawStartPinId\":\"pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_6\",\"rawEndPinId\":\"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_19\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"902.2139035000_132.3599300000\\\",\\\"977.5000000000_132.3599300000\\\",\\\"977.5000000000_272.4374510000\\\",\\\"855.1353760000_272.4374510000\\\"]}\"}","{\"color\":\"#44ff00\",\"startPinId\":\"pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_7\",\"endPinId\":\"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_16\",\"rawStartPinId\":\"pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_7\",\"rawEndPinId\":\"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_16\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"902.0429485000_150.4458965000\\\",\\\"955.0000000000_150.4458965000\\\",\\\"955.0000000000_240.9094220000\\\",\\\"854.4709315000_240.9094220000\\\"]}\"}"],"projectDescription":""}PK
     !M[               jsons/PK
     !M[�qE�>  �>     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"ESP32 (30 pin)","category":["User Defined"],"userDefined":true,"id":"5dd9522a-ac85-4cae-b2c3-8ba3fec8b601","subtypeDescription":"","subtypePic":"f51f6ed9-d8f0-454d-af8a-e11415a94f15.png","iconPic":"53dea2ad-2eb7-451c-84a6-1b4fef66a2aa.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"13.80107","numDisplayRows":"7.59928","pins":[{"uniquePinIdString":"0","positionMil":"1222.61943,718.03100","isAnchorPin":true,"label":"EN"},{"uniquePinIdString":"1","positionMil":"1149.28825,723.61450","isAnchorPin":false,"label":"VP"},{"uniquePinIdString":"2","positionMil":"1087.33837,716.39557","isAnchorPin":false,"label":"VN"},{"uniquePinIdString":"3","positionMil":"1010.89877,720.64723","isAnchorPin":false,"label":"D34"},{"uniquePinIdString":"4","positionMil":"944.18926,718.77915","isAnchorPin":false,"label":"D35"},{"uniquePinIdString":"5","positionMil":"877.46240,717.58737","isAnchorPin":false,"label":"D32"},{"uniquePinIdString":"6","positionMil":"810.20268,717.58737","isAnchorPin":false,"label":"D33"},{"uniquePinIdString":"7","positionMil":"743.47548,720.64723","isAnchorPin":false,"label":"D25"},{"uniquePinIdString":"8","positionMil":"679.29345,714.52750","isAnchorPin":false,"label":"D26"},{"uniquePinIdString":"9","positionMil":"609.50663,710.79133","isAnchorPin":false,"label":"D27"},{"uniquePinIdString":"10","positionMil":"537.35352,717.58737","isAnchorPin":false,"label":"D14"},{"uniquePinIdString":"11","positionMil":"471.80093,721.83902","isAnchorPin":false,"label":"D12"},{"uniquePinIdString":"12","positionMil":"399.14991,715.71928","isAnchorPin":false,"label":"D13"},{"uniquePinIdString":"13","positionMil":"336.60542,711.46763","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"14","positionMil":"267.52956,711.46763","isAnchorPin":false,"label":"Vin"},{"uniquePinIdString":"15","positionMil":"1219.98043,38.22479","isAnchorPin":false,"label":"D23"},{"uniquePinIdString":"16","positionMil":"1149.88995,38.22479","isAnchorPin":false,"label":"D22"},{"uniquePinIdString":"17","positionMil":"1081.94601,34.29348","isAnchorPin":false,"label":"TX0"},{"uniquePinIdString":"18","positionMil":"1011.33956,37.72648","isAnchorPin":false,"label":"RX0"},{"uniquePinIdString":"19","positionMil":"939.70309,33.79516","isAnchorPin":false,"label":"D21"},{"uniquePinIdString":"20","positionMil":"879.38287,36.50829","isAnchorPin":false,"label":"D19"},{"uniquePinIdString":"21","positionMil":"806.49376,39.22143","isAnchorPin":false,"label":"D18"},{"uniquePinIdString":"22","positionMil":"742.00017,40.93792","isAnchorPin":false,"label":"D5"},{"uniquePinIdString":"23","positionMil":"671.36071,36.50829","isAnchorPin":false,"label":"TX2"},{"uniquePinIdString":"24","positionMil":"603.22459,35.48441","isAnchorPin":false,"label":"RX2"},{"uniquePinIdString":"25","positionMil":"531.70319,43.62381","isAnchorPin":false,"label":"D4"},{"uniquePinIdString":"26","positionMil":"468.63321,38.40043","isAnchorPin":false,"label":"D2"},{"uniquePinIdString":"27","positionMil":"397.77164,35.48441","isAnchorPin":false,"label":"D15"},{"uniquePinIdString":"28","positionMil":"327.68801,40.91067","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"29","positionMil":"259.15161,35.68730","isAnchorPin":false,"label":"3V3"},{"uniquePinIdString":"30","positionMil":"31.30189,368.87132","isAnchorPin":false,"label":"USB POWER"}],"pinType":"wired"},"properties":[],"componentVersion":2,"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Photocell (LDR)","category":["Input"],"id":"84ae97c1-8e69-5e6b-4fa6-dfe46d477633","subtypeDescription":"","subtypePic":"b63deb06-c33f-4ae3-8f73-25229955b1c1.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.58334,76.55539","endPositionMil":"14.58334,14.58330","isAnchorPin":true,"label":"pin 0"},{"uniquePinIdString":"1","startPositionMil":"323.30566,76.55539","endPositionMil":"323.30566,14.58330","isAnchorPin":false,"label":"pin 1"}],"numDisplayCols":"3.37889","numDisplayRows":"1.51833","pinType":"movable"},"userDefined":false,"properties":[{"type":"string","name":"mpn","value":"161","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Adafruit Industries","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"a5640015-ff5c-4848-bb8b-6d4b42e5489b.png","componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"GND","category":["User Defined"],"id":"98d6e125-552a-4063-90e5-58c04872effd","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1cdb40d8-22d5-4761-8204-85ee5f97d036.png","iconPic":"9ee875d8-7c7b-435c-a3d9-92ac29f03ab9.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"2.37626","numDisplayRows":"3.61380","pins":[{"uniquePinIdString":"0","positionMil":"114.60833,303.64262","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"LCD 16x2 attached i2c","category":["User Defined"],"id":"db03155d-4b7a-4e64-a4d7-f9e505c5d345","componentVersion":3,"userDefined":true,"subtypeDescription":"","subtypePic":"99708c53-ae63-4787-a3c4-6dca09af2b7b.png","iconPic":"62b25533-4940-4036-93a8-d94b028d26e9.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"45.38860","numDisplayRows":"31.83700","pins":[{"uniquePinIdString":"4","positionMil":"3922.29503,965.39464","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"5","positionMil":"3924.25310,840.40426","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"6","positionMil":"3920.38772,716.32844","isAnchorPin":false,"label":"SDA"},{"uniquePinIdString":"7","positionMil":"3919.24802,595.75533","isAnchorPin":false,"label":"SCL"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Resistor","category":["Basic"],"id":"72c75556-baa3-04e7-55a5-e13f447c8c5a","subtypeDescription":"","subtypePic":"bbfae99c-8036-4c5e-89fd-a87441410720.png","userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[{"type":"double","name":"Resistance","value":200,"unit":"Ω","showOnComp":true,"required":true,"validRange":[0,70000]},{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}],"iconPic":"a262aa33-74c4-460b-b0ad-c746896f6744.png","componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"GND","category":["User Defined"],"id":"98d6e125-552a-4063-90e5-58c04872effd","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1cdb40d8-22d5-4761-8204-85ee5f97d036.png","iconPic":"9ee875d8-7c7b-435c-a3d9-92ac29f03ab9.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"2.37626","numDisplayRows":"3.61380","pins":[{"uniquePinIdString":"0","positionMil":"114.60833,303.64262","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"GND","category":["User Defined"],"id":"98d6e125-552a-4063-90e5-58c04872effd","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1cdb40d8-22d5-4761-8204-85ee5f97d036.png","iconPic":"9ee875d8-7c7b-435c-a3d9-92ac29f03ab9.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"2.37626","numDisplayRows":"3.61380","pins":[{"uniquePinIdString":"0","positionMil":"114.60833,303.64262","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""}]}PK
     !M[               images/PK
     !M[ZR�y�Z �Z /   images/f51f6ed9-d8f0-454d-af8a-e11415a94f15.png�PNG

   IHDR  �  '   js1   	pHYs  P�  P���Dm   tEXtSoftware www.inkscape.org��<  ��IDATx���U��Ϧ��酄H� AJDz��D�P�@T���J�RB	%�^ ����Fz��o��ܝ̼u�}gv��y&��}wf�̝;�ι��ټy�(��(��(��(�R^�H©���m�lg��f��l��Vo���lx*DQEQEQEQ����l̶�l+�����6��͛7ϗ��8�n9��`�fke��[��EQEQEQE)��f[h��r�u��>3��f{����<�Dtsa�0_.0[_�u2[{Q�<�ٳ�t��1��̞=[f͚˾[�n-�{��:u�},/^,ӦM�6D�����K߾}�Y�f'�W���ӧ����#߷���ԡC���?�\���X���@;�f��޽شiS��nԨ��L4m�T�d�ʕ^������M�ӧ��m�V���>�/��2�}w��Y�w�.q��W_Ɍ3$��wM�4���*N�c׬Y��k׮��E��<s�Ϗ'�ԭ[7�ڵ���ܹs��O?�e�-Z���'�{q�t�R�?�[�.�}׭[��O-[��8Y�~�7�b�A�=�S�N7qڀmڴ�^�z�n.Z�Ȼq؀)���:n�`w�k�9��=�|}�l7��Q<7=e��=̗�e���%[�䊒7����V�Z�ntA�.]�^�z��2J0���Eq�k׮�aÆ�|�4����~�g)�mòe�"�'bj���Ҹq㒴����������{�=q�3����GE*ҹ��c�Ҹ����;�,���'֣��?x�`π/Eb,�U��gDF	�!�37�v�A>��HE:�{��������.2v�Xϙ�s�5�U�m�Y��?^�͛�q� �4h q�c��L�4)���8�i����#�v�g������w�СCe�ƍ��'Λ���F.�q0 nK1�22�O�:5��b��޽�i'qـ����nh�c̘����f��G�3:��DI1�a���l;�Fʕ"� ��Q�E�J�[q�aG2D/�hw�-��R`���D��D��̇����D:��S
qn�}8*�n�9�oQ� ��)*�n�y�v�"u"e;���G%�1H��~��r�a�J�[q�����}�cF%ҭ8��d�)��A�y��J���DPő]}��V��*U�w����Ü;��(U�ƉZ�ӗ�S����n;�kT"ݵ� j���~�~=ӌ����W���8Z2�n���r��v�-���(�8/Q�tw`.5QЮ8/5Q�tW����Dz9Ĺ%*���R�Hw�y9�J�[q^��8/5Q�tW���(E��� *���R�Hw�y��R�[q^�����Ap�zm��7c������caL�dt�l�<�E��r�sK�"���������R�H/�8�+��)�-Ŋ�r�sK�"����R�H/�8�+��)�-Ŋ�r�sK"����R�H/�8�+��)�-Q��r�sK�"�:؀5�n[�������z�S"Mϊm�1'̾j�S��C%"� �-���$̖B�$�sK�"=)��R�HO�8�*ғ �-��t�g�C�Ź�P��qn)T�'A�[
�I�bDzĹ�P��qn)T�'A�[��I�BEzu���9��#�5c��Q�8��Ɯ�`��f�AD�ֺ��$�-���$̖|�$�sK�"=i�ܒ�HO�8��+ғ$�-�����sK�"=I�ܒ�H��?�.	�ܒ�HO�8�"ғ$�-���$�s����\�t$I�[
�I�|Ezu��*p#���3Fo���m��6��~l���l]DQ"$�����%� �āْ� �Dqn�U�'U�[r�I�\E:���RE���HO�8��*ғ(�-���$�sK�"=��ܒ�HO�8��*ғ(�-��m�$ғ(�-���=�M�'��U�WP	���F��]3N�jƕw��Yd#�9���Ͷ���]�V�q$y`�d��<0[��I�l"=��܂H�p�9sf��,�-�Dz�Ź%�H�yf�y)�9/�l"=��ܒM�'Y�[���$�sK."=��ܒM�'Y�[���$�s���D�ڀ�AEz$M��'�0�ʯ
�I$��9�6��3fۙoEQ"$�%l�N��l	�� �-a"=-��b\�HO�8����4�sK�HO�8����4�sK�HO�8����4�s��<���ϯ�4�sK�HO�8����4�sK&��6`iQ�	,��8��|%��w�ܢGs���˿�6X%b�40[�t�f��N�8��Ez�Ĺ�/��$�-~��&qn����s�_��I�[�"=M����i��b��\)��$�-~��&qn��4�sK�HW�<�H�����֌��3c˚|������5ͩX�W%b�80[� �hѢ��h�����{mH�8�X�N�.]��N�[���!�6qn�F
F�$M��bE:��gϞ��+�#i�+�q\џ�$�-V�ӟxߥI�[\���-m��bE�ܹs�q*M��bE:��D�Ĺ�錯j����� ��׌���wn���<��3_5[oQ��I�8�0@ӆ4�)K���e��vK��ł��ђ�� ��4��>bĈT�'D����%������o"��|in"=����w���Hǉ��{�H�u�]=��V8w�aE�ǧ�`�@"}Æ��^f{��r]/� �n������\�	��N;�/ɐfc�R�ThJ��>T�3���3Q]��"���R��Sb P��'��k���4ۓ[#��}8o�nvL���6PEQEQEQE	�+�=([�g$/�n�9;��ن��(��(��(��(�@wf����7o�2�����*���T�#�����ߺ����(��(��(�R,��/5����G+�u)��|��r��l����鯅}(g�nvt�l	�דҀ�c�/�6�lo��}�-1!X<��ٚ�qNT7��4��:���(��(��(��(���\�})[����e�f[a�U�E�#�ъ����l;���lY���l)�Vj:��OF[�4"}I�r�f�%C�����q.�Gf����f�H��m�ƛ��s�̑?_�܌^���(��(��(��(�Q>M�+���Y>����̧f{����Dt�(��b6V&#�[ʪ~�w�R��2����Z�x9&�'�ùT�ˆ����s�5_.�-Q���JBi\S��o6۪�ɮ�Z��&���׷z]�lڜ�ʡ�?���z3�ې�{�����?��4q��$�A�A�MR;�)�^W��'I,uko�zu2�����?%���eN�a���D�S�z�M[2ߋU�?mNt�d�S�Ϭ]_!6%�?�L�lgb�c�nHvjd��lE��ޟ꛱�N��'��������m��iG��6��uje�I���s��i�ˌƛ]���>��S��A�[��W��l��R�����g�s���Y��ÃdKi�8`Q�O�v�9��tn����˦-��כ�6T��<(5�����3h���^�����J�6�2~���[ɬE����?�;��.���Of7�'6���Ȉ�l�i�y���Z�����D:�X��3��Z�-K´�`v�JF�Y��3�|�Dޚ�D�J�F䔑3~f��:���6�d��P�7��_��me���.�{�e�v_g�̫��ʇ�7��ҡ�:9f�⌟�bq=���V�dN��$����v�~crE�>��ˀN�3~��OZ��$��h�V�4�g�}�@���Y�9؀�~����d�Tz�ͼ������k sV���Eq`k��eF'^m��\�L��.�������J2
t�Xe�6[�8�HI��9�R�q�5m�S�D�d�>�(��(��(��$�Q�;��q�8�9޴+�Vd�5����"M��6����0[�Z���Dp�r�O1�)1��vs��و�W+W��(��(��(J
a��Cf��ȶMRb�1)<��/2_/�-�����c����P�n>H��{��Rl���َ1'�Jʈ9�\�ƽ��d�cE�iSEQEQE)3���8�>�9�[�V|I�s㡘[q�l��I|��hÑ6���N.�7$�����6�����EQEQEQ�����	LI��`��c��7��a0,�C5��o�7�o�� )�Dϣ���rh���%	Ĝ�զ�Lο�l-EQEQEQE)��v��dS$a��U�St|��C���v8߄E�)��?��~�lgK�1�&s�8�-��~EQEQEQ���vbŹŜ�R�1�}�l��t�]�1��c}&Џ��枿c��gK4�/5��li�\DPQEQEQ%���%IJkck�����1�v1���.3�ۈps`����@����R-�'˖��vEQEQEQ%jȲ��щ���`�u���t#=��#��+��䗚�MXn����̖a�w��.ߗ-ޑN�(��(��(��D�f�����d��A濣b�}/���"�Q�e]�(x�4��B�y�3��y�g���+��(��(��Dk��8eY�.>g.zTY疦f��?�>�l�#������ӏ��
(%�O�k��3��ż�Y�0gc��,XU��x�bq���b��d�a����mذ)�E0��M�A���i�ڒd�ϯo�1�^�u]I2+���ڟ�mL�}�W�4�:�2���j]����_6��K3�?�Wԓ$�xUݬ�i������'4�Z��mL�8���������e���-���?�X���Tl���5�If��Ăɶ�^6�|��s��+**�f��s��n�e{�O�h���0'>KR�9�U��?*[.|�� JV(Q8����v�,I�a��V�6[����Mբ?}�(��i��u�-ͬ�P�Z��Oԗ��`E]oK3��U��i���v��=oY����5f|Z���Tml���go�@�%�~��~��E��NA�b��lWH��" ǚm�(��(��(��(��4�9�rL�WTT�C���(�HZU
ts v�-��~���ek���D��(��(��(J1,6۵R}�I�� �+ʝ�t��\��֚�n�^�,[�Eo+��(��(��(J!Lۼy�x�&��|]QQ1Ib軛�q��c��'�a.�tsᧉ
tEQEQEQ�ByQ�w�m�EV8��;G��OS\.?xzvEQEQEQ%_Ho��T?^0�l�p�5W���`�K��!��d�F���e˖I�V�D)?�7o�F�����%9hR%����D�ڵke͚5Q��K�?�J5ôi�y�b�Ū�%f��TO�2�<���$|��G2dȐT��E�ɒ%K�w�Ȟג�n�:�2e�0@��I�RVS�N��;J�fQ�"Y���+Y�z�t��]�
/�3fx��V�t�^��;q�D�>4n\쬰�1g���\���+WʬY�d��O� ٸq�ןxO4l��e����vQ�z���y��I߾}S۟6l� �&M�~��I�z�]���D˖-�,3؀���'�#����x�;���w���R�͐j�V�i*�KFK�E:3�i�&Ϡ�ӧ���c���_�	áC��R�c�̞=[���K6lX*E:���O>���Q�#��O�%^�<�i�\��?�X�ϟ/.��w�9�"q�s��S�N�6������{�v�!u�ʾ�/^,K�.��SE�̙3eڴi��<xp*E:���>�.�'b���Nhˊ+���F�N_�Oծ][m�2�ڀ2W�/c�vvT;s��b��Ŭ'՗Ţ����tw`^4���?0[�%M"�F:��'�64o�\҂_�c�@�D�+��>#i�8���M�[qn���I���xF M"��`����t+��>#i�8�H�Hw�9���)M"݊sP�|�$��]���o��R|��ó�� ��[��}-���2QJN�h��lI� 60�I��Ź�1i�~qnI�H��sK�D�_�[�BfF�&M$���9�g� ���ܒ&��疴�tW�[�&���ܒ&��疴�tW�[�,=1�s�j��Z �K���T�F�!�	
	���/��e��-i���i�a�ܒ�&�-i�a�ܒ�&�-v�^�Ez�8��E���sKDz�8��E��sKZDz�8��A���sKZDz�8��X:b�@��R}Yi��V2�6VE��uR�Y"J�H� �m`�$y��u`N�H�&�-I��Ĺ%�"=�8�$Y��<s�Ĺ%�"=�8�$]�g�$��l�ܒt��I�[�.ҳ�sK�Ez6qnI�H�$�-j�O���;�l��3�m4cDdZ�Z׈�dYF�c�(e%�t��%����I鹊sKREz��ܒD���8�$Q��*�-I鹈sKREz��ܒD���8�$U��"�-I鹊sKE����|yn�K�*�s����TG�A��u}�޴��$m��w`�$i���#80rlѵ�u�M�)�|Ź%i"=_qnI�H�W�[�$��疤��|Ĺ%i"=_qnI�H�W�[�&��疤��|Ź%I"=_qnI�H�G�[����s@'���f\�p����R���B�����Ѕ̖$Ѕ�s���酊sKRDz��܂������C�E��ܒ�^�8�$E�"�-�̈́	�kѥK),ŵ�W�[� �疤��BĹ%)"���>��üŹ%	"�PqnI�H/D�[����sh [j�UWx�G�����?�Kuo_�(� ]��la��x�۷���bŹ��"�Xqn)�H/V�[�O��}-�HG�ӟ
�r��bŹ��"�q�b�J/�H/V�[�)ҋ�r��bĹ��"�Xqn)�H/V�[�-ҋ��dB9Dz��9` 2ۛR=�&: ��-�`U���^�\�
� ]ʗLT�e֬Y��R���Ĺ��"*qnqEz)��Ĺ�"=*qnqEz��yF@,X� ���"��D%�-V��o�^JET����R�8��"��D!�-�Ho�,���r"*qnqEz��J�[\�^J���b�#PSqn���)���"<�
t��2�d�f�x��м(K��E����l�"�gϞ7\�(ŹŊ�Ry���+����_r���)K)E�5��k���[��
��ĹŊt�S)23x�L�y�c^�n�$n֮]�/*qn�"�c,�?Jqn�"�_�~R
�������ܹ��d��ɑ�s��c�fQ�s���Q�s��cKaR� N���kV&q�?��c�(w�@��TC�.[.zQ	��%y	��XQ��ٳg������łA�"��d��"0�J՟�6]�QCA��L җ,Y����H'C�^��8��ƌ7q�'D:N�4���t�S)��՟�����S�J��ٟ����KuB��7.�c,�e|e������T_"��F�>�f�Q�Ǜ��(��3N�T��+%e�#�������O�a����@����)hJ�***���mjN�1mb�E�·�z/s�u̅O�SR��M\SEQEQE�^0]�4�])Ջ�$����:��7�?��PQQ����$HEQEQEQ���>R�8W"^�;j��"��K5�K�V�򵊢(��(��(Տ>7o�<A��-�ȗt�Z�Î�d��������ӣ(��(��(�RJZ��Z�%Ճ�Ȗ�H�C�w2�uf;Y��4�(��(��(��ToFTTTtڼys�k喘��pm��Q�;�{1w�\�Y�R��,P�=�(��(��(�R�b�ߙ�8I7L��ǎ�蔚��lߑ�r��0�@)��-[V����3-MQ�~}i��U�֯_/+W��_����n�U������|�e�y4�A�I۶m�I�&�l�2o]�iӦyk'Ѹqc�W�^��,-�t��m>W�Niڴi����N-�}��^��[c7j׮-͚5��k�ʪU��X�7o^emV�O��`:u�$ݺu�֭[{�6�|�h��Ki�wa��biذ�w�-�\c�ܵkW�-�Λ6��1}7��u�z}ȥ����y����~��Kн��O�t�����;v���:�\�+V~�?Vd��׃����\�p�l�۷��3m��㏫<����k��������t�\ؘ��;w�l�kG��o��.���&���Σ��޸ҪU+��>|���}���ܻwo���-��{���FPxo���`����l��3>��r.}�]�v�s�}�8w�!�r���^�.���h�O;8ۆL�=���g�g�%�͑	�u�>}�M�6ҢE��6̜93ﱎw<�z�Ĺ�������l1�E�9���~�ok;�����4ƀ���俶.Ŏ�A�������N�XA�s�Y���)�}͹�46Λ�B̹S��T�Օ�K�î��6�1I/0_F���(��^�aÆU~��ʣ�>��[o�U�9�������_.;����?�Cqq���E]${��6/~���o�C=$��ߪ���{�}��U>?r�Hy뭷��l�=���^z���|PN:������^3��ŋ=��wޑ�����A�;� ~�a��0���������ߗ���a<X?�p�e�]���q�Q���/�.]�������^n��@Êk���;o�s^´cƌ������-�<�L�����)��"Ç�ڀQ��?��O���ۃ:H�<�L�k��<�����k��v�z�}�����������%�0}��w����"�#Fȡ�Zy0�-8\�I60�C�[��v�a��?�\_�6,Z��k��s������o/�\r���>ңG�m~�@z�'��.���y�'��rK����;��sϭ������-�m7n�������ac}�6�p����c�y�X�u �5�\#�w�6�4ƕ��{��0�,g�q������
3��'����C��o?������+��\ǣ��>E����/����޳��:49mx�7�699���2dH�X��|���e���^��C�>�`���|�=ό+~��.��w���^{Mx��Pa�������W4Yx�}�Y��'O��;����o߾��g<��O~�9����h�+��i��/����~肃�G�Ƒ �����SOy��駟n������������V�?��m>kE�_|��{��9�	Ldܧ������'���\
�w/ϯ�/ǎ�م��Ƙd���ַ����ĉ+��~2�Ў�~X9����g���w�yn���v��gK�d���X��s�=�#��D�6���wq��iv�]�`g昹�;���d���������sj��ߠ1���5�ﶊ�4.�����k�q
�f��\��̅�#)��/���%�����%�
�O<1Tl"�F/�r�x���,'�pB��q�o���gD�����_������ֳgOO0c$�����'j���;���g�ctc�1�� c.0~��9 n��O����6^h׳�:K�L��	� ��q�|�Zy䑡��\z饞���k�q�ֽ{wO_}��r�m�y�`��c'C���?�F��m}c��I���]��~z�p�a|��
2���>W�z��#�8B~��_zۯ��m>{�G�~�q��'{�`��wt���N���;�,f�m.Qj�&6��*cN����w�d� �\���8��LaΊ(!rd�@$g'�aw��o�y"r<�a ��<��������9:�e��vZq�kώ9����=c�/��6��1�I�q�y��K�(׉��t��~h��Q����<����|���8�x�/��ϙ�'!�*��#m�s����j����1���!�oa�<�^�<�a�h���]�4*Ιg�f�162ކ���?.��h5}�W������	,�����`��O��\�;��p`��T8��2޳R�{���g�}&	��6��/)���3%�"�q
t���C�!���wa�@��f�Q�Ă���5,(R���B �B$�F:RO?�t��2���A�7�����
"
�+�t<�� c<���x�����a�!�0f0�â%@t�֟��	D�����d ���ц(� <��B��'zH���R:"�A��L ��(� @ `<c(Y�A�\�/)�>�|dJ�%uԦ���>�'0P���*�O"v��$�q̘1�F��ם҂��5��%�HW<���vAS0�dӐ5����[8���~�
�_"��8g?D[�Z�w��L�\@q��Apo����y�>����]%�C���B�B9�#��l�� ���`���A��YHM��+<��q@�q�0���]��++^��g���	�O���g���Gy}��ǽ'���x�0L��%�J��c��1�kXLb8��8���]���6p�8W�c�MAM9���=OF��7߼�ﹿ\�	&xm@#"�,��d�������aQ�����1H�d\�o��w8U\这�F�~���+��ɤ��n�(Γh��c�.��`��`���n�?��(xR������,��:!�C�2}�y�|<))��+sί�-��؈[��æA�l.��S"�92��������$�:D�"�~�ɍR`���M�`�ϭv�p��FH�҅���=��8��E����GX�'�A�4�\��h��ს@�.`�3il�"����a�z�����HÓ��,��{��h#|1`Ĺ!CA�y�Q-W�#��	t����|A^�xɭQ�0!�a�z�1��#F0����ta?s<�D���o2p<��<���ԩSe�]w��	D��я~T%���F�a�����F�~���  �=�_�����Iڀ ���]s�;��;,<��#�H��'������
|� cA�v�"�"#&�1d-px����\ѧ,��u�~r>D�0��Gn���F��~�����	J�&}>��W�����'���N���ӟ�T�3
������qA���l����w��M�(�hO=�T��C�mp� �h�;E�-Qd7����3��?�A���0��Z��A�f��c�s��D�x��$���d���Sѽއ�8��e��2\x��Y���Ls҉�s����6p�.[8��xQ}2O��\���f���� ��Tp��pt�^gludpp�Yp,����ta�FT2���p��@��;�"�[�A�{�>���� ��wQ�R�>����Ac:�?ׁ�s�/��3��c�)��̢���æ�$���^	����g��9�o�'	Ɯ#�J�n���U
��1� xs�+	�\��/�����x��@��_�c,��+"#�B:��yn�5^����@�cW�`Pqp"?T��ƙ?E��'���\���4�I�}��1m�C �Z^֤��ii�9gؼS^�v?�U�0�a��6Н�Y�g=�D�������N��F�sCT0��=B�q_]G
�.(�4���x�W���`����������5pj`p�)�nVI� 6@*=}=_���,�I�5����E��4�����}C���K�0�VB ��rAY;.d'�6 �������0�}{<�w�qG`�_���s��{�c��i�S-� �v�6� ��u�1݀��4W�uPF��W�g�����ﶁ��60�ȝ��p���br8a���g�1���OX}���Vl�9��8u�7��&7�s�q�:�Sa���p��de!������p�$��lpl"b�dX��~�v�
t�+���<�m�
���E��� ������l��v��yo������>q]���ڎM�s��A���� %ڊo�	���%(��&c��;׹օ���3n�>L�$�0iҤ*���:��?<�8.݂��Q	t�^(��2M�K<<s�m��I ��ЇL;H	(�@,�M�ȓ<#i�ts^�'��6��^�Ƕ���xح�@��,�F6�:;QL�%v"ሇ0C�ȟ[�2�%|.[D��M���0+�ʯ"c��m=��� m J��`�p�
+E	�z7 !J�C!`�ᤱ��)B�xCZ&����x���}<�6E�HN�B����h>:aΨ|�O��OZ��M����\G�\�9p��`�u! ����8�SG�&ڹ������y���%c�ی��\C2f���\11I(*f��D������mC����a����y����Ϙ^h�Y����`���]�F>�@(�EJX�� 8������8�x���6�f�D�3��﯇�oC>��V���:�]�� ��g�t���S����0��ę���;���IP(<�Dѹ���l��y�����%����!��_ԯXx��r�q�sW�3f����	����)8�p��f��mp�k������p<<{�M��a,rz�5��@`�[d��s�pH ��{nk��� �9��a�j�Q*���۠�i�q����O������8��梤'v�����)�=_���B!��Q���}�R���M�anA;��Os+���1��v#��,Dj0V��|"��t�~Q��/@<G��y���#՞��V@ �0��-��	R�]ㅨ0F}�E�n�p�f�At���kr?��8�lj;"1�!Ftg���A�́��A�ב�e�c@
�����
Ak������7,���H�';ß��0�q��/J!�^K$ڝ�B�@�D��'��h�1�2'G_�ř�B��&h�_�c�S|�~�� '���!b���`!��Z��@|Z��U	��dB�����/�q�b�x�y0������|�u�|}�n���q�afZ���@���Υ���;�)Mٞ!5w�; �y?U�g�BHLq�ʢ����#d� �xo�|���3��V��9cz��y���,�$��:���Ȝ�$�'�/���
�1mˮbkn�Y��w�_�s]�#q�N{�z�;���q�+DY����L
�a�� ��;��i
�E)����a����~�W�9^>��,�qK)��9��n�e��u���%¯�a����j:��-X��.6u�Ц/c�˃dZ�ſdVPZ)��]�͂��G\0&|1C0��~!�)�z?��`Z����lQ�lU��P�K�c$�vS%�Ґn_(�����,�8��¨���l!m�Xq�hD�3br��*�@�mpz.��;����}�x@�<��&��_�(Wh�+�s�d�c�dPA�\��=�0�}�� ��
��6 �b�当)ڌ�MC��a^y��]��
��6 �ڀh!��5��{XH�.�0��X�>Am`:GP8oR�q���D�=�hv� `y�g�K�1��=�ԭ�`�!A=���d`������Ԥ�&�i�|�bo�f�6}x^2M,��a�9j1��� z{.m��3���d
�[$���f�aW	"�H=�6R��2!�N����������晎���9V��{J�)�@�r<5Ϛ��c����޷��'��(���+����xi)n��֍m��
��{��ޟ�i��Ej=�.OA�����9�b�W��b������BR1�_���j���c�s�U׏�e8���p��R���CD�^[�U�P+�|�χ+)|ǔ����]0n�,�:Da��ې��&��l��Dt�_�-��>��1����;���6d��{�n
��%h�@"@D	�Z�s�X�8?�|���+*P�݆ �[���e�o1&�)��\�'�ȷ/�p_����6�ˬ���F�}����"ҋ��6p.�@����~'8�qv3%gs{���w����p*�aUL_b\�ɀ���u��������]�Q�@'��f.�,ȵ�Rw���'����Q�*� �u����$����r�� ��r�%��]����5r�[�fK�	�CH�aƨ���3IJ�9&�ǈ!�W��rt�^�ԇ�q���������?R�q�gW>J��Eb�����^��4D�\��?w3Ӳh�舛*k�K$�TJ7�3HO��nۈ�E�8*��B�+��+�5Cy�����0���C-(�0���q�C��5$�~3���L��Q�?�D��%D�,5��Ka��ZA�����u�u�s;��Bq�(ȵ\S�����!h�s�.�/�?��8'옅Q_��ߗ��@�g�[�aJ=������0}�V1���Bz.m��G���j�����6s�i���₸�/�LE�ɀ��$8I�/$��y��$����D߈�r�d��t{�Do���y���u2s�����|A��������kF�@��c��q���.A����f~.�V7�M_*D��Dx��%�kۀXdUo���)*�1�1Kf�-2KA�\W)dU�Z\O;Wޭo�3�����qg����ডG�f��C�sg*�I��2�A�+8ly����S!]�K����ɸ�ɜ�bq.x�Y����P��h�2�s���-S�K5w)�@�,"4�(��Y�Ѩ�̾yk��Hu��'�(e�yL���$�ϩ�N�Kݮ�[(~�Q�`ϥʺ�� �!��D�~�2�%A�Iq�/�U(r���B�^~��%���V`ǰ�خ��(+T���;@�9��\U�c�s��gL�v�s<�}��Rr?��S9p2����&��F��=�O�� ��%��8�ܔUo�i����_�h���=��צj�$1�����0�1�H�\C���s}�@t��o?F���&�A�&������N6WH�B��G�
�L�N�"l��ՊU"�̑���w�;�@�Za�5b�h!SW�~�Rgjc�ʹ*��=�=�\��4ԩp�8�8v�Xܚ.��AE�f��i�V�������g�n?.�/�wS�駙
s�j�`��G�Y��+�AZ��d)�������y˼��h�xAT��.`�����ªdYa��g��<g�6�]��mSl1F4�jpD����7su"��;G�]�GP�`R��e��s�y.H_��y6�I�l�Ў7���5/��*�@�paXC��+ͅb���f��P�n��;��+,$HсX�W�i<���
���߹D='ےk���yZ��/Q=^xQE1�H���(�F�q�z����6��� pp` ��K#��6A$�%�B7��ؐ;��( �����
X��]ـ�[K!
���͝��U����I�=`(��$ǧ�;Ǜ�V�l�~�0�֝�B�|�s?�8\\�#Ͽ\cF2B�BĊ��L�Y��Ž�A?�_eZ+"���b5��B�П]g�
gS&e�I~��=�u�ZBt�� %����r1�I}F����B�!Ӻ�SI����#r�����
tڇ����*�Ԅ(�4�YE���ϵ���A���q�w.��/�l��8[Z͏��5g��;�x��U���󖃦��v�耰v�c�<�.�F_#rn����P�mpS�� q�L}ȵ�9��|��&�Y,	G��[�2����M�f=;�W��<��Gg�����.��1w7[nk���t�3;lݎ0�s��č ����í47d��T�=��	���-��1�ƻ���4�@w Ƙ.��uT0/	ϥ[��Q%�k`��y��ai��� �׍�QD͙S�/\��5SJ��k����a�Sۅ��G����d+�Zr)�FT��" 1��º/z��B��
1I8"&�Q�Ӆyd�g~�)�� ���V;&�Žu�_[�*.r��=u�ĸ� Ÿ���m�\Qww*"2�:d��m`,�Dʡ��ՙ]�M� ���j���H���E��"�n�$��Uٮ��l�L˭!h?���&ϔu�X.��*K<r�����z8�������������t#�@AN��S��ܶ�Tb撒*�fv�L1����	��%��m�N9 ��h5s������<�l�q�P��#p�q'��=Ν�)W�r�qb��ׂ���w��``� c�-�J��SX���6�2��6���I�v�3�uw�Ǒ�_W�kaӿ-D�]a�S�w"Bş�Øλ�%[_b,�8��d�uk?p��Tkq������9_�Y�p���;��vW!�J�=�Q��d\�>�=iߟ�����7Q�T����ϥ��$N~��T#:oݘ>ڌex�����q���P]ʲ���t�&[���
t��E�󳺒@�&�]�m��ߖ-���$6�N�D��Fw�Ź�TBT����`�8���S�z�鶤��a8�"$�/��r�`�g[�7"��"G�}�0�B����o� K�E��)�\'k�Ͷ�>~�y08�	�X�0�g3AԖ�߈b��kh�#�n��1sS�Q��p�84s��� �2ER�f�'A�1��j��s�9�Q3�-����a`�R��½ɶf2s�����蟓I��?���.�:3�����/]��>��\�\��p�K@ҷ]q��v�p� ��Y��5� D�o��6O��}fs2�T���c��n&���X�g�X�>�9#��H�f��&�3�Qבɳ���f����NĴ�,E4���K���_C���;��$ך�C�1.q�{�n�A�my:�5[����w�D<������0�Y��?��:�pd�W(AT�=����T)�������`<�G5�zN�.�Zh�qo��Cf����	@�	��g' ό���Y���?�Ʌ}��B@�P ��甍6� ���	�@�d�VCX4�l�^���q�p�����[�����:G�5�٠�<v���³�i��쟊�Sp(���Txtٺ�������������NݭFejV�J�@���z��
�h���!�e��@�5"y.
a�G�|�\��<Q�B�2A��h �Ǌዱ�y��͔�
Š���=F'[��B-v�;�8�� �/�Lm�0v���1Q(d�	�O+�p~����.�� N�*��a�`8�B��|ٜS���#��z�-;DOÌ��~��(&mq�#��
���P�I�<83�I��9F<e��AaϠ��a˰��@ց���"��BR�-��l06�A�d�3���n*%\C�T&3���`N}�*��d�-w8ɩ�P�j/L- C��U��,�0pN���P�0H��p�aU(�(8�ê�G	�� ����Z4iЧ)��<� B<�5|�@����\B2�6�x�п� rS�]ш'��]P�l~on���$�CЦ�R�ȟꊈ$J@�H��X�<��
Zփ��n������ങv��@<`l`h`|�E�����h/B�"}T�'ښ)m�c�+ט%�AT��Q�&�`��B���s>�?6׌��ϋ���h���˵��9��̈́�~���-��z�YC�O+"
�R�����G�����o��&[���j:����|�AP� �ɽ�8�r�A����\+�+ڀ��V�/�g!�D�x�pJ2�����D��"H��@��Г�M�>,�9�6�}��r">�C��3QH[��q4W9�؜'�m ����05(ly$�'�=���s�����`��do�X B��E�>@�OP��C�Οc��#S �F����n�:�7�ݶ��#�O�l��9�̄�/dj��k�5D,�\K��G�F�]��D�7D�y�2�?.���yK�w�,�3�g���>\xF�9c	�������8�(�ǳ��*���&W'mw�-׊�B�xg�3��9���U��Eݟ����$��f�;��es�𿳊-К��wx&�~�N�j�����ff%iY8e[T�+�����F��+^L����+�$���s	�F/*0gZF����e���1��^A`�G��@d���zDw�w�9Y)��
��6&�^"`n��|�XOT��te�(!�8�(ڀ�Xl��~!�3ǔ�XHGg+����L�F�s����@�<l��3�6�<saɜ;�ڙ�i�=D��6���dl�=�h�!Sԛ�<l���Cδ$cR��L}�bI?{h���P���$�p drrg��t[A��v�f�W�?����ӆLEq������~[�q�m�?�X��I'C�6П�����@�?�q?�4�\����9�s�	���\pW�(
���s8�������R&�~9ɵZ������(߀!�z���]��\إɂ֝�F�h��I��R(vy�B�@Đi��_�	������lT�+��(��(��(JP��(��(��(��(	@��(��(��(��$ 芢(��(��(�� T�+��(��(��(J�D������0�4i"�����˗��s�����(��(��(�R��D���p��^���[:� �ΰl���?��g5j$��(��(��(��)(�R�5k&u��-z?���|k�ޕ�?��x���1��߮k+�ݯ���θW֮ݐ�8}{��__����7m�,Ǟz��5�_\u�б��}O��G���=\��j[�=�]a�ع�\v���/Y�Jμ�����q�,�Z.?�䑌s�'H�֍+����/ɛo��X��iڤ~��������Q��ף,�?aD����~%W���Y�s����qG��~��9��	�|ݺ��{N���o~v�O��Og.���2XN9��s�4e�����	�|������.u�Ԫ���~��L�<7c[��#=��ϲ����Y�~o����$g����߀��_��T��ϯ�~�M�&�/_�gg���x���ӥs��ƣ�����U�ׅ��� Çu���ɧ>��~G����ˎ�:W~��?ߗǞ� ���$�^yH����o��O�'�qvީ�\qɁ��/_�FN;���s�GI�.-+���ݯˋ�L�z�?��8i߮i�����W�����~~�}��yg|����g/��F�3�q9p��~�n��O��@F_�9��!�����r��O���_���
tEQE)�����K��Y�ڣO��_�Zo�p�����ШaC�o�@�֭�n�wݺ������!���ߛ�S�����]*��8�+y��i��:d�*�6����ӥs�*��⒫�%�7;��?Wh>��ͱ�d=��]{J��d�=��D?����>�W�skԨ~Nm�գ]���ء��x�K����������u�2g�п�]�*��٣���7ᙂ��6����W�gm�43�Y,��y��s��L�Ϟ����ʯ��t����P��j׮-w��v��w��ܚ4ih��̎�͛l�w�{��)����A��v��~��y9�i�A]̱�q�}1g����	�ߡk�s[�f}N�i߮E����iѢ��^�>�ox��5mP����M��X#v�^eLyc�g����Y���ҳʹ����8�>ޯO{#���<���T��ۮmss�E�(��@��8��%ڶm+��$�^��_=��S��}��ҵkW)7'N���zJ%i�9�ے��ٳ�G��7F��Z�j���.��zj$b�֮]+��s���G?�M�6�������J��9s��~����k�I�پ�̿����0��+L�-�ܱE4���>�yd�}�ԯ_Gzl�J>�lT��ٶ�8/���w���h�b�Q�z��(�]��ͥy��l��؎�����'g�}���֌��""~��:}Hd�s���	�G��}�Nͫ��b�v���8�Z�l$�����8�D$!x�G�����z=�/_.����c9�;��3��~�3����EQ��~��'W_}�$��}��5�\�~G�%�s�$�w�<��s���Gn���D�s�޽���/�>}�H��ޭ��6���yw�6��]��s�N�넣��˯M��1G�L��[/Oh��bۈ+�����8ᘝ�W�y.�wG��8�;���7� +Vn+j{vo-#vέ�n6xG�,<26���G�&�3���������Y������eÆM��n���<'J Ȉ�>�ҶE~��9T��~E�z�$�Ջ�8;�,������~6�+�;lG���*У��?@Z�j,�o;��c�f��ь�8k�:�ǿ�N<&�6)�Mq��%;��%I�|��*�%G��k�X�۫W/I���vn={���R��I�kGɨc��MD�'?�WzE����q��Cv�=�I��#�.�ᾑx�u�ˉg�'��}�I����k�,g���<��$y��w�CN9~xd�!���"�~�JJ}�u����9S�b���c>���Wupu��ߗz^(���ޘ.S�W�r�@�m/Q������~[5��>@���k���|0�Y�pe���{�H�q��L8��]�Gޫ�s�_yɷ#;����'�S%���_=�;Үm�Ȏ��e}�e��.r�i�e�Ἰ����e���̘��_�9������%/�o�6��Q� �*Ы)̥��Q�4h�A�(��­�!a�^aq���xNi�������w�.�̓�-zQ����P���{��2t;y��	�v�z�`����Ky���G���<r��q�2㳅^�����	�(�W��<|��8o�+���O�w��F���͉�r�����ޖ/�-�>���yg�y�,�c�z����d��{��9�QF�����GΖߛcP��^�:�ȩ'����>��oI��m��G�z)�L���{V��];��g�y�w�>?G��>}��;����4[n��0#�;ɓO}"�V��a;u����W�.J���Y���9^��ڵi��#�bA �w�Ir�}oɋ�L���v�%矵���������3���g/�2P�>uw�%Mח':�WǼ��7 �O;iW�Y�(q����W_yk����͛K�֭EQ����/3f̨�~��ѱ�]�}���ꫯV~��ϖ��Y�`�\p�%=���ǜ�����M�~�i)�\t�E�V+���w%n���v�o��A�w��o:Z�(�����mq��n=�-n�DI��~�O���fa�7�I��781p�E��+2�z�7X�)lq���n�7M�4�+.9@��T+��f��2e�|���2w�\O��[�Λ#߸qci׮�W0���ҴiS�i�����OJ���K�7���(J��4i�|��7��U�VI�x���+�_�~��������Ǽ��s�ܸq�Jznd4�Y�+��(��~R/�1.��N�]*�#�)�Ct�^�z޶a��3g�g���%s���FQ7EQEQEQE)'��+W��'�x�[�Neb*1:4�\g��ӧO�D�/� ������rdD�kM�D;�	X6�Q@EQ�a��]�[ߊ>=�[���bk�{�4n�H�䣏>��^zYEQEQ�@*��/�(��{��X��_y�r��g��ŋ����L�0A.\�x�夳7j�Hڴi�E�Y��9�l�u{�]wy�؈|�G��Zu������I������(��N���/G�\�[o��h�~�a�F���;"m���<�mq����ҹ�Ϥz��%9����m�`Јx�P�s�^�8���7�-n֯�X�>w�5�񶸡0[��t����8/�:�dm�}�[Jr���7��%	�J���~�m��[o��	�V�Zy��>���2{�l/"�k��cǎ^z�1�#�]w����e�]&m�F����(��(��(���Bj:�����^8
�5k֬�wD˟y晼�G��~X}�Q/���/�|P��N���K�t�=�]�EQEQEQEQ�(Z��>N�t[��[�n�G��_~�̟?�Ko�r=mR.I�3f�\u�Ur�9�x�ީ���_�Rz��%QB�=��-T�W��"6�v�k���ܹ_��(��(��(��h�ީS'Y�t������?��d�}��� ��ȹ礴������͓SN9�[Z�k���n�Iڷo�q���k̍W���?�TF��Ujd�{t�k�*��(����~��I�Z�
��%K�x�CQ\��=��C���v��_�B&O�,q�����Kk�S�[X�9��m�����-�v�7xky׭[7�c"�݈z��~��,��(��(�����\`� ����"�YC���|���9��|�Mo�y�i�ٸ���=o�{��M?��Sc9�|�9ıD��(��(��(�R>[$�����s�W��-W
�N���[o��#GʓO>��c~��(��������REQ�C��k�JR!���R���իW K�@�'�u�[�n]����r�Ay� Dѯ��
Q�f�2�d�ā�;S�a����N8Av�}��2�EQ�h�F����婧���ӧK��hw�v�DI.�f���>�I�@Ǜ���O{^�rz~(PG
?���~[����»�(՟c�l+��2Dn2ۊx���Xޛ�Bޟ�R%�����	tEQ%9 �ɲ�@6"��ߍ7��C�}�С�<ja�СC�'��ox�bmI��ޜ�/� ��~zQ�"]�]��
�U�%��>����Ұ$Ǻ���U�+�� ~��eȐ!�(��$���
9��<��-����V�B)Z�s�1^Ty���x��W��uI�7A�s�N;�4�!,�lc�rVo�k�G���(�f���^�̨)fܴ��O���EIӦ��q�/�G��F�/Z��K�۴i�(��(�}бc�*S���{oo(
]+J�$.ŝb�&M�q]T�`�w�|��Q.�z���{"�o�k�+�RzH�[�p�$��K�yD��A��dI���
"r�I��(�RS��&���B���_~Y��J�$N��&�������S�:tEQ%�|��߮R���*�EQ��ӱc�J˖-�G���(�ַo_O�(J!$N����-��ѷ���^�B>�x��4t�����>}�T�^�=EQ�d��l:��1[)��	t��sГ�4w�\Qj��.X0_j���EQ��r�,QEQ��O�ҥ0�bH�
��St!���T�X�x��X�[	F����Ϩ(���TGKI���Kj��X�]�9�1AU�FRVPPEQEQ��D�:� �K����b͂�3�4MV��R@?3f�(��(��(�R:'�5j�	a�$F�9?��вU+iа��4��(��(��(�'q�u��Dѓ6���;t� ��(��(��(I�i���׼B��dРA��'q�K�.�����'J��6;N�Ν;�Rs�~� iѢ��4t�5EQEQ��vaSJC��߉�� �U��'4HNj�,��@M��8��gPQEQEQ�Ғ8�޸qc�ٳ�̜9S�Ě5k<�ֻwoQjS�M��JMcÆ��(��(��(JiI�@����K�O��E������� ��F�=͚5�aÆKMc��PEQEQ�rS�@'����v}�u�J�:��v�=����O����Dt΃�u����b?\3�NQEQEQEQ���\s�L�0����;N��g���ٲeKO?��s^q�b1=���������?2n����۵k'w�}�(��(��(��(5�D���QG%/���,_�\Z�jU��X�b�'�O:�$QEQEQEQ��H�@'�|�1��<क़S<��������[��+��(��(��(��X�Gy�����2y�don{)�oܸы޷n�Z�:�,QEQEQ�rѬY3/�ŪB,E��p1v,�W�Z%,��K�zu�EI>��<�^z�\|������t�zܐҾd�o��ѣGK�&MDQEQEQJI�Z��k׮ҫW���I����(��ϼ�(JrI�@�6m�ȵ�^�	eDs�"�A�����+���}���(��(�g�ȑ�-w��zuf%�4o�\�I������gϞ��G����EQ�dRE��
��K�9�6��z���%jz��!�]w�W1~ѢEҴi�X���e˖y�'r?bĈȏ�aA���kW� �uPEQ���%*�^�b%�:u�!C�D��-��Ç��'ʧ�~*��$�*o���z���C��qһwooy�n��P��(.R��S�9�_~��x.���V~�<�B���(�������e�ԩ2o�<ρM�-"�ЧO�{EQ��m۶��N;��|1����ؿ3g�EQ�E���:t���>(O>��,\�P6l�E��L�`��{��}��:�\QE�ѐ���SOy�ZY�$2����w3�����0��#>��X6l��v�:���M;lذ��UD:*��T�d�*��??��Se�}��`{��w=��ϙ_C�/a�����r���gN��'�,�EQE���N����sW�����W_�1c��QG%{�g����/d�=�v�,��~�w=�xi���8#�4}��Z�;� �KQp<X^{��/EQJK��e�����Jf͚彀\��q^^֋�Ƌ�qn "����~*�EQ���{�GƎ���!��l���/��c�u�+���jѢ�7���d-��)����r�Jρ�]D�!+� K>�����G�?*�s���S�)(Ӆ�Թsg��/DQ�d�Z�nA��y�r��{KG�?^fϞ�
��xI!�y��"� �w�9�Q�PEQ����#��-�]^y���?��CE)lD�
k^����bl�=�;�s
�Ι3G���+]f+�`��|��Ş(竻JA�n�2W��$��t/$ֈdSEQ%w�y�/�XH�'��������($���:�	���<��?��+���S����p��I��K���?(J2�6]QEQ��A�Qx5
�N��c��O�SMu�j����ڵk�kFEf��_�E�m�<���s	R ��� ���'O-����f"*AD�V���SEQʏ
tEQE�����{��L3�0aBY� `��5��%D5�Ť��E�Y���t�/Y�$k�>"�T��G}T9��?�g �z��C�S�G穗"�a��!�S7s����N�;SO�&��(J2P��(��(5�?�0�}"�!�I��:5n��Ht�@:ԋZ��)�D��R�
t�`�O��%J�O���.�
�βz��\Ȥ���D�6m���}F�g+&���E)-*�EQ�3eʔ��9i�$I�$�O��C��&�������=GB�HyD�).g��;�W@�O�8Q�N��U�&���;��ùB�^)-Ů{N����s��₊�$�J"�EQ�vm�`^6������>��4֬-�F��e��բ(J�0�9���Dr��^�y�N"�vM�N��u��ׅh9N�b��݅�_V�[�.ӦM���OT݂�`�w�O>�������,�ǆ��{IT�� ��P���E)�H:�.� ��ⱽ袋�:Ë��o�����T0^�2|e�B#	Q0a�xQ�Ccl�:W��D=���׊ �ҥ����^7
�`�}�VR�Yf������b��3ŀs��޹�D���@��k��N;UF���w��������͛{�Iu_�����Že��Ȝ`*��(�&��o}���r��R��1�뱾��$C�����y"]��l0.�ㄴ=}f%:�r3~g*zU,̳&M�0�v.."����{�K��/�IG�@_�6���e\�L�	�������.��/6�̙3E)/�s��@�:S�J!A��i�6� ynT�+J���
/kR�e_���,ҳ���TE�4�皞W��}�Q����s�-z�w�4l��(VM��g+j��(��v�J><�1����n2~�xo�w�@8���x����~g��
m��qPd+6��`̘12l�0/{�B�8~7w�\Q�����:S����⋢(J�@z�;z�����C���W��'�.X J͂��V�[k�BZ�?җz��^�(��$3+%�hR���}���8`L1b�'<� $�t��e� ��!��$�UZy&��s��	G�Ǖ�@w�ɥ<�m�ر^u��;z?�I��Z%�,�� A���}���B ���oP��D"�ǍW�jh&� zꩧJu'WA�ڳ�����^��5h�Jua��Үm�{��RJ�Qt�0��#W�#rI�f�O��Q����ӧ�����+�Ě���EDڮ�TڎS��_��q�k�7΋��u�]+#�O;�x�X"�52;(��_����C��mZ{�Y/8[2Մ����{��o�-�Ԟ���H:/6EQEQ��z����}�~�K���tJi�O?��g�G��Q�P��1ɺ��e�1c���=r���y�""�QD��߿х�b�y�5UHwF`ٶf*}�H��{�Y��@;����Y��?����B��B�h�Vr��""��q�T%;��(��(5��|�<��Ñ���#��*8
��F�g͚�s�7�1��mK��Ca8���>(Y�K��[g�o�2�I$�f��i��ٳ#s��t�M�8�2K�{�sBA9j	ϷQ��w�]�|�M�Q�B��ٕ!��Q��(��(5�����[R��i1�vEp����|��/��1���<)��������ñ�l��^/D>��z��bwDW��`Z(SK��r�2F�� ��`�"=�U���7d)��]QEQJ���ɝ�K��SN��B����O����.v@\�[�n]��Q�\�����v�w�;[4q�h+dy9Λ9�6՝v�>��X8D�������8����E�B��|%�����`"]k(J�Q��(��(%��������A�?j�1jGc0ǳY!��~��#�<"���z������Q�FŶ����f��\a�7��R��b�0w8�C�Bʞ�k��V����ګ���e�lf��������8oΟ"qڧ�0���s�����';��q���-,ga�B�� QO�G�g(�R:T�+��(J�X�|����Lo{��	r�:u��R��D��O>��L�<9T�#�w�a9��ý��qC�3
Uɡk׮^�?עkݻw��?��B"��@`���T(��D�9���,O���/"�@��o.K�)���5|���W�Aܳ��"n�
�b �c|��g�(JiP��(��(e���'˽�-g���$�,�t"��|�'��?�?"�r�9���L�:�K�"�,�6a����s�?���X�{&܅
������ܫB*ss���3��B;�^����R����<g�S+�+JiH�@ǳX� �w�? ٗ�Ҷ2��Q ÿ^$/s�+��(Q��K�)�-��MO
̱}饗�NF����˕��U���$�Θ3g���ܭ[���P������_��*�sGIϞ=c=F6�^���҉Z PQJC��~��'�>�lA����F.���*?cN�c�=��gIo�#�w;���r�M7U�����?o��(Jue��M���E���m����X�.�(nu�q�?nH#��Ԁ��r�
*W�À���6C� �+ee�4��_
���ر�����S%^'�K^૯�ګZ[�h���{#��'��EQ��<�mIdԨ�Juc��F�j�#:L���9������i�j)�s�s�-_~�����5�Qo�Q1�7����@��ݭ�_D�����vzJ���� '��(�Pc:P��o�q��IM�宻�"�����u���IRH�夐J*)�( pP�"�}�^i�\���p���*
���
HIH��;	�����|��?Ι�ev�������g>9�g��ٙ��+�OQ���ƾs��&�q_�[�j�*k�;"��Bf�x>��������!B�,n����w�����B�$������?$P�Y �^�NF���M�6��pT�@�D�ӟ��>�����!�H&G�hb|q�]���I�O�����C�]ٳ�8e�e޼y��D���t<n�s̋n'Н�_�Yo^�ˍ��$Dj�3�����*����@���N:)��|z��Q9rd�_��
�]w�]|�ű=v�=
:WQwڶmk�gώ�1�x���+��/���.���pۏ?og�� kղ���u ��o��9���
h���㳂���"(���7��r�-�����7���q�����v��eB��P2��B�:�����p�	Vn� �/G�aŤ��oB��gwȐ!�D�w��*ez�he�[a"R��Ҳ����jJ�9�ad�y���t�L߻woo|\T��$eU*�^����-��fƗ#|%Ѕ(%#У�L;'k'^�?�x;��S��g��r��m�24q���.�I};�ᡱ<֧��q 7�\q�)i��2�d��e����;��._����1W�{��W#+u���CR:����οu�c<��-v�}R�� �6 �Kl�m��}�ҥ:>�Ha�D����&�P ��Ϛ5��=����Ȣ?���e�L���Q�q3B�J�����u�Y�
��>��z�g�g?���EL�X��/�~���`7�p�%�GyD��ĩ�Ae���w�{�-[敠��S�[�lٜry;$i�IY����7h$]Hgʗ+|6M�4�q��\<��WT����>���(��"���@�Y_x�Zn�~�%˥��G?���}���'�ؗ��%{��G�\�&Eم(>�ׯ��Ç{��"0n��!�7n��]��l�/�J�}�Z�b�0����c�f��z;RCɺ\�s	F�8�:DY�uh�
&IiDO�j���y�W�uI���L�Jǃ�f�u�z�%Ѕ(%sd�v����eժU�����בUz����,��=�\�*����O~��˅p�B��zn��K����?{[9���k�B����\3-����xu!�@�3�իW�� �]��u���+Ѓ�#	���+зm�f�;w���~D�L=}d%[�,t�;��K/����>+G�V��.��B�|	�e�*h�����Q��b
.:�.[�>�`eˁ2i,�Vh��Z��S%�JRڤ�(G*Z�oݺ�&L�`�^{m�u7�t�=��CV	��5�!�-�"j�9'����ik�.,�y�Q�]�{I*G�2�'���|Z)��L���NЗ �00z��H�<��kH!�?(�Ny6&/�ȷgs��.��z�'�#.��r+wC3��&����x��ߛ"��0��O�yn$y�WL?���|��&�"����Fl��9�X�;���Đ(*�B�.�,X����#���.�lʯ�y����ri	,u)�'��t�c�=��%t�z\���H���+Wڼy�"�_�8��.��������BQn�~��v��כ��3g��JEr�?�oǌ�0����6�]�6��,��?GJ�Ìq3fL�ƍ�l�`���`ٶ��SWK�'� \0��@��ר ��S2���������Yu!�(7z��i"�W��1�O��̻�P��/d��#b��[�?�<,����~���s��?��ݏ��K/�d]�v�N�:E:y 
4qB�� �~Nn�2�?��:�
!D�qH�F/&�W",������;^�uoN���k���|�	�hѢ���;O� (E曖�իW{���/S�;m�܆ϫ�fn��*D��@�_��^����W�GM!ʝiӦ��X�0znذa&JD%�~�@��2sL�p�.��)�؟ɮ�Sz��ر��@�8oŊ�?e����e@Ԧ���cl�@��@�Dtd�W]��P2�2�l�5k�佸�@�"�w���	!D��`y��M�]}��&��P�>�h�g��-ZT�;�G�>}�r�t�E�:�d���9'`1e��\�T> �Y9S�V�ZD�#��p�����,	І0�|/p3dȐ�����/D�(��\��e<���@8p�	!D�P��.�_�k��}d�-���7�eCe���/_��2S)@t�)v�/^\������:o�,0�|&\Q��oX��/#�׭[g��� �2U�Z���������x��۷�HN���~ń}d�������8�;�? D�(��pn��F{ꩧLQ�����k�s�ڕoY1itP���UY%�[�n�x2�ݺm��3�d�����Q�J���$���&�>`� O�DY����X����s(sw0�]�~}d�߼y�n�d퓒!N*���s?�ۆZ��
�.!�C=�ĉ��L"�B��e�����í^������|������wl���c���t��[kL�~�2D2�Y���^t��d�Д���޲eKd��4��+�G���G�����@���x(ehy�
�ٺ��;�m۶y�n?͗|��	!8�>g�;�����T�8_y�Z���u��/L9�(̬U!Dyp�]�z��s�7l���y�G<��TB�%�����]��8^��mzÆ�(q�ԅY�y��~xz��2�.��s (��6#�������6T�?��@���0u���ߏ�
�(B��$N�}�r�,'�\���R�BT���T[�d�����ƍ��5���D�/_�]�g�(g�������vbD}��sLu)>��CQ�����'��(��x=~^{�5y$��
�(zԐA��
�E��Q8'�E|P]5:`!Dj�i�M�����]ۣ쮛�`c��0���ڑ�����k�z���w8��5���7�I�9%��o�@D?��
c�^�zy}������rP�^W�N��R}��Q��;TT���r�Y� ��o�UPQX$�+������sРA&�"3[�����=�������M����?�z�����Z�i��/,�0��0�ҥKu�cǎ�P#kYH(�����cW��z���9��#_���@��`I��{8�J��5�@B!���~l��v�M���L��R�Y�fy����v��\&�Λ7�PO��_�j���ׯ�:ƷN�<����Ɋ"	 ���T��~gf#�
1?��a_H�@�w�ߟB���@]!�(k�6�Z���~�嗽tĨ_Df��2��l��?�C�;���M�z�)�?��c=#�tlڴ�:�4��������N��@=��۽�����]9B+E]]ӹ�5k�Ժ�J�Q��ѭ[���֧zB�h�@B!�D���L���˖-�+Vx}�q1����j�x1�"�G	x\�f<}���:��<�Td>AW�t�A�ݵ  ��������^˂4��0����
f�ق�o߾�@�w�} :w	\:�.��]��#�.�B�C�g_�d���A�"H�(Id��:��Yz���pB/�-�p�Z��-k���{��q�����p�3���!(&!
��B3͛5��r���D�B���G�	_�ru2�;��;�Nƶe˖���ɜ�9�?��H�7a��c��A D<H�!�10rxW:������N=��5i�)�A/wT}�����H��9��]�v��1"�q��^|�f]�@D�����:��}������ �p������9lذč]�K�.5!D<H�!�1p�wO��c�L�ϸq�j��օ�S�dz�����;�I?���E�ͬr�� �����̑ǭ=8��ӽF�E�+�={��R�}�}!�9�"Z$ЅB!
"!�i����y��@�e6��`׮]��)��= @0`� O��af��E�$�ī��ꍿk۶��T�ȃ@�x�@B��{���c��1_BTd�1�b�;c��� �FC�1Nm�ڵu�~���;��|tJ��%�fv# Ea!XC`�y��d�`,�"^JJ�c�B��E��b�䆓�g2qGB�� �$D���۰)�R�J˹?,�q�g{ˍ����7�3��H,\��O'�Mz�0�����E�;cܸo�{�M��Ο?_&`1�����ٳm�ȑ5��$�8O7PQX/����g��r��1�FYX*����-��+{��"��BT���8q��Ey���UN,ra��%}ֹf�����W�`k��#S��_��}���S�L;p\;��S���v�c/��͜9ӎ;�D�t��ڕ9�x$V��5�.���4Ȩ#�پ����ĉ���K�|T!D2y�WL�L5���Tb3����!D9;�d���9�A�+dÝ@����37�Eq�3�6m�g�GB�P*���ٳ���9s���A�l���N	.!�K�:}QW\q�7��.p�;묳��N��������{�gB�Xe�و�y�H�[eB}d���Ej�#ɚ4i�e�Î)kڴi��*&�ꓱ���S�N���"��<�TP9@�;n�Iy*>��s�z-��J2���j�F�ŬY������$J��{�v��WG6BȪ�k_��N:ɮ��J۰a�	!��.}��$������v�-3!�B'�)�g;L���G]���Qd%̳a�Hg����_�|���GaB'��j
|r�Q��A�s!�A":��������;�`�AT���n�A%�B�j�~�i��K�QGI���_��&��	"�s��՗����Ƃ!z�N�p�o$'8���^��~�{���o@^�S,Y�Ąɦ����/�K���0o������G���B �;6!D�ٶm�����݁W��p�l&��r�'s޸q�����Ѽ�ش�r����(+T�������8Ĺ���M7��E�.]jBQI�@�4����H�)=8?�� ��'�5��O�w>��Ts�SA�R<i��!�"=E�g�y��w78����?��.�(���B�#'B!��N�������M$��g̘a���I��h�s�B$��l��5���B$��	tf�_����'��Τ�߭\��39�̂3e[�j��cJ�O?���ѢE��l����M!*�}"z��"}���^?zǎ3Α�,�u���,Dq�s�{���x�T�/�(>E��8O�O�X�L�!pa�;��Y�n]ڿ�G-->|�W^?}�tB�J���1cLd��(9�ӽ�Sǣ���G��������;"�
9~�����o�m���3!��s�gJAP�㭀�_.кLZ����Gyd��)x%Dr(�@4h��p�	���>s�LE�(a�t�b��~�WI#j¢���ϻ�X�x�no�����O2av���W/Z�ݍz�7��x;�*����\��b<׹�B$	'��:�u���Í�9�G��$��(6����CЌ \���$��WUU�g?�Y{��gMQ�<��C^��H�B�V~饗��s���7��Mf'�x�q�&�qC�-�m۶�&�̝�P?��
QL�UH�3|�!ЙG�GZl���/H�Q1�Dfh��t!J2,Aw�`�� K0в{��X�z��D2��:t�~����ٳ�8L; ���2�B$���)����ȭX���J�qB�&I;�$�+>[��9���?\�����:8u����� L�B��1�"�lܸ��[��^�zE>Þ�LS=�"9�.ЇfI��+��o��	!J��'z*����y��=��#ּy�з�������X�ӟ�$��)'���N����?�5���u���.<w������4�N�v�����#�17fR�ҥK#�Ib�ѐ!Cj��}�ݜ�����;�]�����?Zh�4
���rowྊkԏ�}fz��?ޖ/_nņ� �YL�<+D~<����G�d�:물z�ƍ�-,�EFm��/TR��ܣ>ׄe݆]v˝��s/��G{�2�B�j�-[�IY3F�q�dҷoߞ�P���Oi{�o���2J"a�?(�0�-	�+�\r����رc�s��.ԁS!ʐ�6گ�g�}���L�cҤI�ZZ���"nذ��uTKQ
���{6o�<�[�}�I�&^�wkz��=A�LkC2�l�o��� @�^�,�6]��� �����GyĦL�R0�!��a����9��1.A.J��;w����~qW�Nh�,x>��\�b�|�H(�	�h��]��\p�w��@"w�8�t;��sCߞ�;v�$@�M׮]B����.�}���+���	Ȗc��)�+dߩ�$/�H&��{"P�"�������'*��$>��Cv��9����e/�@ӦG����Փ�X�q⸞&�Cѕ�{煏>�����D�ٳg�M�<ٛLУGo>z� �׭[gk׮��!Dr��[����Z�ψww?��]ֈ#Qh~x��	D�@\oܰ��*�)ʏ��u��.m"<���g�K~��І)�m۶m��R��Z�h�	�t���T`����f���<��6L<ia�0GA�!D2�Q���-ר���($�կo�۴6Qyp��ڭ�m޴�>V�K���׳��-�������]��:���ְaCo�b&�i�&O�3�
ڴi��FW]�o����	!ʛHz�%�E��w�n�>SQ�t���v�|Û�*D�����8��Dy�P�KFq��KwU�:&���"�(�"ZЄaL=ˍ����)�I\��މ{	�pt��-��<��OEv_���v1!�eˣ��k���&D)ҼY#��Av�����s�ze������q;�j!%��&����&T�LL��$]�%��w�{ ���0a�M�>���Cd�[oق�[&b_��y=������/���z#sa�9����bp�w�ͺ��y����'���*IB��~��'xV�3ƛx���>�4^!�H%)��E¾�S�|�a�{�y�?�7I(�fq��kX�fm�^C�6m�~��U���|��ެh��;u��]��=z����T�ߗޡC�TK����:�(��66>cZ��0�9���y��7m���
�
!J������BQ��u�����e������y7v~}���Σ�TC�w��ŘTCEVӦM������A%&~-Z���y�1��ќ�m߾�wߣ]�v����m۶mi[�"iH��|��B��c��uE�Vѳf�{���Qj�v�w�G�m� ��s�NɠI�&^@�y	D�*������D0|ǎ
�	!��B!J�L�fdJ�N�jC��J�Ӂ8[�x�'�Eq���k׮ֲe˂>���F�k��f�7oVE�H$ЅBQ�˝)F��	wB�R�)S�x��-h������5^��P�NK%�q�{����{��W�!�H�B!�(	�N�#��������[�PgC�S��F�4%�d���A���@1`�6l��S����!DR�@B!DI��w�U�kLV�f�:Yr���=1��b��B��az�Lǎ�^p��|�3����l�bBQl$ЅBQ,\��Z�j��ts�ɬw����ȸ�]G�#���A���={z�g8��V��M�6Y�@�{챉Ț���g���^�=-�MB	t!�B�[�n�6�ի�'�3A��~g��L�ˬ3z���B��9r�7�-.L�b�c.Y�Ē s�)#O�3c�`cd�|�]O����c!�13�-��m0{�l�
!�F^���;8rr� �fzsR����6�c!�B��	��3gzB��:�<U֚Y���fC�]/����!�?�裂�8��r�����ݻ��IG,��oi?�� 
^O�`
kO���F�>ג��͛ۨQ�l֬Y����lx�G���~S�*-��$'�N4��0�y"�<�8	q`�DH$RB=y�9=��Ñ��e�MQ�<��Sָq�зg!|�@a���B���G}��>J������2��k�z��T7Z��Z�ܡC��˘խ\���eӬ�(�&8UUUE`��#F��Y��d�������`}�3;Az�Ɍ�a�"}����|hۈ��B$��aNS.�[uN�D#i�"r��=��cB�����7Q~w��6���Yo�w����I�+�$X�`��I[\���4�����:,X`'�t��؈QʾY��B2Wq�0g6���j���֭[��/A�"p��!���rw!D�����A�$��oz'�8LRDeAI_�Q����Y8���y��O>)���b�#QJ4n���:2�8�� $!��sɘF	�l#��u�3��y�-������И�RS��q�FϿ /2�.��	2�C���'4B�EV��ɥ��=���s���NB�^z��3&�����P'���:��ի���C�b_|�M�<�+�+�5��5Ѥ��O>�8��ݪUK��}7�k�뮻L�׷\�c�(�ƍ�z>�]�vy&qd��_�Ž�/� ���j�d�I��u��m�%�LI���-]�Ԓks_>A�*U���&��!D�OT��T𻨢�(ȶ�}� ��q�Ξ��{ݎ3�<��ϥI�d��M�G�y�}�nݽ��b
t�#�?�u�6+m>����qA��W^	}{�:��$@Yf.��0��|f�� ���W_m�&��Pɂ �ː�=��z��׫g�ʹ��	�e��q^��q��$��=��?<�0w��&�T0��27���'�lB�Ҡ>:��qP�hu6p�d��I9)=��|�sP�'JŢ����Y3���C�j'N,�8��֭_�����x%�^{-os��{�k/�4i���"�<���w��&�q�1�Dz���y{�ŕ֧W;㴃b�(e�r���l���.NPk�QI0	k`�9oٲeE�R!=c��iޙ�e�v�&M*��B�� '��QXʕ���I��{���a��'��ؼ��;y��|�A��YY����^����Q%QӨR%��j���x�v��[�|�n��t;��L�F�Q��s7%ӅtL5�\:p��P�]�z��X��Ʃ!ҩ&��1�ד�nB�7�e"=IY�8��DeC9�!C��I���4Y�CQ�$?�s�λ����{�ڵmj#�w1�8�S��F�{��UWݻw��A�Z�Ĺ�`��U�����6ڦ��B	�2��?�~�9�ؓO>����z�wT_fA5���E������hؽ{�F˼�+��}����
��<�ch;)$��z�������?6Pj��[�d�.v�֭�r�{������fH�������rZ�>��_�!���Τc>�5I����ٳm�رY���2u�TB�B!�.J��u�m��J1������
��}�C�U�Y��ز�x��RdM�I�Z0"E\q\"����Q��5!{�m�.��y��%��*��)w��r��(B�B �.J��6mL�E�=�bC��]�vy�m1{�1KJ:f���'�y=�lٲ�D��^�j�r�cx���>�)U�X&�p�`*������K�.YoG�U���Klڴ�+e�DUUU�:�+��0Q�H�W(���ӟ��~����O�WF�:�rHB���yO(b�!uxޔ�F�W\��{��P<����#����qcC�v���$A��ag0���^x��ŧ>U߾���&r�є�fd��9Nq�֫W/o$�ʕ+m�ڵ&�N۶m�f����O>�k#�N������ՍM�`Ѓ�[*�/��Le�"�H�W(,Z�9��C��(y����K߽ ��šy����fM��	c�����y+]�t�~������>�H��SO=emڴQ=,�r��{�5�X���C��ꫯ�}����	�k��v[�۳h-�@�ҩ���ֳ��mL�F�N�<q���!��}�����_���S�F@��@��6�m$%�<�@G��Z>� B�����{�V�|�����#&%��G	ʻ�;�m1Ӻ��+M�Uʌ�$s���lԈ֧W��w=(R�SBಝJ��g��s�s�'�N�{0ˎ�ܳgOQ��>���+��*c�%�qҰaC��c��LJ�c��ȔE��"N�.���s"+�q��P����K��<���B���ү���c�L�s���2Fn޼9m�������J�dG������"L^)gl	|�dr�'�C[��yN3B�tԧ�+ݼ`"�Q�'QZ�K`T�#�I�q��&��<��o�!�������ܱÒ�f�җ�oݺ%�~H!ↀu�-�/#�w����>�)S���ѣ��\s_|�v$�{�T�	t*�J��%�m��c�� ���g�A����D�um�|;w�u��yn�B�dS����.�,�/�<���?�zq�
�9��3&�ue��A��[��E�'�����%�sϿ��>�������l�A"D�BB�_NKKX�+Z�0�:�㪯#��C=/���T𾖺�8m�_��;�eDoж�k�+�'���6��A�c���{/��Y!J��&q���o�w��E��Q��/}I���A���E���Ӽh!�(֮Ú5U%W�p��ʅ`?t1[Ȗ,Y�rM�;= ����O��0�!ۤ�����#�@wq@���'��`�&�G&�O��aÆ��/��	|!D2���N&k������'���:�+o�D��BQY\{�9��5	��\�Aïb��*�$;�4�Ø-	�J�l��9\̅3�z'3�~��QPxG��<�p�S��U�V�"����H���k���\C����w\p�<؄B!�^_ʦ�0G�l۶-����ݻ-i�G�R��'�(��]6�N;ARF/�f�g��K����79d��e5��0N�* �{��U}=�$ЅH.��sb8����㏷iӦ�ܹs��]�A�L���=��Ç��!j~饗ֺ�����&�H��+������ʤs��_�&>�r��7�� [��k��.��~!p�և��2���/Ȁ���b�xg��o�\���k�ԢIeC���?� ���A��U` ƙ��+��"ل��ܧ�r��q�#2G���8D����{J;�����_�H��w�iFg%���I6o�ܼ���O�a`s�wد��?���>xߊſ_����0ˇ���ͮ��0���Ki����W1K^���;�d|�V��Q0Y��[g�>�`���׵kWo���̯N��Ǟ��*/��_?��$��:�d���T��g[w�So3�1�L� h\�0���A�q_� �
'�+}�(Dҩ�7�FǎMD]�h;4=j��9���3��8w�.�^��{��R��Fz�y������z��K�������(������v�\�i;.�� ��8�;s�ٳ��	Sz](���8���$)��	V�R}�lV���g� N�D�Z�BF��c��%Xb%D�/�c���D*��3٬y���6o6!Dip�1�x�<�3�&Tĵ;�����ӱ�L��8`t�Q��2w��;���!8�� I�c�dHr0Z!�.�� :u�h'�tr��L�6�.\hI�gU�u�>���K/��4��>�=���Б#G���� �D��B���q�F��<̡�4�W�j�?��w�^��`x��H�!ʞ�+_�q�>1��g̚�hq�׬�֭ۥ���_�"=�ʑ�v̘1#��g6Șo޼ٖ/_�#�fϞm����!�d8s+Zylݺ��8��S��~�O���WR�E�44V4$Ѕe�wmڶM��z��6O�p���ʭ�S�TP���:A��\��9b
7�`_9�˓&M�J�Y�R���ʅ�r��v��e��{���5��E%m���&�%���^���\n�^BQ��u� ���謷����H�رc��2B��|�z�q�7�l���r	sL, ��\�T��arp����3eЅH6�%�իW�B���+���c���������B@�7����:��X�<y��jpA��iǢ�e˖^E	��<���<ձ#i���@B!DI���7m�d۶m�Ԓ�Ĺ��?ڇ�(_$ЅBQP޾}��#���o߾��YuzqU.����@B!b`��m֥sk߶�կ_|��Rd͚5�Fi/Bì��)zs��ֿoLY�L���B�� �.�(+p;nݦ�}��?�{`����H�7�.ޫ����ի^��>���5|r��[o�e���e"Y���g��;�nGq��{��v���~�Cy�U���޶m[O�7iҤ��pjoݺ��	Q�0*�Y�f�������	!��z����SN9���,ę�*���8���;�^u�'v��/_���5�f�S(�����e���«Q�ƶ���]v���	j@ �r.�w~��b�T�~g�����<u�M|�2��:�>���\�e�\�.�@2��$ЅH.�%��Ν;׺�l��&�Ʒ�~���*�=o�����|��m&��5;m��_����&��/�	�1��~��
�!�($ЅB�"1s��
\�ٖ-[�SO�;<(V�B�		t!��0�%�}���7�xÄYӦMc/��ԧt.4T���k?�%杧�~����.n��J�$����t�x��o߾��ke �D�=j�PvdEmx�
���3!�Ȇ3ELŉ'�h�5�~fjA*o��N;�;��Tv��a{��5!�.��ܬ�ӦM�������߾z�p�E]< �?�V��!�"$Ѕ��X�n�����Dv֮]�}�nu�����.��;��>�r�/N>�doZPƻ`��P��]�v�^�zU_ްa��X�� ��>��98�������������#��5B��%��V�\Y�zp�",[�n�z�b����/�-E(iw}�dy�����}fl/����?�1,Yb7n��w�ׯ�L��iưqN-D���7߬���#8@`��`|7`���kfŋ���s����	"�"�pOգ.�H�%�W^yń"
�0y�׼����{ѭ[�������3-��z��x:����#Gz��4c
H�;j�}�]oƴk'�ׯ�u������o�Q���f���`?�߿�-_��3ܢ7�B�"z�>�h�zhȐ!�gLÆ����*�fΜi�'O��>��D� �.�B���{����=]v�Rxʾ4h�]F�B���ŋm�����]<V\��TSY�޽�q�N�:y=�{;�ɇ��o|���/�F �1x�`;묳l���v�-�؜9sL��B!�(9��]��a۶m����tB�xw���S�N���<�8�ymdΩ�A\e�iӦ�S'R�s�M�L>��;��N8ᄬ��eg���v�M7�s�=g���@BQ͝w�aGuT��?��_���$P��!^6!,|�]~��?���֪e��V�*��ڰaê�����3�-Z䍛��m�q��b޼y����2`Q���{A�{9��"2]B�ƍ�
�E@����F���z��y睊2��u���$x6���E2!sF�;V�x��~�z�j���B�j���c͛7}���淶o�>K,��X��}�,^��HS�*Jf�f��zn)�D�q�g۷o�6��s��5�6�y��g����ٶl�����a>�V2Żv�������y0��{������ċ.���u����Ӿ�9�c�=��Kw���������2Q�H��|YT�z����	!��T�d�9��ݻZ�0�>�,{�ڎ;L$�#�<���k�.�j�uǠ�@^�`eE��8G�3�����*�$���wPR��g�Q�=��g���n�-�d���~�7��?�x/�U��y� �^"�;|��Z�s��@BQ�P���Q���	�W_}51��;�O;��B@�/}�l�_��ܲeKY�z�]-�X?QXh�q̝;��-OWBP����=��#��'�>t�P����f�t�@B!DY@I�I��Lzǎk��"���mn�(<��Ӓ�KKM���"�gϞ�t�R���������X�j��҆c���ڞ���_|�N=�T�k����B!J��Ntc�
Jz�e4=̈��9������
Y>(x��n�\��LD�/[�,e�p)@U A  %�^������wN��b�*���B!JJ��B6�Գ���V� r�]�PZ����*I�D���ZP��*	t!�BQP()g+f�<�l����/���]$,]U�oaZrZ�jU���J	t!�B�,��"�[�n�m۶�Hr�A9��|!��j|X������Z�={vE�Qɂj�÷0����^�6�%}E����T!��R�V��d4�af�9cٔ)-,��#(!��=d1��s��ئc֬Y�z��#����
v��ǌc3g��	5]2j���/�O<��h��������H���(m$�KF�=��c&���W�.�m�j��axb���7�<����m옪�����ƌ��Jf���^9r&�{͖��S��|�h�sb\F}�@�-��d��m�>w�{��g���@��]�v���~d�G�eӦM�Ɩ	'�w/�����K�,I{��c�zU0y�d����B�����<N�CVדּ�I���O��V�7�ʗ���;vd�-����b�E�S�@2a�+d�q�g�9B�O�>�����#Gzb��I*�v���G��������kC�����7Q^H�!ʊbD��}�ⴿc��X�#ɋI!D�3p���U��7�qR���/��!`�i�&ϛ�r`f��1�#�I����;��Y�B��B�B�dEoX�$МU!DB 
���.����l�\��Ea�ԩ�u��1�m���oF ��۾}{�qo�3}���Xb,�Q"�^� ������~'L�`B!j��=a}�t�cz��/�5�:wln"(�ElQ������<(���S�\���s��da�������\��IIw�g4T���Cݖ�nL�����L��eǛ7��=����7ߴ-[��B	��(o�֭k]�I���B�d�f��y�;�܋+l����W}־���M�2阊B*i&��>7hР�2F�8�gk�AD4�Z�3N.��t�o�t&� �U��Jf̘�e�۶m�����HQh$�KH?���׺�2��'�B��ᣏ���xֺvin����D�@����*��0x�֭�wa_�~��:4�NI5/���$]*�͛gC��*�i�b���&��D]!�(?:W�A�S^�h�L��ׯ__-��L�G���[Ҡj�W�^YoG�õ�����эc{�r����{��\K�B	t!��#,���T"�D��7�|�DeB����3�t�͈ZW���,�8�ѣG�9�.[]̲�t���Ν�͓�6��w��6u�T+e��H6!���B��a���I��֭Ï�E���{_Expw���RpJ����S}����! �sD��Lz�1^)'���������X�re�=s��Lz&8��J����h?�B���`�B$	t!��#d����b���s���w.;�Dx����J��P~���ي	���Q�FU�:mٲ�'���3��&M�T_.�xԺB�y��9���k�Z�A��e80K=��j.f��W@ 1���*.!J	t!��#,~p\Nǁ�X�0�/��V�Z%�T��a��9��>*��zl'����i]:i�Z.$� -p0�=�Nv�qy��=~�+�_\�<�$���gcѢE)*Id���a\�`t������TT �]f�,y�`�"�H�!D!���ϟ���z�V*�x�V���/����F�	���9�={��!.Z��g2c�2�8��1�Z"�ƍ�	x�U�D�~ ��m��f���3A��l6�;�V���`_ +�~�2���}B��A�D�w��u}��5!D|��n׾}��'I�������c�L�废����/�W���/����q�D�s����]F�@�W�.z���!���5��JW��q&ie�a��q�ب�ˠ{�����[��|(���Iv����wI�BH��\�4�DQ����W�b¼��H6]�t�qy�ҥ�`��;��[2���v��٬Y�2����	�N&=[&�@}��}BȠg��������7o������;	e�����A:B��
�I�&G~�7n2!DraL}��̃>h�6����6m�T����z���ߧ�~(2d����K�-�����+^�9��A��^�f���M�;g3�C�*f���Ul�A*C���yҼ
��!�^�P*w��כ���ر�~x����>I�}��G���#�����;�j�/��s��n�Z�68�����W_�~�<����/������3RLW	��d�1�"�OfaNb˖-��O-Z��z�m۶Y�����4{��b
tLd��O�0�8���@B�:Bc��ŵ(/�v����9ǺTp���)�J�]���qM8�Nv<,��J0�_&�|J�5���L�ރBC5�spwB��}Iu!J	�
�u��֭[����B$����Mdgɒ%&�Cа+X��9��b~��8���Ϟ�]�vY��M����8Z%hs�����S���v�d��/����2/"�H����^v�e��'30q��P�q�=����!��_LR����}̈́��?��?v�/c�D��� q�9��A �� ��ā����l��s/e���>�т@f��w�ws���y�|h�`k���F�X�`�	!���BT0��N��ad)B	�H.A�DE�&��.XnLﶟ���b`x���R�Oe �|�	�0�C^�Ν;��@ݷ��*艎��W����
�Ȣ�#�}� �?PE���v'��ƠB$<DTش��&�H��)d��)�J
i	!���!{���={�Ly[zn�e.{舻�S5��2�-3��kd��k��n�ƍ�{"ԅl��u���;��qB8�L�Г�*�>������IZ
��J������@�"�d�A��뮳	&d<��Q�n�Ʉ�Q��1#i��\��'W�^m�t�`̘1Y����k�,�:t�P}g�;�+�y��>���	����'F��������tL�($|�l9�q�&�(]rVnnA�8+Ȋ��0���Ƅ(�,RQX��~{��k,J��
�$B�d3~��9<^}�5�)G�L��_�o��{��q&JJ�i��ӧ�W&��a�X���6I���8�Y�u�~��t�^s�-	�H5��O�3�T�#Sf/�@�8��q��l���	�p�s���d!D2�I��\�����?٦M�R���4���������?�|��"���7I!�(u�d�݈����r}:���e+�{��uUe%DB�ei	8���_!�P��~�ڵ�0/$P2o�<��-[fI�*��0NΛ�����}��6	!DzB	tN�<�M�:5�/7}S��~��>^��B!�R,s���y���"�.�	 �d]�t�.#֩R�]T�;���Ȏ������ƨ	Q�d�Du�cη��H���k�_}��5"78!?�쳵�_c���$��o�{��z��nzZ��2��V~/^:���k�ҥ^)�+�ޟ�lRQ�N����B�Y����:�<�&I��+�4�N���rK�e�_G����BQ�����6vLU��!�Ej�w�Z:�]��᠉b�}و-&���e	����VR�/�JȠ��ڵ�h�B���O�÷T�#5}��H�����z����F�J��%7BF!��o���Z!^
-Ѓft��.Z�(t��]Ʈ��?!�P�ɧ��ӕ���we�Tg!�K}f�>���<�q���n�Np�~%E���ц�B!J��lNd#�[�l��sG0ѦF��ͫ��
s�1��C)��L0�e�����"l5�16���f��"B$��Ȏ�����ID.���P����'?��	!�(m�L_m6��=ZYӣx��l3p����n&{�#P�6�/��Ll�8'����>;n��`8'�H.!ЅB�b���l����[����ԓ�؏�/ֶ͑&�3{���#R(w��C��O�V�����?��G�<_�+�`Npc��6l��]�*/��oT`H�Q�H�!�1��G�g�ٜ���ǿm�Z61J�S�K��6x�b��-\�Ы��ѣ�'��B92fv���j0'*�3ݘ�u��y�!�)�G��?�=�u!�
�+W�Q)P���,
�WB�3o[R�Oy.a��b��	!�(��x���;�~v��LDK*#��uq���ԝlz���~`DS�jݎ~t2�;w�-[�$�=O�xл��?)��H��}��J������#����@��?�r�� o�3�(6,¾�N�B!ʃ�7��;��r۶m���~�t�S'k�Β�tN�YN��J�Y�j��(�W��!��BhB!D�8�HUIE���L�H>P��(5��9�Y�fշG'ad�C��B!�H�!�E�3��;d�)	��q��G{[*�n��e��(h�V�䋿O]�<$ЅB�"��KF�� ���3&kk��py�fV:��2����O�{X���2�	��ڵ���"�H�!�1Ьi#������lm�;Ԇ�얨�uʔ)ַo_�s&8QB�|ٲe^�=.���j����5~������C�״iӼ�B���sqO��D�YIT%�0� i.�B!*�����6vL��±w�^�3g��E���e������)F��_vO� ��Ni>k-ͬB�q��!R�H�q�7on�$��!�B�d��h�T0���:#�
	��X+��Ax�l��X�tP!�~�
�3&9F�m��JT	Qd-q��
ԺF���J'I#߄B�rAҰaCO$�aM�ϔ�O�:�2��/�aϞ=)o���߆���]�ΝM�M�6y[*�Rp�q�U_^�`A�}
N;�4	t!J���/3'2���l!F1��<�� )�BDYD�q�w?�z��A?������J���K��l���I�N�n�B$�P&q|�)��o�Y�a�9)rrT_�B�J��W=bG�$���k2�.�xX'�8	~�8���������"�����n�e=��J�!�MhwN��5�J�8��}�ᇵ��d�ɖsp`+�)���������SԌ=���ͳo}�[�q�FB$��o�%��'wnH
�]��з=p����A^�����{x92n�8O�糶`���%�$���=|z�����3�� �m۶��ƨ��Ъq�1�Ԛ�ޭ[�}�=z���{��B���5�c�dG6�͹��t;9<��Þ8O��z�M�0��8�B$��3g�I��Gq��}��=!Ά(g+�)\���!��$�?v�Xۼy�'���S��_;���#�p;�����|��^2�*�`%k�?]�,�4��$e�rGO�3%E�;�M+�BD	B���ˌ#p��Hdlٲźt�R}YO2��H��.kn2��tS��8Sf�B��%ҹ�!�A��H.Il-8D�B$�w���ʖ-[f¬S�N��z4K��di�C��!T�I(�׬]�v�ZG0 �ҳgOoKf�s����@2y?�ر�F�"yH�W=�P��N8��!�H�	�:^!�0���i.u�`̔si�;��3YEf������+u�80d�gϞmÇ�(�y~��o�K��_�֤W����6l��˗{-�)�1"�i"���E�L�l$�+�'�x|�������B#��ӵkW�bɒ%�?�)G�����:'d��e��&Z��� b^W/.�]�&M��ݻ{υ�nDe��ׯ��#ϸ57rM?�;T[�^��FF�`ԋ/���NP�Θd2쯿�����($Ѕ��`�֯_?ّ0J6�k��۷W_�a���QlN�K6;N�,z��r�< �/7m�+�m&�[�.���j!Di"�^���������`�!�H&k֬��|�3՗�ؑ��pF�;"�]�6�����֣{������W�+O&d���>O�x����$�E.L�<�	 ju���@�P���[ߌ�~�V�����ǋT�Er�v�N�q�g��G�Dq��<��+V������Ʌ����c����.��md�ٲM�qcb�(��r�@���k��+�����3��e�]V�vO=��:���~�{��S�������Ϯ�L �[n�u�X�V�̬�����+���ω'ڐ!C�/���� �`���5��qL��e˖՗�;�<�2e�	!D�����t'�3�U;(	v&q��㞉.D!�2�Y�f֨Q#/�B���f��}��/�(-$ЅBQ80mv��8e�p��N�{�}�Bą&z�1��t����P����B�j���rkܸI��S"��L$�Ծ}���=#���.��y7Zˣ����[XÆ��.u0������0�-���L1?�a�3g#s��}�\[x���֭[��=�u�N�:y�z���A]!D5��rJ�Y�٘<y�WJ��?��u�o�b>N�~�]����O��?��:}���ꓭE��&�-=��sc� d�ɢ�A߽{w�8�|�.#*99~��4G��5�����~�k�.�R�`���ý�&W�>�h��mڴi�D!Dr�@O �H����>"!�������4Ϧ�Zg�<�k�L��(A���3��[]��Cg.��%<(�nѢ�'@��e���g���;v�o�a;w�,�jFd�#����̞=ۄ�E=b8�;��/�r?��Ÿ��E�)���)���ٰ�M�d���L����{�S;�ql���g��c�ԩ^�(���k���r��� ]�t�6�k۷o�Ɩ!֓����cǎ5�c���'�@Љ�&�Q���	N`���~p�5*!D2�@OC]��B��9�6��a�EP\ ��~�@�d�%��UUU�'���ܚ�������Q�.8@�Ά<3��f�۶m[����L8��A(a�z�V��aÆy�	�Y]��R��������.Ŷ�g!���4j��VdA���{�1�HG�?�Ìf��>h�9��ጐ$;� u����i�n�:�ܔ���?e�6�޽{[�=�q�����Q�� 4gΜ��<�!B�3��Lu �_B��(��hfs=���t0���v������¬P�t'gz���˴�q�ۦ3fq����Da��T���ӳ�������7QX'��k~舶b�!�=����7n�a��`��U�Voǹ� %瘺�:"���Y6���A�<>�<����2D:��d���%g��"�ݻ~|��H6��\ĳ�4܉q���$�_��۲q��燾�k���۲1z����y�y�e�'�^�z��O�]��r�ك��/1/�7`1A�K��U0���޽��5'���M�l˖-^�<jXcR�����;w�:�,���M�ꫯz����Qg�q�����_B��Q��|PL������M���<��6s��H�R�_��5�_��0ʵ(kɁ�n�B�РA}o�1��x�|��U&r�����)�=p@.v���{��T��3�~�����h7f�ϟ`#��tw�K�|�ln�^�Ҍ���ŋmŊ�HG��ʪ�� �P_�h�w_ł����^��o
BDG}ʪr�0ѓ*�y�}�E�g��I1j��Lℒ5��K��J��O��?���1�uaܸq��A��^8(?�cRSH�-g���33D~]�2<�"J�q<����^@F���TB��*�֬Y�eԋ��"����!���	C˖-k�g˵u@/�{��iB!�B�2��֧�Y�d����F��{7��L9Q��unD:I+F��"L�P�N�>���ϟ{ �D�cРA^%�%]%�!O@�ɥ���R����7��~���~��Z�����mĈiO�Q!"�]�vM[f?��O�n�(E!�"�`4���ls2Ք�#��d�����8��<'��ݵk�z�!jm��1c�x%�a3�Q�m�6�ӧ�W��7T)�:ܴ	��unCI;�sw{m q>o!D��:t��aÆ���m�K/��Q�����.d�3���^����B�L(1Ng6��r�xJx4~V�j�*wxߏ;�f�m� 	[V�8'_��<W���`O6�¹s�z�b>h�G�K���e�b)ywA������l���k�!'���%J�(�Y��8��������VD�������B!
ʵ7<a-Zd_��|5=����̨蘃!f�t��11�5����G�����#G�t���:���G��/4��.�`����СCC�-�J���11�m���^6?��v�)��Ô�Gϓ��R�|�"�E��sm߾�	�tzv��y;���-	p�x��L!�($k׿a[���],��-K5�#�S\�@�B��b��yP�S��|�r�،h�k~��1��N���(�,��d~&�Ѽy�POx&�d�:���g�߷���Y�f�&�����)�;���J@�>{�|zvof�;i���-^�����C�EQ!��׿��~���Ȣ�=��H!����}����u2�n|>�O�%r�5-����A�S��g��5�,n������qSϥ���q�gV��YFP���#�l\�3gN�*�`�;�* (��uD9�U���e�l�<����߆[�c�Y��w�G6��6e��CQ:�G}�.��"+&eL�0��BQ:�iEpSbܢE�Z��G��N𲛜�|~�8Tk[���"΃�։�t�I��5��`��K�z��:<Z�=����TT �y��w���k2�.+N�ĉt�#��eJ��8�F��U�j;��g+_+�V�E�����N=�T� 퇃l�
eaD9�r��`���j�٨�ʀUB!D�à8"k�꜏HC��U'k���DA&�X�����W��v�~�����s0`�͛7����l��tf���[�߇�˜o�})l���4�Ф��]��N����%��z��}F����Y&*��	t�g���J����k�Gaʈ#j.\h�Ǐ7!�B�ÆK�G�Qv���NןKOq�@N��p�$~H�`��j,Y���?�Í��̥̝*
�@'P@�&S��A�\J��$�y�$���g�]BK��AU�߭�Q&*��	tX�r����?��n����4�0���k�U��BQ��gN_����)S�k׮^f�%��c^��L�U���ϗ.]j]�t�����L�0��E���H+���.IPM�>���x���Ae�H.�e����	
��ST�����;��N,"�Ҥ�}�{���B!J��1�Je�E��&����A7|��i�,=WR���\>'�bMIf�`A��
Ȓ�^�Ʌpw��T8,Z�ȫ �c服������O�͘��D�Pt����o�ٌd�6lX���D}�5���C!�
�J�����jq\��;$�����,9�"�	���<^:u�T���dɒ���kC:�g#(���R�y�-û�7ǎL��
���Ç�v��C5	��M��
��{�~�﷋�ˎ����ښ��ɿ��XF�d����/z��;���K��g�y�n��V-Ȅ"_|��2�'�bI�q�ָqv��m�_�c���&�!ݧO�׹Qc��|���b�ɚ���Z���O� ЪU���ON0 MV:N�9昼Ĺ���t�|���0y��xc��}z���({��m��-��ӫ�o�U���&1�1y�9��g�a��ַҺ�������W���FB�����,4�����K�'O�$��.��c��ޮC�5)$d9,8����1�c����=����,+z��U+K�f���x�y�9w䂛S���U�����kF?SI}�L<�ЧN���c|]�Ϟ*?Μ��f��$���&��Iz�(\�PO���d��&*�D	t�����{��\r��y晵Fy�a���K/����)@����/u�S��{�,�I޽{wϘ,�q
F�4��b�H�ܘ��h�Z�P���.�@�I��0d��p�#�.�ٶm����#���o�0B/W�"9�@A��M�RyD�Q����`�� ��fp<&.H��N�(�<���{��I��\'�p��n��{lĈ�F���D*�N��pf�;w��޺~�zB���'�t?D;�'��Lz����eT0�DA�Z�=I.�/ƨ�Z����G�	u�߸�*�o߾i�]?6��c/b�`oZł�,a��<�u&+۹s�}�A��E"4�%C�	>��w=]=[;���]����~X��A�g϶O���?�q�"7�>��2!�������#���
tB����'f�D9���Ȕ�"8c5��R�h��.� ���.��nXXg[���-Ƃ�!��X�R��(� 
Y�ѣG�]݃x�dk���fٗ�����9$'T8p�m���<�Te!y�v9�,\����<�ٹ���J?��h˔�S*�z��Q����e��{rY��1�lժ�w9W>!D�$^�����Js�0�f�
u[*,n��f�v�J�X���?g��;i�$���M�|ݖ+��[<���Y��n���s{�����,�� �(����c"��i �('�lډc��(k��ɱ<g�
<^]c��EdQ�'ݺu�`�Z1�@����2K��f$UA1� �ݻw�ϑV�`�z0ۜ	��,��|���������L�B�F�P!*20a�0�΢ɇR�q�ƙ�N�@aX6o�m;��gS������v�w>mW]�i�@����pCa��f�3!�~o2�.�e�s�~�ڃ✪!�%�	q�kq��l�?��w���[�.�i4�P����@Ɍ3�2s����0LI�e泥O:� b�����%��ʨΑK6�}��E���|�o�V�FcքH6�BT�dqr-�ɇV'`ٲe����0���K=�jHU6%|b?������N?����8�v��ի3�s?��ŋ{~6�0-�)%���#�)��$
��3V˵Zp<� �~t���>�T�s�W��/��a�y���W;�S�����B�瘫.� �=�s! �u��P�g���0�B���F�9�C�/΃ '�;�Äy�={���1}|�zH�ǣ\�u��q��.A�0��rb�F߰{����ׅ����z>���j��	�!�s9F�����gA�<�A䯲U��%O�w�B�{���o�87n��)���A��E]$Nr�r���'�r��@6���ϧ�.��>����Aq�lF	���\�մ�_rp1�`�|"o��LVX���\\�!8[;�2�`R��:·�V����8��.�j��ʘ1'��Q�D���EO'�o���p���Qo�sq(Gܧ�A��%��|�.�-ǃ���s^e�D�m~اy܆χ�7�=�3,�T !Dv$�E"��.
*�E3������r2QΆ�,�.��Ҵ������@g��*���~U�G��'��ϕ�@�=��l2�a��[���	�ɮ��.���xX����y\k����w�Ź�υ�r6�"b���@:�#@�X�" 
F��C�\������r_��梀��@���^�2q��%7�H6�BT(,���tQw�3�Qy{%�"4��qy�[6J�7kdW|c��p ��pRm	���D�1!b�_��1/�2_D��.������:(��*��:Yr~����-"983�At.ؚJ�A�K䣄�o���5���61$H�} �Y��@u�m��Nߓ`Ձ"yH�Q�yw�l,5#[���w����O�훚���|uf�Hf���Ƭq,�ؖ�
q�L�5k���F���g���8D �_Ȓ�-v ��/XM�h��y��dr��U�g�e�*0���gks���}g_,d�"$Ѕ�bW����sg���B����x��8�����Z�<Oh�a�ڐ!Cj�+a��ɸc��ׯ�o��e~��8p=�~�D~���z�P����TUU�t?<��`Z���D ����>��@EF�6m�����iϞ=^p���q�G!��B�	�`�SO��}���& ��i'���cr�6�iӦy�ܠ��%�d^Î������{�Ddج�!�t����4�	>G׫��$_S�~f��G����Sû\����
�d��x��l�?{�&E���2�������� 	�ΜN1g=�g�p�����!f0爘83��3�� A�A��ͯ�֚������<#���t�z�o*���!���!^D���ɥ_�~�����ϫ�{L	��{��[�"b�]w��D���V��AH�ڰaô@'2�p�6�NqF0���	QO$�\���b�!�{6�K�ӯ'�%��zs�yP3�$p�rC���R����rԨQՄ0��Q���� .j�AZ��~p�p���� ��4	3h2y�~C�b=�ɤ��瞺K*�U�dH��5z�h���o�����N�:�m0x������3���<xpࠏP�ܹ����#Gָ�2�;�s���3F	نe`
5���vnV�^�v�m}��՗K� �AZ��Z̼��jŀ؝5k�~���ǆ�y�������OwyM{|vk��'�ܵ���.�jC�����Ĩ�+.B�$*�/��Ru�ᇇ~?�A���o�]80�g�~���+�P�5�}�y睧�}���u�a�.��B�B��q�E������R7�p�g�̝v�I���W�ű���y�%B��dh�������(A0���Z�<�4��LVŹ��0�ĥ�A��E�q@&%�u��k߾}��v�$A=�lI/p��$!K$���.��� d�L�������֯[n�Eu��-������ܱc���8���������i�^��%��_|Q5n�8��3Q�|���裏Vg�}��_B���6�5�D|��󎁱��,�v� �q�L��F#.M�;�f�%���e�����8�V��^��"W����	Y��/א@M�\[�k�8/�a=g�>�ϣ�p��T2(������E�Bvɔ@���Kt}�؋��#F��Q!-��k�Ճ�_��W���n�Z:��	�t�G}Tw�y���D��	�ĉ��m��m�Q��4AHD$����@L�>�C��fk���@�a��F]�	�!E�_�Yn]��kfn���%��IB�����v��Ejh���ݏm��&�R��h:(B�&u��!~���W�L�ΑG�YsL�K��9%M�K��u~��Ԑ!C�@L�8���V{�9眣'��z����_x�Oq�`|�}���c��I���SN��\��o�Y�H�>` ��	�zV��5�)wc����
5�>}�(A��`}jZ�n�8�w�uW�ɝ(j������	6A���uR�ӊx�)�D���~`�4i�$rG�B`�5����:t��Ax�h7�5�Cy�m��w�s�vGwAj�tvW|�z�Z(�j�*��~�?H�ҥK���te�����l~�a�vο�:�=z��5�n*��[o�u�m �9䐼T��Nդ�_u�Uy�ǀ ]�8 h$�a���Wm����7տ'���x�	*n�jA�$@�����/j�M�5/��n;N+�ɾ��F�d� �ZgW���{��3�ͅ �f�X�l����7�����)6͞��AN�,\�Բ��9hӦ���H���*��΀b�44��H!Y2����O�uW��Mf4�s�[ٵk�j��@-8k�^v�ey���g��t3�T�/)�� ����j��A��A��>��7�|Se&���̈́	� � $i��@�1�#���ڑKއ�oР�v�!��Q�F�0�qA�c`?H��kx�pľ��n���o[6~�`l7��y!Ni�K� ���'v�� }��َһp�D죦�h��{������=�����p!��,M�ԁWp
ћ���PydB����Y�Ć��@*��I��ѽ{wu�T�z�y��WZ�^�
��Q;�
t �%�.� ���^������u�A�Q�O��-#�Y2,��Gv�1�5�B�g?���n��X@��I��#��y�1��L)B��r��oD&b���w�9��n�/���Ms8s�8֨�������R^�
8����A(?�tı�!|�1�xֈ{u@�c�=<�ׯ��k��N�~���{�6g���]�6�K�Ξ��0�-� Ba�n�E�Y�Ĺ�L"��;w��"8i�n��$j���%c�"��7��:۷������=�L��� ��t,/��5�A�(s1۱����.��c82�~��K(! ��%/B�H}4��9K�~�T�޽����$^�����\�΀��f[Ҩ\Ђң�m���;�:��<G�.�~��W�^�{�|뭷J��Fl���O?�����վ�7���$ �c8��]AH�)\�e�\1OD>i�mDup�췩�Nc��<�C�G�IM;/w��b!Z�#��漅@���//(m?8OdX�9��[��@��P9d&���GQ��~���IʗA�E¼��1#��ⰵDt�t!5G@TOrm����o�޻�Kzơ�� �l)U�s�4�xcuZ������w�|G�5�Q�h��3��"J"5���h;�]�m�R��ĵSD��b�����$`v���@GPS6@�?B��������k��ū�#7*Է�j�_�>�жmۢ"���~���qK'M_�$�4�]i�c帙�.I;	AH�L
�SO=U�Q�͠o��h%�D�U��~��6�L�~��{E�Br �1���d��T>͉��KN	�s�黩m�m\�}���oV�IF��to2�#&�b���m����dD.��UD��~"�ԛ��m�4�٭��ڳo�'ׁ�,6v"��6B�t��ŵ�sI:/9��G��ؙ��&_s�q^���Zf��O����sA�\ʲ���3"��mG���%5l���D̄���Ck��6��C��&�4&VA!���j��M��.T[��3����c5~�h��A���D���D9m'�����I�Pc�L1���T�B<�w#f���=^Q]�-J�@��X�"/m�+ha��m�������[kԨQ�"�,����ӫ~&;��x��t�9Ŷ���
���wf�:q�	Be��@�9��g���;�s�9G�+�0Ȝp�	:������sn���}^�ua^�`���˂�D�<��ɔ)SB�7J��PX/�P�[إc����r��.Vs�P9L�6Mn#�'�n9,f�IK� ���A��D��ԕ��4�Kc��`�W=8A�4�w���F�� ���d2s��B�ߤPf5y�d}o�����6���loj�;��m2��΄s��w�3�<SG�mX����y���V
��7M4lq��~���罇��Ͼ��k�ߏ��k��;�pp?�������NSB�!r���C��#t�+x�`��J�{���}�>]&�N�Y��6I�:T]�n��gl9�SPZ;�;Ｓ��A nq8h�w~�Ro^��)���v�������˹��� d�Lt�?���6Æ��[oy�)��[n�%p`fP����������U^ 4
	���:�3��;A���[Cf��֯�E��&����@d0�6o�\�0]�����4[��Mll��
S6g�pӅ<��v/�N��D���,Eϱ����2�p���n1M�8vĿ���l��$�{l��w���s�P��&��g�lD|˖-u�eU� d��t&XR�]\^�g�yF�x�y�Gx_x���[o��~<�w�q���z衼���\g�G�#������Rخ���j�g�}�'� B��g�}�!�Ml�q�n�p�����͞]����y�j���J��*i�t�nذ�.AC�9D��5���d��5�M�$���b_UDt�_l �� d���w9�L$R̹3B���k�;���,KS42+5
�<w�ر���={���6`�E�iR74�ZR͎�s��Y"�Kd;HQA�,2!�8�w����������w�qռ�={���t��o�>�g��ÇW���)Eh?���y�Ǩz��t��O?�WFZ��?^����G��?Y��C��{W�Hky+A�H�_o!�;�@2e�z�����6��IZ��zaU��DX��N�(���t�����E��H��P�6�����-R�N��j��ܸ�?I4&�W�n��ҢE%Be��@'%ͮ��+K'M{�M��}�V��LW^y��ѣG����ٗ_~���bA�#̽R�h�ƒn^�i���S'�|r����'�|Ro�����ҍկ��)�'���`Aj��	���Z����wT�kQB�ǿ�ڎ�Kc��0%w:Qd�r	A��=&JMVL�6mB�Ax�h̘1UN �)�A`[e�
�P��.Щj۶m���~�W<�����WG}܎�������n���>Z}��G�<u<���P��+&��;,T�w!���ڑ	�K�.�20^`��;������Ӑ���?8W_z�ķ3��J���_^���rX6<�/�AZ>k���܌��(�5���&zt���J[����s�Y�J���n�tJ�3v�qG߀�A�� �J&R�]0���~饗���I��I4;J��!E�H|D�<�@u�7��/�8RzԀt�=���~�i�Y&1{�a�*��U��K�y��ف�5�� �ܕ�d =#����4K�0��r�h��u��R��.4�-T�'d��qW����)͈`R�I�6�Ҁ�e^��;��H7��b�& �$�z^���2�.�;z�Ң�6,�ÁF�ƫ��%̒�����:8z�XN��Rɤ��h�'T.q6�L�:c0	3�ѐ��1�|
u�tt�O�>�.P]�v���N�B����ޫ���:�C�+����֭��~�Q�g��;Ｃ�¶��W�~΃}.�Y/IO� ��1wȐ!J(?�tm������*M����9�ȑ#S]��98�S[ �8Hj^'jM��W�%��NhժU���l�^R�L��؁I-�����gdwq�^Ď*�aI7**�D�I'��Ҁ��k��/<�4��s��FD��O�^R��u#q���o2Qu��lC)uGt"�k�s�y(u��t�P��W$�X0��P�����ϝ;wV�{�����2���������+���vvu�;(�f��\�8�A������X�AR�M��1�D�a��� a�-Gj=6U�.���m�]�w!�γI���(��EY�f��Uf,���	��N-�-7���#P�&}���*�e�lP��X�ک�!�6�_.�yeI��'By9��s�5�,�������gv����t��hؠ�j�|3�ݶ��l����J��paA��'5�D�"׆(8"��4��L�8� o8���a�� �KLP�=e�ű_�q��@@������l�Y��|��B��&x���dϋ�s1��dp��(���������f.�97i�f���,�_W]uI�M��U��ᇟ���MQ��VB��	t����n�uGd4hР�簓�~�.]B�W&��C��B���R���)�Y���5YHY�V���n9V�޹�����U�4�D9�z�6���4�.i�v�Ӆ��l�zr�'kn¤��كv7w2]��!�d7�ddH?��	Ĺ}mh6��s�f	�P������sXm�UԹ��V-WS���� T>"�k8�H'=�����f���n�ܗBu�*�A"�%9��}����6�$�ܫt��a�d�oZ���x�9m�fo�f��M6M����hXp��nn2���\��8\��B�ԣ��`_2�ԝ�Y�=I����k��q	gϤI�B}� �|���f�A�0;��D5k❩�%?��"�k"�Aj1[�����꽽z�RS�NUiA]�����ʀ�o֤&[˫�9"�h9��r���,��}l�8��Y����ei
t))�d�P���D���{��߾}��N:zU$�����8�q���nU?㌰;�������t�� ����7LD� T���&mi@$0�@����o��҂(��ʁ{�k��=MO�B��i����}������7}BR�bG�Ӫ?�����4K@!��EOj91����Q�馛&�9���]֕mu��!�Һ\K��{R���QF���^��܂� ��⫥�}���:�e���#�����[n��{����O)A!���z4'*���US��5�����v�8"k��ֿ���Qϼ�0�_ޏ����I�� X��j��<K��QsM� �h^8]8�$KL8�'N��	@x�N�"9X%(��sS� ^k�s��5b��w�����B�9f��fŏj�5�C�F�߀P("�A�*��c�؛�!F�~�钾����N;M�Ͱa��{ｧ���?��~����@p B���"*h�������:#Ĉz	��A��k�#)�H"�:L�=	���9`�iF��S�³ۤI��8�e
��4�=P�@������.�`Z��j�2)������gd���l�����ԥ��VY%�y�����3�P{�.d&�Gy$�{_}�Uշo_%d�]�����������Z�x@�߹`��X�)�Ŀ<ܒ%�S�B� �h���,�e:�ч�7/ޏ�D����_>N�"���g"��dʔ):�܈@��QNPh5�M���>p-�,���K޲v� �(|Z��۫���w����q�M��Zv!;�@}��;�������?�wG/P���~�)��J�"Ѕ�����>��z�~��l��Ð"l�� ��
[\Q6��f�/^vgw��&U!֨Q#�"{"��:���$aɴ(ZD ����=gB4ACܒ����ڵSC�M�AZ�p�q{]o�!:v��+<�����^�{9?��u������M>�����c�P��E��Q��+x�jC}�WGY/p%z#1��oFmmb�����_��j<�`�Bjٲe�+��/�H:�pl&���_8���p6 ��D��L��֦,
�a�����݁�6M��8q�����ħ�Ԝ}s� �i�?N'�-Z�T~��r
��j�Y	p���w�?M�@g�Ȱ�RIs���TM�	�?��O������ �C�ƍUmc���F��2�M,i�ʭ����Q)fɳR����J��'r̒]�QBs2�@ҽ��A��I�8����EFC؀����r�`g��LJ�ܹs��#H�F����2A��\;�.d�J���w!s0��v�m��;j�(%d��~XpAP?Z*��Ν3G�Ԝ>��#��9r���WY�#�R�w���ﾫ�z�Y�� �| qf�� �8:ޱc�j�h�-�Y�"���t�����o��.8fH��b�-"?�K�D�M�=�AҬY�j����	�^%ddg��]D������bB� �5��Q������$m]4n�0�]�Dڸ�Q'�ĭ�;�K�⡖���I�6�e�b���,Qd"ۤ�S��m۶-*�q>f̘�9 ��Y��{8��8�u�mHoO�� ��@g@;�E��D
-ua#� � Ɲ/�n���Z%`�8�ˀ��Y�:-���~�v���:�@$�-�h^G���[nY��M7�T�H;+��%=;��>��,?�����.kܸ�^v/jJ;�Ĝ��.'����N;K	�@�{u���ܔk�>A��ZƫݣG%���^�z�z/�`�AA��m�F�5Ĉo]��KM5���i�-;��c �lCğ�n�^�����3:��9 ��6t:����vە���4v^aJ�'Z�lY���*ӦM�D}=!��jڴ��1G�sSSN�#j��O�<x��j��I�'� ����� H�� �  m���JD���,="ӝ:uҢ��A��战4�Q`��O�9�"�Q�_�
�A"�8G~�&M����NV����a�� �>�����
%��'"�4�+&[�h3�,�Ã^d�9�H�G��Py�@��0Y���l�߻|�7JA�ab��o߾��{'D���r1�ԓ���v:2��^p\�(Ёsij�	g�!iڈ^�5��8c8'Ժ�o�e���rV*6Z� ǃ_����K���tD��R�?�MÆc��C=4����#�L�.�ӟ
�DU�#� � =�cǎ�QR����R��rI��}~�[���(�2e��Ҙ�:ug���7�5��81�-��a�Z�sw9����@�5���Ȓq� �>j�@g�f�f���J�)@��ׯ/�+ ��=���w�u�����[aA�,:���c�6ѓY�f�����L���C܍7Y7�4�8�kh����oTq���h�%��,sEM��:�s���\"�;�C^�E���I�>�a���T�h���q,�I6W��w����Ym�Fƈ�x����9q{/�U�!Bq���Ǔ��4)�sJݙL��0�~����	B��:�֫��w���>��������������	�<L��-zK5h��*�O�qf�G�"@L�pR�M�7��������!u9M�
(��+m�~Fj�j7��9"c�&h4(:�bj����z:;�n���gG�Y���d����ؽ�ya>'By��Y�	�_�~ړ~���ə�x�M��6�s<��px�i&4��{�N�� �H�|����[w�L�s�p\�`���W����B��&��)g�s7R���������.�^��
�eݰ�2(�B�6`�v5�+==(�����_�i�F�L�p֚�	��)Љ�<��S�W^ѓ/]6�=�1!v��Ew�qzy*^�_~�G;DC�lC��!��Nl���m�:ut�h�#'�K��:�Wk)B�`�  M�1Q��w�]�,��%�6�püϘ�v����j�4���ID�k4@D��=:P�c߶hѢ�܈�D�Bv�8�Nt�gϞzpe�!M�Զ�_~9��00���G�hbu�e�i�N�P�kt
��DڡC%��8∲n?��s���*!s&�ĩ(�&��G���~"�mG!vC��ी��NM�Nڬ��P��#{}y��t��Ӻ�i��g�w�"ݯl�y��|�LP)� �d�N􉨵i�¤㵤I����#�hc�eV������[oia~��W�z�#F�	4	×�e��?>ۭT��Pc�6g�����oR��\
����jպ��ߧO�&�B�a�=���tu��a!�U��d���N�i���mf5"�~K�	����(G�3�ז�Bf)A "�H7��y�lٲ�����	��=J�4a"�ݫW/������sO7�^xA�r������W^y��O:�$��K/隰�����5�
L�A��ڮ�����Q�F����t�'MV�P[i޼��G)ufDɜ3�k�/Kk�a�P����}�>�ƍ��D;Y����9�� �+;�SU�z��۵k�E�Wf�-��
p	��y�s�]v��VE�G���ץ@:����I��v�w� ����;u�˸�6,<Ǉ~�A���Δ�!L�:Sc����L<j�Ӏ  Ml	j� ��>��ǉ������Be�}C�'v���(D��)��kvI�/��� d�<�N�5�(��dX���%-���n�A{��@�v�a�m�tӌ
�NAA��w��v�u�~MI��!����"����8�Q.��t��I�;� �g؊��=�#�Y/���N��đnN:8��8��5�4�����>P_��;*AA�g�pMT��W�;w֑t����8��Z*�L��X0A3�x�f�|?#Y��m2-�I���M�yڝ�������e���w�މg����3gN���}�ݪ{��J�.�u�α~<X�|�ɱo�%�&L����}���g9tI.Q'Y��4��D��f�;��:uR~��~ٵ�[o�u�*-��+�pH���Hz�������X� ���
t�Ԩ��#^.aL:]����[׮]��<����
��-��e��w3Fâ�ե�\�*�w��_� x3}�t��N�r^��m�喺+:Qv���29)jԤ>\/��:�x����@A�%[�-[�ԓ��F^L=��<�6�˽V#)pD�hRw�A������6m�T����E)� %A�-�qb�i�oD�d�!�Ӡu��U�d��-\�0��pVӼ�|�����j'��N�&2J��MTx�%��vA�>%��?^��5j�H���￯'"��i��{��mȐ!j�}�-黨�;�쳫~/� � ���ŋuI"��~ V&M���i@gm�vLf^X��~�bw  "�����~K��Ί����B�!���.B�d2�}РAZ�ge�p��D��~���P&���B��!U(󤶯g+B< DH�eI)�F�s� @��9��AN��C������~B^��9����u��%��xp 0�M�VU�.$�رc�P3`A�8�i��(?�c޼y��-AGkl�M�E�n���q<"�Aj6��L���5�@'�AM� � �5k*k��7߼*"�*"�o	9A�f�9�βfPh���1���?� � D�F��A���	t:�BR�.)u����� فN�]t��l�͔���޽{��S�*AA!�dK� ����ԟ۰_�Z&�����U�&M����G��5k�;\� � �&s�&.n�UV@�G�)Br4m�T�y�ׯ�:t�^{�5%Bya��R֡D��9�t[�"YX�]�?Ȫ3/kd�dHj+d�}��GJA�Ȝ�V�n]�Via���6� �0@}��ת�ByP׮]� � �PydN���I1��:t�k���W� d�nݺ�iӦ��
KBJ� � Be�9�n:1���O�Zj���馛*AA�0L�4�*�l�2%� AdN���O?��c�:�ҐJA��,Z�H	� BX2'з�b�����N���Z*+|����I܎;�A��:�(ժU���3f����Uh�r��=/X��gϛ�P����o�~�S�N��XA���6�A(��	tD0K����P�B�fj��-Z�P묳��2�a���^{������jf&�SN9����~��������~�~�={�jk����|��u���p�|��g:��湂 ��;_��� K�:�瞺3���k�]������=��C	� B2D]~��U?�F�}'���b�-�Tm���2 &O�\��d�y5�%��o�Q�ƍSK�.U� dk-[����f�2e��b)Y����WM�8�*�cǎ:�\
�o��jܸ��;w���r�?��X�^�X:���^{��g�u^G  Z~IDATRX/��b%� 6̭cƌQ;Ｓ���#�8B7#:��r!��M�V��,\�Pm��U���{�A��:u��� b�UWՑslv�,���YJ�d�>~�x��{�U���V[�,��c�Qݻw�⸜Qt"?���:��cu
Z��>�ȑ#�~nР�J��?I�r=�t����^z�J�!�v�e%T��8��mڴ��O�)�a�J��ڵk�'�A�<�O>���R�d�;t��I���1F�J&M�Diذ�������2c�%�PӘ>}�:��3�=�ܣ3�����r�m���8��>K� !���r�Q	����]w��	B)dV�ù瞫.��Bݡx�6H=՝z/&���?_&DA�,<X����ꫯV��g���Ml�c�1ԩ���qml�/����{�b�B��qFﬧ�zJ��T2-�7�tS-�o��V-��ׯ��H�����裏V�Z�R5<�{�{��[���8��������A�i�؅H���G������w^s�5ڰ6<���������_~YgSԞzq���-�w�7�Xj�0�mXr��
��.�@�;V	��[�Hq�Y�&�l�V_}u%d2�<�@��̻��v[Um�;�P�_��=���w��nj�m���?|�p�!#�,�/�q�	B\�	t��Q=?I7���;��ftD��I�|�r]�N������L}T��R�P��7�{�V��z뭧{(���8�����a��N�^Щ��^ݺu}�3��������e���A(DS_}�U%T8R�@���O�?�ߌ@g���*��qn�x@	��p��ĊU���'Ї��7o�x�M�N8��z�W��E'�$R��n"�l�m۶�[�n������\!)p���~�~�7߬�����3�8]����� $]�?��c���[�����ү_?5z�h9�9J'��.�L�����/����Qz�G�Ν;W}߼y� �b���J�������WEc���i�g�u��p>���A@��K�
�x�IQ�{��y睧����t������A� YJ��t\,X����@�ǽ_�Zゐ$d ^q���i w�W��N:I�1��LA��⅍����c�!Dى�� 5��:��t%�4�в^�-�ܢ'0�KW�R:��bN�8�l?���� ��>W��QAj./����+칟�&^^��@l���Z�&� d�L7��u�ֺ�Ͷ���S�h�C*��i"�g����r<҈t��O?���:\AA�R�W�%�\�z��YUsD>v� �P�8�k���:�s�a����y]�H��FX������p&I�9���?�c;v�5^�� � B��x�ҹ�]���N;Mww�'�|����+���� �P�H�n�x���G�f+&LPS�L�MW�&2�+��~{�tTI�A�J�Wϣ�ᇴT�д��Պo��j�js�r߳K�N�[�;�)\��ʳg��Zn^�v>�|�ک�M����V����J��U/�6�������Z�������i���멟~YG����9��U6~U+���Ze�oU�U���MU�w���0���=ե�J�#�V��.���9���y����8�A5r����ԩ���=�ڒ��j���Y�)�����N>�}I�j��M��ςW�i�d#5��J�N������P�}O=x�ڽs����Q5iu]���Gs��'�R����SO�-�d�/V��X_��|��tH���;�N�_W�J��SV�G�R�P*-�Ԣw��E����E��Z-��Dʉ��^s�5� � By�U������}*QsA�ZH��.Ԣ7j�H	Bh�Ǫ�e3>�쳼�5�Y�dI�{Y)�����d���|���>��.�t���;�`���qr	� � ��.5R�B1�{��U�3�8#�w^s�5�U�8 �wR�Q��k׮]�����RAAA(� �P�3o���w��>U�׭��?��:h��c���?��}j�zm�4���?���6R�u��:kľ�)�-P�<4\�����&�3N�Euj�U�ۡ�����!�>R,�����٧�V_=~3i�3�C��T�>�Zm�x#���;���8��,�r���;~�Zc�:�vP'��Zy�«݄��eߩ;��F���V[mUu�>۩�N�VYee7��9M�,s\-�5T;gw�Ֆ��&��`�R}޸���[CuXkuğ[Ǿ��zv����d��?�6��P��Em��ڱokƇ����ꃏ>S6��N=��ڳK�ط��?�{����':wj��?��Z��j�ok��9��G�U����sr�Q�7�};˖�W���?Vu�p�����ժ����Az-�t�nݺ���s��Q� B�|8�su�1�i�d<�Cu�E{����mQq����5I?�5����\�"�fK'��6��4`��ꎛ�,�I��?���9�5v�ܪߍɉZ�z��OՍ����%�x�����l45{��ST�v[ŶD��Gݫ�6�Xj�<�����&p�{o?&Բ�aq��M�2_��~O���m�#~���2w��S_,��t�ʴ�Jn��r�5/�5I�0����i��s�`��O̝�#OzP;o�@7��a?��:����;�gV�n��y���8��g��u�Ķ-���\�v c���:A;��b����a�=��pF�=[=��X�]�`#��B��#� �P����^�熛���o;����ߜ����w�;�R����X����U��Ĺ�_~UW��em���x�w�Ĺ��ȓ�ԙ���v/�F��߯Vk����?�nW�SC^� ��3��mqnx�I��wT��ټ�m����<qn@8���T��8�x�bu�m����&�="=.�>�87��л��wP�KXi�f؈Y���/X�n�9@���X�ý����Ĺ����_W�j� g��ύ���Pw?8L]r���lg�7�]w#�������7/�-������sC�����V��$��&��/�z�Fm�v�m7U�aM���~;�{�C� $K.F��Xo��9c���w�q`���E�=��7߬�$�q�f����*n��'V
��0b��0A]y龱l#܏g_�����Ē�I�r�'_z�G�+oLU'��FO?�L}��@G�".�0�p׎�K��!��[�@G�}a���9oq	t�_���8	XʬTX��Ȳ�aS\��g���v�5���Z�����%0���_���ЋΏ����&�����]^,��k���%og�3�8c�t!)b�8�����m�٦�t���=i.�v�I'�:�����K[_TJ�W���U�4�,�e<Ϫh���oU%�l�2�bŊ���&�6���ӎa?ƌ���ꫯ�7+�WkX�l�j�9zFn[_y��]���b�x�?��,h��3j��ف�?��<���
�w�D���3}�H��.�Q|;͝��-�;�M�������	t�I��~̚�����S�Ǩ1�E(vKж�g�_��s��Ĩ�~��_�x�cw���>7y�<���漹��L�6_-^�D�1f�G�~��,_~�:��믫m�A�>~4�3պ�U?s���;vsO}n�D���C��}���k�c÷�z;��Υ_��]�n���>Gd|�L�4'�s&���|>�vܱyᢥj����1���r^�lK
!)�;L	� ����2i����8w�45�y1)'v�=-�w�s�1�4��>�*�sD�f}�H��ǋ/�W�v�CX|���P��Qcf����w?�ܨ1��ے/�	��9s?��܂�_t�<��ؼ��y�|j[���P���#̸Y��<t�j޴A���M_j;3>\�wL�&�	�܇3��i�.��󥁟�h梼m f��?g�w�7��eS,��˂���+W�W�߃>7୩y���0�m�O�5��?7uڼj��t���Z�di�����k�� {�	��˪~~F�{a��ٹ���|rO}n��Yy���?��΂���>��^�$�Q���1j�FV�<{n��hػ��gU?��a�熍� �o,�<{���3s֧y����?7?��W�OV�[N����T�#Y�"�k(x3y�٤�T\/� $�:묣�[o=U[Y}�hi�mڴQPi��*�n]���K.Qi��V[�J��ͯ�WX>������e�g,���K�꫊�o�>���G~T�12]��p����b8�h�;���_Qy���
��9ڹ�I�+,�t�UE�T��������WT�{�~��Ͽ.ꞛ;oI�����S���k���~����1�"=��������r��WT^|y�~E��#oW���t�95j��P�N��o��i;[l��*'��M�0A�Ya��膇 De���J�l����?�,��N;)AA��D,!�K��{�n���[�{W�{ｧ.��2%By�+�:N��v2kY?Y<W� � �l$Ž3s�Lu��w*YD�����`�~���s�9'3Bx��j��Ѻ	�믿�<�@�8W� � i"]��e�������Wg��:�5�7�|3/����j�}�Q���kĳ�t��<�<��;Y?g�u�j޼�5�K���N�'�xB	� � ��tA*��w�u��h�����i |ǌSm����~[���;n�5zc)AA���tA*�ɓ�wlAA��!]��: �K-_��,ۧ�w�u�ͫ��B����wHMu�c��V+�����믕�]X�%���Wj�UW]U�oŎSB�0�s=L�G���K��ra�M�k7[�6�y�[�n��Ra\k����<p?���jE퇹�m�q�.]����3��F("Ѕ��C��/���w뭷�
�X�B-Z�H�7N�&Sk`)�����o��V//dl?��3�I�&U?w��M2Dׅ^�ڷo���v[�T�]�}���Z��SO�'�|R׳������SOU�;w��ov�ɚ�~#G�T����z���:���y��1��������[���U?}��j֬YU?�͚5��;ǰd������4kd/^�X��NS�w���a8q]�L���������"]�}7��7޸�oӧOW'�t��gIw�����{�Ua��_��N?����q]�ߘ�itƱqo��A���cնm[��&�h�
������{���W��~t��I�y�y�c��`�\o��t�#¯��/N&üy���^Ծ�w�q��|��j�ԩ�Y�4iR��y�}�Q��v�U�����/�7�P���U��G���g�}�U{~Vc4h�� �������.\X�9ל�b`�4���g���K�������e˖ꡇ���g�Ơ܏��o������nj��7����8ó����}�F�%�x�l븟���NӦMӵ�<�A�����yu���={�g�Õ���Ξ=[��A�y^O�a���]�vUs<��s��o��,�k׮z���5l�P;�9��|��q�-���ۅ�q��k|}�wԌ3�!h|e�:�S?�<t�%�膎�l��>.��fn��65lذj�a|����!ǀӋ���Y���o^ :x6��<���&���{�9���rD����0��}l���F?��k����7s?1wr����b���W�_}��<'��<3.������,�{�y�W��^!�������|2ql��.E���K/�sd�x�g�%f/��u��'W���ɽo�k�����?�-�u�\0f06���+����v�7����1��ls^����믿�:���8ٱcG�馛���[O���9�9��/����Y�]3Ot��Eߋ<[Ks/2Oq��<g����~�=���|~��z\�y�X��l�ͪ�
�i���
<_�í}������_���e��x� '}~X�c�����.T$�4�raPjܸ�~u�Qz ������̙��V�ZU����O1�3��� a�vЃ�^Wa^��1��=��*��!��㏫����s��LR���<���n�����\��iӦy﵍hѢ�jݺ�*���z�����D���7�`�l����+!q�����&�0�ɾ��L�L�.�38v����x�E�4�︢A|w�k��̵�3B]X��]G��Q��)���<׽{����9O�{�wh'�12�i�~������ 3���G2��Q�0��k�3��2め��=�.T�=��~�?��t���X��h?����?�8��ׅ�ϲ�8ƣ���߰���j'�� �AX��.��b�	���8-.��"��Ѕ�1��H>�3<��s���O�*�\�_y���%��N,/���
��G�q��q�ת뮻.��<�a������?��ꎁ�8�� z��;�B�}u�{�ˠe�(A�g��F��w���9m����mp��=�����w�8���ް�j���|ÿ68Mq���xn@<;6�x��3	Qn@���Z��n��&=�{߾�K�bn� [�ˋ{���ϯvp��=����{�ˁ<�8�x�Lv�ay�L�~v׍1��"s$���`�c@��L{ݻg�}���`�fۼ�7���g���kႣ��!�e��B��@*�#��F<��@�W�(���7�|s��O8�_���l�>�^n��D\�Ν�EFF��	�h/�6 �a�-���-}<�� ���`"�#�C"	p
`l�ae�f�.<�x�97nF@%�x�k���`cB'��b�	�CCgN��������?m ������\c�!��n�cǎ��5�\���B�"ƍa���v���]~ 0�Pb�!/�/8��L{g1���θe;%1�lq�=��%���"�9;�g Q�$���i���`��+TVa�=���A��6(jd[�#8x�>��#��1��`�oŤ��\0V�\`��%&����9"�̿�r�v"����_��y�駋���^�z����`��N������,la23���x"��b�Ȩqr �p���\l#�[����/�8�Ɇ-Bf��#����?�����p�]w�:���q����\2q�Ī��m��m�1� �|��2�p�o�����L�N7��j�e4Qh��a���V4p��6d>0Y�@�s�.��R�10�a�C�9���[\��^��,�>�i/��ľî�؍w��x&����u�NNn�E�9��BqA-���V��S�e�ź<��?7���B���J��]'C*'�B0�䍡�dI��L|L�n���0�A��D(1N�Z#xR��x�(��-Ι������I�Ў�/0�2�X0��<#5�uv��I��%,��hR�0$0܈0���&?(&�+�8�`!�L���9�Kc�����d�ͱ �86���؈``�r��( �
ƉuL��7�R��r+�/#�Ah&s�"`��~������{q6�=nxf��`pp?"��(b�]��+cs|�X�<w6D�2�4�d�Dp���ꪼ� 2�v�.�h����-�Ə�)�M��5��,�k��ۆ"�C�%]!�u�XyM�6�&��.# �s��*"Φ���#��l�@$��_�8��~�3�Mv@����y$Rǘ�<`G�p�"����G׀q�B��=�p��#ɸ1��A�/Ay�H��ϲ8 ��W�!7��gڌ��S7���9��x��@1������5Z��8�8v��GF�s>�/��q�y�g�̊��=#`��5��P(�u�<C�%DZ��3w�n�h����f&K��/� � �ñ�d/p���Ic7"�q�{��Ɯc;'d$�}�(�m�e�8A���S��!�H�)�yv�: ��䭷��i��K�Is/qo1�e�q~��P���d/G�'M�9�u�36brL*:�����a`�u:c/6��	^0�2��U�-��a�5�s�O�
lG�&P��2�0���,��}�5161s����ݻw�ך�A�kF)����}�Xm:u~}�{1������Pфx�Љ�L���^���2J:'k�܋B�)9����ͽM���^ܙ���	�ŭ�2 
Ic�87��<D�����!�z��m���n�m!�x�0pb`��go�c����c����A3�#
łw��&����:/�F&� /���L���Ƥ��75^��ӭ�����baܺ�8@����1���LM*cF�0���Z63�کv���б�㏲�)Cz$�<F���DoH[��A��!��j�^��c�8�����Xγi��wSf�<F����u��|�=>�׊q���&`����yLݠ1�1j������&��:��d�`�Ï��Z�"������1�6��('�kTgz�$	�<{_hD��p��Ӄ1LA;ͷ�3Ͻl@4!��{�Py��}<�8��L��&�9`ײ{���ᖲ �8R�f��i���!�책�krv6�-�-F<��<���!D���g��<��ݝ��g�qD0�ѷ�c��g� i��k��`��3V�w�6|����a���P�/�^���-�����	�7���3Y��~�����J���ۊ��+p.�ӌC��9{�k�˸���̳�v(_2=p�q�]��8D�m�1���1�y����w���`����G�@�qc�Q�1�����c��f`csS�#p�ٙ,^v�WD���bt�A�>,\��s/�I'�/#u���y�|�{q����[We�,	t�Yt�O�D�P%��<�;��E�z�4�:@�&����yf0q�	7��u�[�� ��6F���"�Ů8wa�m��E&m�'b�׻X8^�i�0`Ȇ�^p-01�["�Nq��B<2�a�0�s~��N����];L<��T��� {��&	��cֈ?"Bv��2����#)��B��k8�܉� �ϝ����6@:~׊�q`�)�$�X��`�u���A�}�q�"����`��'q���S��(�9GƏ_�-)�8�l¸��![L7�(�?��jG�q��<D��iFƹ�#��/p!p1��9��ܫn�k1� ��u��(���ט�c��D�:�z/�! *l��Գ�i�gt?�c(��_&�n�D�����'�mg�M������s<Hp��os�p|�ı��̻v�*͘�:5��t��A��R��87�/�v�0s��Lv�-�C����a�]�P̽HA��{��ʜW�E���d�ؐ�Z�L8و�r�'r�Mѡ��g�W�&�ܽ��F��K��� Y�ss/F��N�3��$ݡ[�\����7\�͔P#@�! ��Hgr7�3�>��n�IK7Q\&>kғ�\lA�����2�b a`�Ej�� M��[R�l�>���f�x���s���}>�s�]F#O�Q�$!���l�P��q�{I"J8/l�c�#M~�Ѹ�M��!E�!�=����4�����0B=0��^~��h������k���Y�1j.���Cq�L�����9�Wt���8纗R��#+���$�O�{=�'�B�-IFp�&otR�Iۥ^�T8e��Tl�Ydg!jLd�("~"�d\0��5�<�qt�}��϶('�h��%*7Nt#�?�4�D�ӄ���J���u�Ǚ�}`j�Sm'ύת�۹���-;sW#�k
X
\{�
�l�'�d�p�ص�d߸㰻�~McA*8� ����dzv&&mv���r��v$����ch� D�+���6�o;ӤP���A�s���ۯ���=K��}5�����܋�����@9:O#Vg�N��7����_��O���܋\���P��!���0� 2�5�ň1��)�@���L2�ۀA�t^F"sԗ��.�6������&�l�+F��ί����x�upp<��b:6�!�芒fY*�'�5l��H�cҴ�y�y�{�1��I�F�-��kCڛ1<0.1���h+]��dZ������B$�TJ��v-4�H��m�q�K��Z�䚷���D"&��&?xv�+�#��$׏枲Ũ�;=E�p�)�q�s�@���5���7�Tz]nc>R���*&zn0�+�!��, ����Y��d:�u��m'P��f���-\�i����D��8��>�X�����~`�v��Sܮ���z9�ߙ�D�0�uW'�9"��ˡ��WvL���c�0s2�D8�8����@�0&j�[~K�{��0[��y&s�r	:�1�Pfg�p1.�Yn7��P�w�INR���;��]�#r�r�i���*���\�̝��T��IN�q��O:í귦B�בȲ�x������n�v�9\XhXC�,��z,��k40��ua��@ېFEM��ZMt8�u���;k1��^�~�Q���J��m�6�t�0^�(�)`�����i&s���I�� ��m�?�+c��	ᷮj�Pl7�3���#�#��5��Z:�k�� H�F ����H�U][|��G�tK��=�S�jq� �E$�̽���3kGeqz���q��b�8�&�u�s;ۆd� z�eDR�+)D�L��L�W�C�	]
Ac�Dmq`�{��.7J{�r�?R��d.x	T΁_3.{��~����ĉ���e��)��5�ǹ�Q�'� ȴ4�X�/l�0�P�1�/�����X��8}K̜�5���-�$(9@�'���L'�#s����(E����9��t" ��^�x�(�@�5zl��㵊#���빓OkhB��Hmz�Z�xG��`t"lL#�x&HjOm��a�1�(:R��F��-@�UP::�&��@��������10� �^��r]h�ը`��P��?P:uƅ-j��G��+�:AҴ��-��T�m�&Lbq�(�F��Ƞ礱Q�]J�T���f7�[����Y��8!�������+��KQۉ#����-[�	�?�}�v�#9W�)�Na�0g�mq�~9���L
wq�G/#�(Qe��uK���čN�56Q���g��X� Pr��E䍒-�
�T,�W�{��:jz�6��ˬ��<k�;Ϲ5�a�2�r�H=�9t�Z+��vɄ8=�n���4�r#���^+h�c^R=�n�}�^f�Eܹc�[�f���J�!��d���8I��J��^܋��G�e��{�1�`4�#hcCD���V�!���R0S>e�˱����L�0p��Ix��^�N@c�es�"i
t�P����t�];|�������s�x�xB�������`jM�0I��	c�^�٤�]7Ig2��4�.�z�Oj��4`��N�#��^���>�����>�}�h5�6�Jq�Wn�0��*�6�]��"��8[�`v�b���;�z�@2q�bmwS�a�G�h�`����`���L ��}��"�&���PJwp�)N�D������,j���O�=��- �gH��8?\a<ktNO!�NG�����Y#���t۩���sXdEm�TD���}����2Y� ����a�Bd/���q�)��&�c��2'�m����Wc���q��<sl��m�������S�j�O �������FcD:MI�#��id��p�6�����&s�^Y|��k�y��L
�7S�mlf�S�]\��ǌ�b��������[���b���N�w�?��[�cV7���c�q�-��ݬO���kR�9�)�$�5�^��c�i�<��҄q���j�xR�M��s�SR����=TF���]�s�`ƍ���:i
tZ4�;�*C���܉?\����fvM<!x:m��'P?j2"nZa1��QC*���&�@F蒂k�e�]2L1d�"��¤`��AT�0�Xg�%� ��oi�F!�l8�c���Q�.��0bm#������8��;8?^��x׃� �@3%D�J�7���:��2"�:<R��z	���k���6���c6M]��a c�f�}J�[>�A��0� Q��'�k�Κ�Rh���Rrc�E�QJp\�ORM�p*����_\�G[4sn��;��`��6���C5L�H���Dn9�ꨐ�E�U��ōt��̽n��	�w�?���|���^`���g2NC��NΣ�ZY̛F8!p�hHg��h�D�<�m��c�����k�H�N�8�9g�1"�8��pv����y�v���m��%l�_�m's���$�|��O��x�]�	;�^�ͼ�{�θ@��q�$c��v�&� ��M~Yn�xBe��>��.����*��cr���&��P�N<�
��^tm�t����h�߀M����b �3j�&J{��q#�gj̼�Ew��DK�f�����L,{R-R�p8����ذ0q�*���S�8{]��p܈""��2t|_\�|���[��}���Ǒ�N�����Kj�]��A��emS�ԦF����&8�0N���Rja�H7�ߎ(!���k�Ltܮ%�pD��C����
ҽ���0���Sb�DY6��?��lÌ� ��4�c�2�8���&8 �w��'��c�{��%�o7#cq��r����޸KRpH��N�yc��-{<��಍w�20�2'1��5Υ��{���j7
�*-��A�
��t��!��]�g�{�8o|���Ku�!�Q&�~8�2��l���%a0eCo���A7���>�\�Cc�HN1�'<�v�*��p<����1�o;�qF؂��7���6P���N�����ΠĮ-X��-�#��I�����a�b�3תԠ�?�4��ћg�O�'�#Lv� {�o8=UXRԫ6����Z��]����,�s�rs�)��e��IC�3�"Η��H�z�{uTBf����fҤI:�O,�"�	�b�&hi"ۮ����h^ͥ�(9*�=�I�A�ҭc�t1��<c4�ҏpi0b�Q�xH�,&����J��m�fY����m�t�g��J�&�5�14M��� �m���j��DT1f0�x�	�.�+�	��)�/���&?&w�$7���-��id^$�&e�ԇr��"��=i/��8�p� ����M�#h8��y�Qt�!�#߈-D,ƣ�8sr�x�1C�"��>/6�o��E������v�r	�1����^F0c�1�I��3 ��n�3e!2w����w�=� �$��"B�+c!��g��\��&�Ƅ8-�2nw�ÍRc��ںݠE��a\��7 �l.����t_R�����&�I��;�<+^�+E����>����a���3F��.`.@�b�l�K��P�Fܯ~s��q֞�ql����bĩ�;;�se/]�f1n�ktS�[H��0�r���9š`��pԺY8<���s�83khc�������}dΘfad�p?c1O�u�<WQW{��y��d��'�j�D2���2	�8$�=cJ�#�>�6��i�4s�_�wz����N�fcN�k�I��)C�FqW"�����q�����4.a3����v�Fj��R���L?�D8�x�qLp�px.�����?����@n�������a��c��9��ғ�+�G��� r����"��w�*!��L�WPA5@0L^�a��vR�� 5�K����ƀn��e"sk4�����q����K��X&�ΫL NL,^FKa�x��kG½�h�bA׆��\l]F�_U�I<�n��t]�j4�Gв5�1`���0��&g��GH%4�����QJ�?��&����`��40t��`�0ϥY���:-�Rz53�?".0ȍ�x�ܦ|�8LLm"��1u˦ֆ{��~+�8gA�NM>����ƃ<�\�R�_0��kܻ��uډ|�uaǡf;�l��=K3<#��L����Q�)U�����O=P(�����_q����9���t��R��e�pzu����q��-��6d���b
�v�d�������s��ӔPP�`w��6��o`{��8��,3gq^�-�X�~vr���j�V
��G�F{<��M�Qds�H!'�kJ;�`d�6B����	d���!)�	��p���)^�SP�Þ�>���o	�B+�}�]��ˮp{�ظٕl�9�P/��v�E�P��wU!��3�{�u�Is��"I�N���r� r��I�ĳ^k�����(�P����I1j �w��S̀AP�i�x!�"����I#ڎ8�Af�q���D���F�m�����,D��D{��(l@ qވ�1�;UȪ�����F���e�+kX�Ǹ_�*M-g��b��0k�,a �SL�h����G�&����QQ�U��#ֽ����{�1�I)�M�6���jþ�u�<O����GM(�l���/8F�.��3��5Z�N���l���@�g?	���0(�g���1�̎��}E��6��ތ�j�פ��c��q#���[�u�p�a��-��U���vO��iD�q'��%v����,2	�m��m��m���̇I�v�6NQ7+�A�$`�8Fq���������=�CG�]���A�G�d�q�4p&�g�q#�r38��.d�a��N�a�::�5�c�܋z�*!���]�*��}�''�N���J�		"=�H�Z&E&+4�Fغf�c�({��"�	b��+�}^�/L6�l�oY҈��=@ �h`pdBa�c��^��c�yK�5PnD��f�z�n�}f��Q9ƃk@sMp6���n�5���E�\�(8�i�5�x����t��'dUD���ɉ��\qΨ�
cP�����6�^��d�/����)� ������"�mGc���c;"�q���"�{��5�_;��<���|&�@j�m$��ٽ xf����G��dR�Q�!j
,���~�;�*>Ə0�ǆя8ǩHd��Ӂ��vJ���ٳ�~!+�ke90D�W��W$s���Srý��=�9CL�dI$/p8�%Ŏ�<#A���e��Gz��ky�[y����g����s�ߺ�6�cQ�kw��N�ϻ�8��y�R8��+
q�s���3��e��o��h��\�С$�4K���XG~{����'�������������n ۏ���M��|�O�� '>��{��{�~�s���E�]`;߱���Kn�Qn�����`�+��!S'�:���g����L�y���8�#��ƌŪ����O9����ʛ�HJ�3�]����t�[�����I�@��0��7S)QX&���0(�t3�c^�kwc:���R#�L@4��㨥�랍
}1]pÂ؏��1�Ô��/�~�]���W�q�q%J7�H)�j��Q��#���܈�����u�6=,a��(�/�u�v��0��Lq���=d)��yġ���8�����)�7���;�Fij�\���+,�(�5?p.
����Qʽ�̈́�.v:��ġ[h���Ӊ��
%��s"����$�?)�>>����wf��S�9�g)AAA�T�\�*�Kr�.*��ג���]�jW���ܷR� � � B)L���_G�
'w_���J4X��>5��CT���܉'�c+%� � � �&z���\֠�<�/�[��%�EU��{�~�W��*� � � ���o��1~���E+��M2-��S��^��(=]1vR� � � B1��i�h�Hf�>�Z�pK|� n�>+w�K[,9��&W� � � BtXZ�Fr����[���q�I�f�|�ud�UG	� � � Q��{�Q5��+��k�eR�S���������v�xYo����+���6X�����b���Rk���J�/��R�e�����Zw�uU�|��7z�ؤ�_��Ze��2�<a��(k�Fe�5�Tu��UI��W_���9���p-���lY_9)x&x6��k��H
�%I�~b�`�H�%Xg�uT�:���#�+����9/i�.]��yN��A��_}�4�u�yIQ�^=��j��$�	}?�o��G�`b&AZ������/_��ļ�=��Y~���%�/��bX�{MV5��ʹ,��0S�@� �n���p�#�.T�|�I�߽�����*���]'N�]�c0���Z$��ŋ�|��$ӤIՠA���k�$�p\�h��;wn�ߍ��8Ҙ칟&L���B��j�J?I��4s�L}M�Q�Fj�7֢*Ip�|���j֬Y�7�oӦMS�K�,Q�'O��8A�s?�5>͞=[K�l��f���#A�q̘1#��F�7k�,�k�5�2eJ�
1ղeK�L$����'x�ㆱi��7O�q�ӊ�>}z�"g�v�m��\1mڴ��O�o��>���%�������l(�FS�̀���8�W��.9�q�Y��́8�b�-�~�TZ�h��?N�΀ܺu�D�A�����6m�$>��F�m�V�7.V���mܸqj���͛����v�)�l��~���t^�!i'��=sq>��s�H��6ܿ�HG��%v�g�E\"=Mqn�g��8E:�!��\�喿�$��s�$3�lpܷk�N�;66�n�9�ܤ�=����*N��8ǩ�d��/�)��\ߤ�$������D$:�8�d�M��{m�k@� e����H�[�},�fq
��r��AM?��È�S���tz��v1X'M�T�H7�aZF��S�q�6q�t#ΓN���n\"݈s":qGQ����)ҍ8O�8E��I�S�0��%�����8E��i�Hǐ'c�T(��~Z}��S�+p
�%�mq�&��q�t#�9�4�S�q�&-�4p���T�n��4a�\HQ�c�V5���ޮ�	��F��Pӏ��(�8����]�`A��Q.qn�`-U����%��%�q��r�sw�������%��%�q��r�sC"�\���H/�87p?C)"݈�y9�C��K�����8D�-��A"�\���~�"�N�Fy�h�-��%�^��<����*�r�s``3S1"����P�H/�87�*��-����r�sºX�^nqn(U��[�J���RDz�Ź��t��b���[�J���RDz�Ź�T�^nqn(E��[�J����~�(�9Ie�N�44�˝�L
��qʋD�3@Ĺ�X��qn(F�gE���Y�bDzVĹ���qn(V�gE���Y�bDzVĹ���QEzVĹ���qn����?F���g���k�mlg���^�X۵cl㔦$-iӢ��6	�U�CQS��B���*�)�����"hR�&@��@ڦ���6����^�6�����wwz��:�̾y3sߛsߏt�fwg���޽�{ﻷI�"�J��nEΕz$݊�+�H�9WR�t)d�17��,ѥ3:T�H~��%9Wj�tkr��"���\�UҭɹR��[�s�I�&�J���8��Y�s�I�&�J-�nMΕZ%ݚ�+�H�59Wj�tkr��*���\�EҭɹR��[�s%%IOL~n�&�R����p�R��=<���2,ʹWҭʹG�UZ�ɹWҗ-[FK�,!�đt�r�đt�r���%�V�\�#�V�\�#�V�\�+�V�\�#�V�\�#�V�\�+�V�\�#�V�\�#�V�\IA��a���,�A�V ����`:e�,'*�X�s���[�s%J�UV�ʹRMҭ˹%���\��t�r�T�t�r�DI�u9W�$ݺ�+�$ݺ�+Q�n]Ε(I�.�J5I�.�J��[�s%Jҭ˹���Oᐌh3e�.
ؘ��;�D��IgK�~.������gr��'�^�\�$�^�\OҽȹRIҽȹRIҽȹ2��{�s���{�s���{�se<I�"�J%I�"���.R��ɋ�+�I�9W*I�9W*I�9W��k8�l��cv��i	O&l����8�(c�+v�A<<ɹR.���\)�t�wOr��K�79WJ%ݛ�+��.x�s�\ҽɹR*���\)�t���$�J�����Z���Q*���\���xG�FFF\ɹR.���\)�tIG��\)�t�!eB/r�$(�)�\������~j����W8�C�C���@jx�sE%]2}9or�H�W*���M��t)�h���t)�tww��sE�\�J�����K�[OOyE$]
�]]]��\QI��=�g��Jz___^t�ɔ"�.�����\QI��N��=�t�����$��{C�	iA��J�T�Je�G��n�.W�\Y��������&O�_�l
�-��{#�W9W���-�� �I�,�g!T��y)""Y�, �x�8,EDd����,<cE�%<#�����UjKI���Jz?]�p!�*��:��;�S�(��*.�M1!���lr���Zc
     @V���1�]j^>��e�uAk)K��Ĝ����s�\�(#��H��r       P�����=A��
c��T�OX��7���:s+����       �<V������r'(��@SW�^o���0l䝝�'>H_�fR|��cT��       P2 ��Th��7s,��RA�1�L<ب�.��D����yO       �׷��t�r����h>`��Kw���)�#���<��b������       Hc��\VE�e�&�u�#�,ӇyCG�qAVr<���Ԉ�%�	�v���3	�;9�N��;��)��z�`�w��Ү��d����mb.�;[�O�ˣv�,Y4g��]�����L��۝cz��Q�rAtz�xi�8l{���hj�X�w~�7����W��9Ñ�9t���i#�L�8F�D~gpx_��i������j���V��{9�[�y^G�N����Y>�O����m<�GH^a���銩����u����MO��G�wn�DO'/L�7O�MO��v�����˵��}����!��]��sl
��[�-"�m���� ��r�d�_��r˯�~��֛��w~������q�6�+D��eY�gr&������6�q�@^��~h�iA_��!�PEF�F&�����8�uA_ǂ>�c$�;R`�{oϟ=\�Zln�0-��m���فV�v� uU�̝lZ��ͺ\�Z�r`�iA�4�zz�J7����K�3�ZeI�yA�v-vi�-�Վa,G�}E� �xote��=����[7�O�F	��3��W�Y���P��(�8eٽ�%}�|�8�
       ��'�{�������9��Y;\.�Oq�C�&[������49�O���        	d��ؽ^`I�C�}�)��m��̡�'�2'ox/�ti�����u�����Q^|��       �;,�x��:v��d�G���亶+/TzI៩Ђ��� �#w�A��(��]�T�        Y��x�]��� �ٽ���	o��7+	�#wp��X'����Z������%ߡ        ��g9�c'�v��d�W^<����{��^���S�ο���Ia]�������m�OF���$/����        ���P��v����x_���s|�~z���Ȕ4R0�d��k9fް��o�]����?HM��A���ǧ8�       �f���E��;����;���>^<�q*�f7ǣ򡢠�	��;��?^���e���s��m|���cJ��2*t��v'�      �w2��#�k2.ڟ�+^�)6�n⸕�'�͎r<��zY~�j���
5�؉���'�y^ޖ��}��)����?F�p        �^ן帎��>�����(oKo�BK~;��L3���ø��'�y��]����9�7s����"/���=z#��i����&*��$��?0��X�D�N#ӌ��1�qZ��h�����4q�Ә�k����.��>A��jz"��1��d��W;�j�@��d��'=��OO1�Oc�&J�8�ݘ����1�?=Y�'�XeY��F�&_��0���y� ����%�����C^�~���ӥ�~W{��KORA��di1>�'�5^�=ǿh3=�×����
��ˠw��� ^�==�9|��z�����%�8I�흞Ϝ�0)���s�;/Ϝh�Dz���B��>?�kχg.]�����ԫItBM��G���3�sYHO��I��g�~�!.h��/������'�od��y���_O���fe 28�=���t>��(�l�ҡ���q/o� /�r<ñ����x��ߕ�3��(���6��        xEj7�EO|��Y�����+�cq�4�µ�=�e�DM�>!S��_>pz����y��XN�!��(���o��=��!90�����WP���w�1       ���*��9d��3��Ex���t�o+���Kc�����/��?Q�˪�.����>L�A�Rs��]        @�E�l�$�ೕ�k�u��X�e��         �p��Av�}��KЋ|�C^�_M         ��z��4����؂�+9������{�	         q���;Q_��]$��Y���?~���9�?H�Pgg'����oxx�����3������J޹|�2M�4�<��c��T�0�_�pog%=�t�ޟQYHO###4qbMEJsHZ�4���|��|�p_�:u�N�>M 8~��7��Ts���υ+���y�Ɓs��%z��i�ƍn%��ٳ�u�VZ�r%͛7�<"�+��B�'O��k׺������+}$=M��s������Eoo/-\��<"�=���j>�[��&L�4�j|<H���6Ќ3�#����glOO-Y��<""�m۶|A~���n����{��a�L���gwuu���iN����^{�.^�HW_}�[9<~�8�ܹ����*�=�YS:7���-[���ժU�ݻw��Vғ��<"r.��<oA�q��ϛ�վXW��+�<��dr3FX (�%�̙3y9!�_�&�*��Ν��,a����o�eJ���M�U�ED$��I�ʹ���g��.r����?�5�(�*�����o��M�U�O�<��Y��%]�|׮]y9���M�5��W�
�$]���ѣ��E=J�������ǣ�Xo��r>00����K^��ח���ɛ�C΃#��|~?Η�ͤ]���\ �(�r.h�/x��r9N�8�N�K�\!�&�r�x��r94��$�r.�5�&�r�x��r9�ǒ'I/�sA���$]�\�C��7I/�s��$�T�}�z��R9W:�_z�t��u�y�z�t�ypNq<�����C�9od��7���8>J������˹�I�+ɹ�I���\�$��\�"��\�$��r�x��Jr�x��Jr�x��r9W<Iz%9W�Hz%9W<Iz��+�$���+�$�\�O�9�tk�ߟ]�?5������.��/e�w�9
p�IO��%�IO��%�uI��sŃ��'�I��sź�Gɹ�A�ǓsŃ�Gɹb]ң�\� ��ɹ"�a�'�Jz��+$}<9W<H:�<8�����n��$���2�m]@`,Kz59W,Kz9W,Kz59W,Kz9W�Jz9W,K�.�gϞ�߳,�q�\�*�q�\�,���\�,�q�\�*�q�\�,���\��Ǫ�ǑsŲ�W�sŲ�C΃���3|�g=�,�����?�s�$ cQ��ʹbQ�k�sŢ�ǕsŢ��"�5I�E���W��fZ�"�ȹbM�k�sŢ�ǕsE�˒��f͚E�E�k�^��+%=��+%�9W,Jz\9W,J:�<(��n��ߟG�]IМ�w�\X� �G�k9lX��$�V9W,Iz=r�X��Z�\�$��ȹbE��sŒ��*�J�I�G�+�^��+�$�V9WJ�'7[��sŊ��#�%I�U�K�^��+"�r�W��fS��+�$r�	��9�6tB��Z�C�������+��a�d�^��+$�9W,Hz�r�X��F�\i��7"�I�W��ވ�+͖�F�\� ��ʹbA��s�ْވ�+$�^9W,Hz#r��}%4S��sł�C΃!2��cߛυXa"9V��万����!��0% Ah��7*�J3%=��+���6�ʹ�LI!�J�$=��+���6�ʹ�LI!�J�$=��+͔�F�\i����s�Y�BΕfJz�r�4S�Cȹ�LIoTΕfJ:�<�~��g|o�Zi���-�[,�7��Tx7ӱ� �JzZ��s�TҧL�BiR���+VPZ��sE%]2ʴ)�JzGG���r�Cȹ��5k�PZ��s�T��"��+*�i䥰(��r�4C�CɹR*�i�.	)�J�ܹs)-v��Aǎ��RIO�Z��s�T����R���4+�CɹR*�i]�y$���q+ߗB�<���w�^<�	O�K�����)=�L�|i�I�6[�o��V09WT�-ZT��ۖ�DC#�.���y���ɘC"b#¼t�Ҡ��JH�W*D�B#��Fzd2��
� �@�F�K�_�#4Z��ۛV%��_�O!�\I��顡�`�������GI��G�ȶ��'4�SE�OI_IG���H��ɳ)��t�ȑ��=�J�<g[[[)I$��sJ��tIOI��~IO!+{)Ƚ�Օ�$RR�#�%�QI��l����ŋ�k9�銳��.�'_Jj#����y�O�����;9��-��<�4��߹s'yF��;RJ�0�&Rh�r� $!	i"������L�W�g�#�J�4���$*��D*}B��h"UIT���H���{F$M{�xF�9d/�f ��==ei��.��8��e���M5��i^<͢./����a�e6�       �nE�e���c�d�:��t�$�Y�e��[8��Eү��       $��$n*�����U��-��t�Jm��    IEND�B`�PK
     !M[�����"  �"  /   images/53dea2ad-2eb7-451c-84a6-1b4fef66a2aa.png�PNG

   IHDR   d   7   ���   	pHYs  P�  P���Dm   tEXtSoftware www.inkscape.org��<  "pIDATx���y��U��w�{kJ���2UBI !�DA"�Jd��->�x*v�zK]�G���(�����2=��L �		�TU�JU���y�o��w�͗�M���֩���θ��9_L��+5�W��5G4�(����e֬Y���&���RZZj�g̘a����e���2g��:u�����Hy�AY�`�L�8�ʎ;&��s�9GƎ+�x\>l�K�,���+������r��Jn^�h����K�.���l-���2�����;O23�dpp�����om��ӵlP���csg�h4j�w�ޭm2m.�HTzz��^nn�,\�P�G�����7N�ϟo}���[�)S�HQQ�����ظ�=��q�����_i�s�|[��ͺJ�� �	F�1a�1c�Xx�XXɬ�l�S�Z=RQ��Sh�Y0i޼y2~�x�q�+�a,�z�@���@�!MK"��ŋ+���l(�����ٸCq��r��u>�A�H�,[���g�V/-.˗/���?''����͑��?_222$;{��5//W.����-�YY�V�H��u��6��q���0�4wh^�ȟ�|S,� 2k�]��!�h��Ha�X���%S
��92a���˼	ݒ�5$�+�����d��.�Ȯ#AY��-��)]})�ɲ2ڮ��!�m19X�i���ʧ���PC�m�P�e)%ʥ�ڥ�:Kꆲ�3 �guȎC��8r��䳋:ek�rNN�jж�������dDe�y�,�
D�d��9]��4G;V�� �O���7��w�ebn�O��AQ6��Wf��-�y�_(=��_5�i^��7���� �n��͚�I<7�-��5/	) ��7*������D�o0�T��֮���2�5uƴ^@�^������ֵ���j���?bm�,�IMkz�����ֲ�����BY��,�+�g�2AE�����o "5:n��As�m�%J�2��О.i^���K�!�5wiި�� d��r�[���G����$��:�|i�[�Uy^.ӦM��h����`��;Xnb��=���w���#2{�,9�:���z����c2w�\�l�1���*55��6�8ioo���F����ri--&����V˴^CC��1�YiM�Dӆ���Z9k@�2SJj2$�KU�QC�4Յ�E�ޑ#�U�d��)S���E����$Bt�$�W�ieD��r�.S��7��G#c��[��1�d����	F8�yn,�f�k���>��!uuu���ۍu#
��"E�¦(M�켌z�nkkS�5����ߔ�d�e�_6���@�2�eMM���!�������̥������˨G�C�����{ƟX]ce�G?<#��GOOOr<tW���ѣ&j}��-�&� #�7J�%�5Y����VF�CHk֬�ɓ'KGG����UV�Ze� Q ```@e|�TWW�$���.��@HXO^x�!�	�J�-2�����I�&Y�|�)}�0.ϔ1(�� ���\������A" ���!��7s����&�qS�  �{�����ߖ�+W�a\<�����e�]fk���\7j~D����I�OwK`�"��k�O	̍*!> �۹s�Mj0,�Hʜ
��ar��Ƃ $�c2��ȑ#f��t��2�ji�����Y�����7�'��(q�5sչ���ː��/c�y��qP���q*��Oo��:���3S1�ܦM�nEEE���jY�b����R�|�4�^s��F��!P�W�u:���L��
۷o��3eήd8��x�y��7�>�#C5P�@��:~�������p�|�W�Y+�Xc ,F���Ha�!��ӧ�5��HΘ,��Ҏ�"J }:^�X{z��6����+=�u�$ѥ����1ي �'��I��ի�c�b��Ա�y��Ek�_�D����3f���
���?6?�#e�	��C�i�o���}��GM����ʰ>J���/���۸��;�AE�����7��"9����p�O�[�t�\��+�y�����wݩH��}�{�$�.bq ���A~�ؘ������Ųt�4y�߶�u�_&ͪI�n���޸B^���5C}����?m��CG��l_������4�c�{���d���!�Z>K��@��v����Ȗm�r�Wj��2sz��9Y���۴ϕ�g����������{[+����Lfj�Jԉ���?6j$�%�s�=&b ����M,̜9S~������G��&s��G�'D��wݭm��&�QJ�ʯ�_v��u"5�Tt��%tx�������,�}�.,6N����Xd��=*��&���ϕ���R~4OV_|��4E��[6WJFd��OwTT���k��õJ�铤���RV���Jsg@�\8K�VFd����{��4��sR��}Α���[���5Wɡ}��}KYe��_����,+�!b�u��OJ�=v�%��ۏ�裏Ј�;�cJ�ӟ��a��_V�8 /���YF���Ɔz�U t�	n�K�n8�O�K��3S��ʄ��f���~e����}�����O��.��⠽�û����uލ�=���$��=	`"*r�z �y!=H�"��$�cP�"=���Fl��,Dy"���S�����-]�0�"LsLe�Ͽ�zx���G���:a���z	�7|\��immI*g�h�o��v.&�/��GB� �caڟ��C�yb{����3k�-��w�}��)���@�m�f��e �o|�V��q@O���$bS�'��S�k<��To�����C��M
�瞓/}�Kf����@☄^�nD�y���Q=��w1�aEbQ�j3��wl#���N3Y�.���@F����{fـ0��[o���r�k&e�@��{v�R|4)6|�,��yHߵh6��ON���|��&"`�c���φ����7�h����ȸ�~�/��3�! ��'HÄf.�f>�"R"C�B�;v���b���$wn�'i��L楗^2�v�ڵ��� �I���!��#����Sp�#�����r��9�%��O�ؒb�b�*����`����ȑ�!㤫���l~2�""��  Y����(u@\򤓉6'�A_n��;iw*.9U�.�z�	�|�<O�x�(y�q�7ʖ-[N@��Z[Z�M4A���:��T),��|2�7����(0��f������;ԏQ��tu�����7������%Ͼ�S-���7s[�bE@ڎ��!I�S���snIe�p�W�g֍�{6\�8�H��b�' ������N	+'�`ee�Y6tx:�6�������֜�C�u�2$��Y2�S���x������Y1ɻl����͔%�L5����������N����l�}(���l�aY҇��F�wR2�S)1!懄>��C�h��;s$��ݻ��S�?l���g�Z�H}�|[,Y�Rٻ���d�6�ʴ�C*͎��<5i�U��7���y�ޛ�`�&�2��D���@�H��	�aU(n�!�0Q�D\��[��l����w�+W^y���]w�e�qx'��P�٦��xA����ʖw�J���7�"l�|���Y5�ӓ�R�ψʄA����C�y������1\<:W����b�t��[�\����l��C�J���|g<�C-�9�ǽ��+���j�!N"�sVu���Ǩ���=�|O(��UY{�W_s��^u�������;,+�Н��e�ª�ќ3g�\�z�4V&�Iy��/��֓Ň#���y����!��I������APD��r��>����5����o���f`�Hxd�.����c�=&�<�ƫ���@�QW�R�u�� ������G�(�w��Gy��-���o}��ҧ�xB���ԔdKK�E @<2��k�Qjk�l�K�_�{A��X�Es�X�����"X���J��,J�p�ъF�<��~��%A��g,���k��`g#��<g͞=���m.? Jc�@�G-	0ʭ���$�p�"s��0�_� ��hl��Y3gK_o��< ��כܣ�@��nQ�l�Al F���l�ٛ�Қ:�d�x��a�A 2�|
�1X�w$?$�:�ebD�;� -�d�B/�����
"*�S:q�m O�`�'f{�j�q� ����=��s<^��,++I�8�)/�/���V&��cǪl;��K/M�E����6�S4�I&7� /K��l��Om����b�X4 eN��7z�Յ��b��aB��d��1@8�t:��Aux��
s
	d���|�:7���e�$�D����d�V�ѣUI3��VW�Z蜄N*Tj�8X����d��ܴ^������7����[o��a^�r�/_&6�ju�;������3�N�p�U��&�5B0�SI0`�.N|˙� �}�T��$�J����+s&���N�?��(2�Y��e�I"�W���_�w� ۷o�쉾���O����ig�%N��|��f�r���O`7�A[8F֬�cGsR%��C�$c8��C��������Ɔ���$���Mo��"���p���ş��v�|�o8�	����roy�Ώ�U�O�+�/��[p��c�:���t�=�q�ֹ ۴i֗�+_c�u��t=�&��0)��t/��(��S?]����yx���.� r��jY�l������-e�?���vp|���R�|�9���9���w���,��}���[! ?�;�ԁ\)�� yg�|�s��=���w�A�4�L֭��&WVv�8��1*�6�i�k�~J{�{gg�^�[�y��4I���7������:��ks��3��;��9pg�q�<:aTd+¹�x��K��͛7'�x4ł�,���<��}�D��L�l��T��$'�f�d�o�vB9�[�Α���H�����2�x�)�;���'p�w(���c�9�Q"��J=t�h�*F�4�/�d(���r8��d`s?��1 � y��ǒTw�Й&��c�G���N�>������ma���+�P��$Qq�vJ(yp1,
InR;�����c�vGd�Xsd�i�h82h�E� <�n�р=j
`38,Ɯ�����?�`�<|�� ')';C.��Hj��)ڧ�bF���F���a��uE�}���i���T퉠�E2<����pVcS�mK,�ܕ�P����'�|2����;aSz�D�I�&���9Ë&!68���IZ�z�W���k�R���&;'�޸�''�ᦨǲ\�x�NH�|ox�c~ZнW�7my�@��k֬U6�ׅ֞�)�/�~?�����s7�f�IvAzkk�9��p�4_=�u�]$-]�ޛN�ׇa��u1w�+e��.p�CF���ew36j;6H�_����P^8��s(�M*"�L������{v�A�+ s�z���D
[r�v4	J\�r��;�q,Z�0����+7�؉�R�� W8��)�Bq��8��<��.�8^x�tɈ7'KV�?_j�e4����z�'��)w��_������?��IC�"��X'NYpD�#6n��qԁ�	@�N9���Q���S��h#	MS�(5N%uu�I�F?9���5�u�p�D�� ��!� )~P���x�D��� [�.�-o�,8/6
��@wR�?��S�?�)ɞᐃ�w
;��q��h����'���������@� ��������㔢�%��+/�T� 0,�����\;�0<���{2��c1�`��	XZ���hYă��ڜ�FY�>V�,o���'M�'l�~���7���w�5'	������<��AO�cN��ku��w�<qB}��7��htPuG����U)zlR�q�=56wʿ?�S.��̓j9!��9έ�(�a^�Dc Ġ���)���n4J=pF�k�)���ݵk�\q�F�t�����5�\m�.Qx[�l=#�)�Pf͞m~D{{�����x��\���QnzY�1�LN��\�i�X[z��!���ALn�;���� ��p
F'5c ����j�(����Kd����M"䡇2d`��s��eQǘ$�w��i�=��W��&�1
��%8 44DT�u��2��	@���l�u��C�w��a1��@41�v9q��n�l$���W���XuHը8b��2�@�'�Һu��.;rq�%r��!���{F���2}/:g��ٽK�[�%��(CL�TU�*��Y�������"��&I{��ɣ�Wn�Z�C�xh�nG����{�X[��X����ok�-�h_]�6��i1����O�S����p�5:{��g��?��-�@)sWJ:��/���"�1���{���;� i��-v�=��E�{����?�)�o��¡?�@�D��?����K�ͪ�I�wt���XnW1�.1��a�bU1�_��I����nR�q�!fӦM����&ĭXڀ��F�|o��G�\�`!�`�V+{�|b'T�9D��ܹ˨������O�: ]$����Q��7s�-��C� <��g����X��Sb�.��q���+A7����o$�d��#1���o��V�����0�pi�3�''���	����GW	�p�ȯ�s<�& jZ�����͕g�:��񹤧�F�?%B��v,@�'�}h(�Is_�|D�}���ZX��@"J�;(??��=�#����T�`�|��7n�h��������0�&��S�T�2���|��=	 �D�'��]P�AL�Y�s`<8D�!�p�� �."}BC�����{��6��k���g��!?�я��1 ��<|���;����H8�{��N��wؠ ����C�	���loo_�T��t�b@�7ސ@x�!��U�M�v�r PW�(����%�䉿| �a�46u��ͫ�6|"3�Ȣ�)��3[e��n�:<$�^�(��fI��,������_]-7�ܜ-�-xz�����-�o�{���������3�d��VG�to����er��.�Y�Չ�hė���n��6�Ǯ|�~��X�'�0�GM�{':�`g�> �/��5�T����-�
k$ l���u���޶mۓN�By��]��;�j��˃m��m��?����v�0a����N�R���Aff�|�����I�1�m����6$/m|��|����[�hlD�}`����+)���7�R��ȯެ\�f�������]}I1�KB-���C�9�湚�Y�pe��w���I� �.��rS��^{�Ev����N��'f�肛� Āg�t�����17n�`�n��H�\gN��R�!�T�}��_���&ikm��7�r��|RbD�q7�Ζ- CgaX@$lJ���{���믿a��H�K,S7|85ÁA��f ��LD�2��/7
�W�O2q}�w�S��$���<ŷ��~I�fͅ#a.  ��t��������"���I���Y ���=�nx�׌��N �{LZ���C���m|%"8>4(�� �4��-��Q��}��Z��BԀgNUr��q;:��q%��z@
Ҁ�p�K��bg{��PX/D����`�:͉mO�7�e��!�X���apFA<���i�����|�t�Ꙥ�$��&
�6l�`�P���2Bh��X< g�hD%��m0�$��@,�F�S��v?��~B�2 J=?�ȸ����pm���[%�M�Dz&�OK�i�)�!�Q� M��� 0�{Vv�����^�ó�se�v�.#3؛��갽DA4=���������fZ��tE���s����mjb$Q���`���)ត_���Civ�`p��ʘ�#,ħ���Iܔ�b�'M�K;��_����7]���\�!-�
M�ć�-ґ�"P*E��@r�R͗i~-T�u�	!�˦Ș��-c2��`}��� ���.��L+��]j*��R?d���E�T$�`N�1߄�y:����w��<3/N��V������A9gZ�mJ�±�"��i]Rѐ)�pf���Z<�[��f�$E�}K�xj���4D����H�J��dQ��>)��+%U�F ��̊�ɬ��R�e
e9�2�`@ʪ3�:��e�ȸ�9P�mđ@�?h��|#�z���B�@�����%�e��2�d�G�C��=h�
�b���w�xW�e�ǝ-��3h���dN4��Bz�^c����ײ�.��� ^`�O�뗺6��z�(`R��}u��?��`Pv�N���}q�?)�_��)���nv4��U�%����hB��/�ٸ%��\f,.�$^���o������˅�g5�)�� ��H�{;��[%�#���+�C|Hٴ1���Xd��c�x_m �"i�Z�d��Tei��F+�q$7�>-k��my|bQz���ݨ���|s���Ղ�z��/��ޮd�|���̞�;]�\�(+0�tuv$O��QVh�X�x��_�h�-��.I����Ҏ�F����2�^��ʽ�3[�;��Nb�* ʫ[���%���9�DZ�Ȩ��D>�?��M3����/g����PrX;��B^��4r�= KBibY��~V�&|���o"��!\�s�X,�CY�.�@�a�����n�����8��Q�E�B&��_%�9���O-R�a����e ��y��2��_q�Oq� d@����������    IEND�B`�PK
     !M[��F�} �} /   images/b63deb06-c33f-4ae3-8f73-25229955b1c1.png�PNG

   IHDR  �  D   CzWF   sBIT|d�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<    IDATx���{��y^�'�U�Y�s�����xYD�F@P��;�Ჱ�ll쮷]5aa�V$��uB�n�0ܼ��������,������Ow�S��2뒷�#+�T�S��\��WY��Dd����'�'N�y�����   @�	I~>�J   `!���3�<S:   eUK   ��OK��(�   P�S��zs�    ���  ��ޒ�g�|b�     ,�7$��$�[:   �(�  ,�?��ǒ\-    �'y_��(  �2j�   P�W%yg�V�     p�F�/O�����  �9Sp  X<_���'��    �QM�G29�����   p��  G%��M��    p�U�|v�ߐ䇒���  �<(4   ,�z��L򕥃    �#xO��%9(  ����  p��d2�ꭅs    ����$_�d�t   Ύ�;  ��v=ɏ'�=��    �)��$_����A   8
�   ��'&��I>�t    8E�$��I>\:   ��Z:    g�w'��Qn   ����$?��3J  ��)�  \>oM�I^W8    ���I�M�/(  ��U+   �S��$ߟd�t    8cK�{6�*�  �S��  py��I�i�f�     pNjI�x�^��+�  �S��  p9��Ç�   �h*I�p�V�S8   �I�  `�}K���ɉ<    XD�$oI�II�[6
   �C�  `~U���$�t    �@~ �ےJ  ��)�  ̧z�wfr�    8�}I�<�A�    <w  ��SO�I��t    ���]�/N�+�  ����  0_���7��    s�?fr,m�t   ��;  ��XI�I�R:    ̑&��$/�  �kSp  �kI~<��/    �Ї3)��z�    �:w  ���$�6��(    �سI>7�ӥ�   p��   xUoJ�3Qn   ���	I~.ɛK  ���  .�OL�I~K�     pI<��'��g��   p2w  ���S��?�o.    .�k����@�    �K�  ����I~&�[&    �o-ɏ&���A   8N�  �b�=I�M��J   �Kn5ɏ$����   p��;  ���Ln�|�t    X�$?�䏗  �D�t    �$_��2�    ��z�/O�t�_*�  `�)�  ���I�?�iQ    ���e2�]�  �0w  ���d��I�T:    ,�Z&��>��g  XX
�   �L����A    �$I5�I�J�   �(�  ���    ��;  @A
�   ��OdRn_*    8��;  @!
�   �K�    �C5ɗ$�p��  ΍�;  ��Qn   ��R�d���;  �9Qp  8_����,�    <%w  �s��  p��0�&i�    <�i���$�T8  ����  p�� �r{�t    �LK���;  ��Qp  8;��    p�Ԓ��(�  �w  ��񇓼'��    p�(�  �!w  �ӧ�    �۴��kI>X8  ����  p���   `1(�  �w  �������;��     �B�  ��)�  ��v    XLJ�   �H�  ��)�   �bSr  8%��   ���&��$��A  NK��H�ٜ���jY^^>�O�s�ھ���T���륥����{�ܥ�����Z���۫�jZ��}�W*��ۧ���~��888H��?�?ooo/���^����� {{{�֍F����[���������h4�o��`������\ �9t��O%yo�    �J�  ����$�:�z�  @9��˩�j���G�V+�J�XI��l޳=9�P}R��V�ssΓ��GK��j����џ��\F����=%��_���e0�^��^��ce�����*�O�?Z���ߟ�����?��E�n�a>6 p��%��$?Z:  �<Rp  x4�=ɿKr�p ������=e񥥥Y�{Z����l?Z@����I�z�~��>��ۛ�f�ƙv`��P�����p��x<+�-�O�G�G�?-����������t���?}�i�=  ��n�/N�S��   �w  �����L�7� �mZ�>߽<�>�P~�>�{��<�}&���~�?+�O�f������|������y�t���� � v���$?[:  �<Qp  x8o���'� �"x�ݞM,�N+�N:�N_^^N�Z��?�����d�ݯ�qMK��i�w�~��$���I�t�����i����f8foo��G��[I>/�J  �
�   �Z��'���A ��f3�Ng6�|�|t��t���������3�|� xu���t�|�׻gB}�۽g:�t�`0����=S鷷�3J< ��+I�P�_,  `(�  <�+I~*��(�ӳ���f�����,//�^���j���N'�z=KKK���v{V@o�Z���'m .�i�}ww7��`6I~0�����g?{{{������z�{�3-����Ϧ�pi��䳓|�t  ��N�  �u��D��(`ѝ4��t�N�s�4����v�=������Z�V�# �׫M��N��n�{J����l�t���݌F��`�}4�<|  �>�  ^�R���t% ´H�l6�n�ge󥥥c��ѧ�ޯ� �㙖ޏ��f��"�����b���M_�P>�I����A   .*w  ���'yO�/.༴��,//��j��jeyy9�v{�z���j���dyy9��˳������ ���������������eoo/�����z��ݝ=�ۺ��׻���}M�ȯdRr�t  ��H�  �d�$�J򕥃 <���v�=�����2��~����������Z���(  ,��t�����S�N�?i����́$��$ۥ�   \4
�   '�'I��t�r�V��I�G��O�����cէ�wOTo6��?
  \�~6!~gg�ش�����z��z�ٺ�������f8��(����I>?�^�    ��;  ���A�?_:p�M'�7��٤����O���G�]__O���  \D��(����&������l�۷og4������I�8��j   9�
  p��&��J� �G�ٜ�ϧ��z�>[wA���z��(�  �lZx?� �<t�ty{{;����G ���%y[�q�    ��;  �-�7�<������GK��v;�v;�V+�N'�Vk�  �"������nz�މ��'�O���g`��#�W�  p(�  L�wI�a�j� �hN��~wY�u  ���j��.�����F���a��I��t  ���  �?��;��J�y��%���������  �ˣ�㷶�2KǇy5��.��\:  @I
�  ����I�/I�t(�R��J����-]�n�S�8�   ���������3{L_O��G�����$_�䟕  P���  �"{K�K�)N��&�oll�ʕ+'NS_[[K�Z-  �� S�oݺ�����>������i$�ϓ�`�    %(�  ��%��$�J�W����������euuu65����N'����t\�  ��x������������v������[:6���$_��'K  8o
�  �"��$�w�7����t:���x���W�\I��.   .�n�����{��O��O�O��ߺu�td�f��N򋥃   �'w  `�\M�I>�t�_�����F666f���$��֯���R�Oq   �G�~?�nwVx������f677O\�֭���ұ�/&��$)  �8�  ,�N������j6��	�G'�}LK���   ����?�?]w�������ұ�x�N�I^.  �<8  ,�z��%���A8{G���b�݅��E�����j�ұ   f��i���+�-��z�ܾ};�Ѩtl��J�$;��   �5w  `T��;��J��4����fcc#kkkY[[��^]]=�����F�Q:2   ���F������N����������lmmekk+�oߞ��}�v���JG���D&<��   �%w  `|k���t�k6�������FVVVf��	�G_����R�OX   ��5���v���9�����N677s�������&��$��A   Ίv   p���$�t�E�l6��t�n�����+W�̊�W�\I�ݞٯ^��Z�V:2    ����+��z�ܺukV��.�z�ܾ};�Ѩt�E������!   Ί�;  p��Iޙ�Z:ȼZ^^���F���f����r�ʕ���fuu5���Y__O��,   ���A�������۷oϞ777�������ܾ};�o����N���o$���!   ΂�;  pY�5ɏ&Y.��»r�J��ַfuu5W�\��766��   8�2�t:���Vnݺ�_��_ȇ?������(�W%���A   N[�t   �3𻒼'���>��e_�e�c    �@��z�\��+W�[�h4�L5�?K�B�[8  ����   p�>1�'Y/d^����
   ��acc�t�y�L��I~G�    �I�  �L6��X�7�2O���JG    �$�U=��$�:�'�  pj� �ˢ��I~k� ��T,    .
Ǫ�SI~<ɕ�A   NC�t   �SPI�]I�`� �h}}�t ���V��T*��\�TR���y�I�ﻟ�h��x|���px��x��x<{߫= p~�zd���G��5�~�(   �G�  ��^��(b^��3 pT�VK�ZM�Z�-�j��.O���'��_��>��%��`��h��h��p��p8[�ߺ�2  fuu5�jՅ����g2�O%���O  �9��  ̻�1�_(b���3 \~���G�ZM�ј-���4�T*��q/�ii��l>������>2^u��I�  ��R�duu5�o�.e^}y�oJ��J  xT
�  �<�#I�n���m�`~-�O��G�^O�V�MV��J�2�o������-�������������� �e������x�J������A   �3  ��zs��I�hc4I�4��Z��1 �����~R����A����I��� `^mll��h���[�|4ɏ�  ��� �y�T��&Y+d�mll��  �R�+�7���s��L�Z-��V��V�eyy������X���� ���988H���x<>��  �OE#ɻ���$�_�,   E�  �7KI�e��P:�e��� 8k����>}LK�J�tD.�J�2���ݦ�����Y�}�|ppP - �q
�f#���|F��g  x`
�  �<�d2u���rY8Y ���4����,--��lfyy�$v.��*�O��O'�O�M} ΋cV�ꓓ�H��N�W8  �Qp  ��7'���!.'����>-�O���̻J�2���Q�� �yr�����$ߙ�O�  � � �y�g����!.����� �B�V�Y^^���R���g˕J�t48W�+��F�Y�}oo/{{{����h4*� ��:_���I�f�    �E�  ����%�$;eN��Z�X�}yy9�fS�^E�ZM��J�՚��{����^vww3& �cVg�o$y&�;J  x5
�  �E�[�|O�f� ���� ,�Z��V�u���h4JǂK�~��fޕ��W���^:�eUI��|8�O�  p_
�  �Ev%�%�Z:�e���"�T*i6�i�Zi��Y^^��x��f��f��u��� �^/������x<.� �(VWWS�V3�JG���I~ �g%���Y   N��  \T�$?��SJ��VWWKG �SW�׳���v�=��^�VK�NP�׳��6��r<g?�^/{{{��� �b�T*YYY���V�(��F��%��$��  pw  ���I>�t�����w�j�X���j�V���<�J�����,//������fwwwV|7� .���U���30�9I\Q  \(
�  �E��$�t�ˮZ�fee�t x(�B{��J��I��2�.�z������݇F�Q�������n����݌F��)�Ӷ����{�t����%��$_Y:  �Q
�  �E�UI�z�����(p�U���d�v��v��J�R:PP�Z��}p�ڵ����������eww7��tL �1������(ޖ�W�|C�   3
�  �E�$ߖD��8I�ET��f��v����%�v�UU*�,//gyyyVx���K��Sx�9��չ��$O'yg�    ��;  pq��$�I�*dQ8I�EP�T����N��N�cB;��*����wOx�Ny�ǥc �auu�t�ERM�$�&���Y   � �a#ɏ$�V:�"q��R�.�W�n����'��F�Yٽ�����tD ����#,��$ߗ��%y�p  `�)�  �U�|W�O)d�8I�y��j�B{��I��(	X`�j5����>�A��nvvv��v3' �
y"�'��I���   L�  (��%���!��� ��J��V�����t:�,//��gj��g���$�u:��j��0��z��׳����x����Y�}��+ p�g(�&yg�/-  X\
�  @I_��ϗ�����JG �9:�}ee%��C���x4�pg���8�����3�vg�L�g4���������~F������f��[7��I��#a�lo�?f��=��lo�3�Y�^O��~�}�'\�X?���I��VVR�V���tR=,��z_����v{V�-/��lN�7��^�R���|�J���u�\k�S��OL/�i�Z�~�z���쾳�c�; �#����I��$__:  ��.��c  `Q|f���R:ȢRp�q5�ͬ��dee%�v;��_�gaZ���L
�;;���{{�z����������x8����ϊ���-�O�ݣ�݌����2:8(���x0�`k��=q��;�DgoV��TR_YI2)ԧZMmy9�F�X�q���n'�ZjKK�.-M�?,��:�T��Z�T��&?��J�јl�VO��$�Z-kkkY[[�x<�����ׅ ��2����M�KI��t  `�(�  %�)�$Y.d����ÚN6^YY���j�����`{;����`k+���;��~���w
��nF�A�;;�"s�7{���x8�`kk6u|t�$s�lF��)�o���V'����;e����Z�T��YѾ��6+�ז�S]ZJke%K�zvG�����'���r}�ٜL�w� <�V��F���]w���T��#�/gRt  87
�  �yk&��$�+dљ�����j�t:Y]]���J��j�H�dtp�a��a����V��ެ|>�ޞ�lOZ���po/Ý���&��#�v`��F�I��[�%�=|��N��aٽ�nO��G
����Ia�p�}��J��Jm���N��N��u�p X$����y�f��l-�{�|z�!  �s��  ��o�������� �5-�O'��,��4������v�������ome��u|����d����J5I��1Τ��K���g��g����:�_m6Si4R�t&����T��f��k�v�N*'�wX��	� \p���
��}r��M�I���   B�  8O_��+K� �V�i�ۥc p��j����dmm-�N'��(=�4-}����wv2��ɠ�ͨכl�ٙ���s�0o*I�Ӳ�t��i4�F�~F�����Tj��d�Ng2M�՚=���;������]Z��M����������%��$�t  `1(�  ��O&�_J�`bmm�� \�z=���Y[[K�՚�n�zw��oo�ylme��3������t�ay}���a���`P��\G��9�����t��=]�R�Φ�W'�O���_��k�S;�0_�tN�� pY������1�J�/
�   ��;  p>5�?OR-������ 8c�~2�p���ͨ��xw7��0����z������E���n�Ψ�/�ҹ��~����Qv��hrW���Gz�ѸS~��_?,�O��G��WWS�;�p�9�u�T���$L�g  .9G�  ���I�t8� ������e��;+�����^F��d�����p�����po�؟UM�J�N����*� ��J&/��d�i�}T0W	�~?����77���VkR~o�'e�Ng��#    IDAT��p�zd�|�p����� s�1����=I>=��   ���;  p�*I�'�o+������L'�vv2<|�,�6{�v3>�<�j&��i��r
���wt��8��{7����`�y0���pw���W�VS;,��WWg����kw���Zg�	 x-&�_HoH�%��$n�  �	w  �,��$_\:�rr��L���^/���nݚMP��ܙ�~8i}���v2>���R&�OieRr`~-��2)����ڛxh��(������}�N'���cS�k�Τ ����]�I�%f �Ð��3���$�M�   ���  ��/I�5�Cp2�w�Ѣ���>������[���[[�F�����I����V8 ������$��)��������J��+W���H��Q�x�a]h.�/%�{��   ���;  p>%�w����w�2�log�����v��Y������_��dԟ����3)�w� �eWK�r��'�fRv��y�R|��L}uu2~m-���IA~u5���ɺ����j*���%g����MI>��J  .�  ���I�$��p
��Evt�zs3�[�f��;;�u���������NV?m�$˙�[��X,�L�����4�n&���%CqjF9x�����_m4�8�_�t�,����_��Z�u��N����<��tT3��'��$�^8  p�(�  ���I~[��:�w�Ӹ�Os3�â��p��tݰ��p����wwKG�p�\A։ۣ 01��i9�I�Iv2������ٿq#�7n���F�%�z�����������h��j��땎��]O�/���${��   ���;  p��!ɗ��ks{g�Q�����3���`k+�۷3��N�����������GS�dR{'��; �O-���� ���$�qԨ��hs3����ܷ�h������z�kki��M�76R��Hcc#���4�^Mui���lmmM�����I�E��,�  �$� ����I�f�<܁�����������͌��ܺ�a��a�wg��V�#u��2���N�:| �y��Ȥ�ދQ�<�Q���͛�߼����=~6���<\6xTkkky�J�ൽ-�H�-��   �O�  8�����o��0��3py����LW���`{;��������o�����x8,y��2�Ծr� �����N�A&SݻI���=�d�j�1��ʝ絵4�^�L��r%�É���Qkkk�#��)�/$���A  ���|  <�f�Hr�t���0߆������ܺ���f�_z)���72�vK��-eRj7���TO��d-�n&EwS�9o�~?�/����_~�}��l�ѩ�Ǟ�\I��T',ǲ�J=�w%��I��  ��>  ����$�^:�IA����q���߼��[�ҿys�����+�L�o�ʨ�/��TM�Τ��(���R��wP;���;���G%C�	�n�n��{�U���������k��{���I	���4�^M��`�9�5w^��@�?7�  ��;  �8�l���t���j��pƃA��ln��p����w����R^y%��Y3�R{;��P^=�F�Lu�N�2:��`k+����~���ݧ�h���ө��+W�|��;��]K�Z=����Pp�K����&�K��   �I�  xToN�J��᭯��� �ʸ�OssVV�>�߸1�Ⱦ����_NFf�.�j�V&��f�, p�j���� �����1����F�o�x�������a!~�p]���TM��"k�[!�L�]��   �G�  xk��f�S:��+xp�^/��7'�[���f7o��֭��J�ne�햎�T���j&�A ����z&E��$��������y�U��w:�_���իi\���k����ki\���k�./�SbX�5̭J����M򋅳   sF�  xX�$�N�J�јz�nw2q��i��	�/��A�W:&s��ɴ�v&�0`U3�Hk%�n&E�����bt�t������O�ј�ߟxb6���w&�_�����9���gX�\�$��$�'���   ��;  �>����Spg��ܼ���/g�p���+����sp�f�ne40���Qɤо�I� .���v&��${I�%C�7����F�o�8y�J%���;S߯^M����T�k�Ҹz5�����rI�r,k�}j��H�奃   �C�  x(�ה��qR�y7���OZ�q#�/�d�:箖�(���e �̖�LƯv��&�95��$���]��zj++�I����+W����.âX]]M�Z�h4*�G�eI��$�R:  0� ��d�w&i���YYY)�k<ep�V�_~9��i���7s��+��J^y%��;ZSV#�R{'�ɶ �H�I֓�%�e2ս_4\>�� ��|�gNܧ�j�y�z��x"���'S�_����_�����9���S�T�j��u<`��I~.�ϗ  \|
�  ���&��$o(��g�;%��ɤ������b^z)/����l\P�$��L��EW��b�N��L���E�b��f��g���'n�6w&�?�T�old��'���i^��T\���X]]Up��$ߛ�w&�U8  p�)�  ��|v���9K�~?����߸��728�:8-���r��Μie2��Y: \P���A��$�Pިߟ��l���g{�^O���c���a�}��'Ӹv-�j�@r8���j^x��1x|��I����g  .0w  �|Q���tNG�ZM��)�96�2x��%�χ���ۥ#©�$igRlw  L3��L~�>4��b��I*�ZW��y�z��xb�|X�o^��ƕ+眘E玄���'��$o/  ����  ^͛�|{#�.�N���[����~�ľ��s��g����d5I�p �W�$��>��d��{��|���_z);����l�N�o>�D��zjR�����SO��nH�e掄��7$��$��p  ��Rp  �{�\/��c�S�^/�/����<{�?��>��)�]-w�����Qˤ辖;E�a�D�i9:~���g{�әL{�����i���<Ǵ.�z�w&�]I^,�  ��9   ��[�|V��.Ӯ�x<)<���������ǳ��g��U:\�LJ�$�o g��d=��{7����h"����y&�g��g[�ZMcccRz��4�z*KO=��'�L�u�K��*����1�K�u�X�ܸ�  pw  �$_��ϗ��s2�r�����ǲ���MJ��?���</���@uN�Ȥd�. H%�J&���lE��x4��͛9�y3;��+�l���f���f���%��)���K�s���$_[:  p�(�  w��$ߞɐ=.'�_�֭���},�g��,?��";< �v (��IɽEw�^����lo'O?}϶j���Of��o����/=�dׯ�Rq_���1�K�'��$��t  ��Pp  ��&��$WJ�l88?��������{���~�����_Ϡ�-�R#�j&e: �b�ݏNt�M\t�~?{�=��瞻g[�ٜL|?�������
��������֥VK�Iޜ���Y  �B�  8��$���!8;+++�#p���t?��t���}����y&��z<.�v �����0�F�}���>��=۪�z�O<1)�?�T�^��,=�T�_�z��9�֥�d&�W>7ɸp  �Pp  ��0�_*��e���q��K���f�C�ί�j�>��d����F��L�r ��Pt��h0����g�����V��Ҽv-�'���ߘ�7�i2����1����$_���s   ��;  �$�O�I���p��<?�~?�8��>���O���2:8�pw7/��A�W:"\J�� p9(��e<f�ƍ�߸��~�ضz�=�����O��o|cZozSO<������t:�V��F��p��!�O'���9  ��� �J����6�\rn�|�F{{���Cn��ϥ�k��Q_�K#�z�V�  ���ݻ��e� f��e𑏤���[_m6��������4L|?3�J%+++���*��UO�]Iޜd�p  � w  ��|^����Fs37~����O�d������B����v5 ��:�3��v�a�8�����3�=�̱����,��i��MY:Z|�v�P��E�}a|B&Y��t  �w  Xl���o���1��t�����������/����q`�Ԓ�&Y�b; ,�J��w2��>*����^z�HzwM|��Z�I��G�W�J:�nX(,�_H�J  �Pp ��u5ɻ�4J�|T��t:��1.��G>�_��o���ϗ���I�}�p X<�L�t�lgRvWt.���nv�~:;O?}l}���շ�%o�3�P����p��$?���)  8� ����$o,����tR��s|n������߮�稚d-�듬�A- `�}`=���.�|t����_(cn(�/��$ߝ��[  �c�;  ,����J��|9	x
��<��w�Ə�X�$�0*�Lg]KR+� ��jI�d�}a+I7ɸh"����K��l��r�9���~s���*  8_�] ����I�^:�oee�t��6��w�C��Q;���W�� ��i���$˅� <��h���+c.8����*�Y:  p�Lp ���L�L��`�|t�?��|�]���/��a)���3 ��j$y"�^��$��q ^��sϥ�ɟ\:ƅ���B��$�O�L�   ��Pp �������t�p�7���3������_.B=�Z\� ���L��Mr;ɰl������r�t�9���B[K��I>+~� �B��   ��?��-�r�|8��<�_���Sn�sP��L��� ��N��'وc�Ŵ�쳥#���g$���!  ���8  ,��I�Y�`�9	����>O�7�����Q�R�$Yɤp�~� �,T��frA�J|� .���+a.�@��I�9�C   gO�  û39��s��wv�o��z��Q�R[N�T�+q�
 8?�L�<��������͌vwKǸ��"�_�ߙ�u�  �%��!  \~5��AyN>�����ٿq�t����ʞH�(� X\�L��\��$�0g�c+���k�Z���cP�'$yG�  ��Rp ���w'�[�Cp1�����p��~��y���/.���R�
g �j�]e��a��JG��*�J:�N�\_��K�   Ύcu  py-%yW�u�C&�����ތG��1���$y]��$��Y  �V��{��2��P	���-���$��t  �l(� ���-I>�t.�_�pw7�?���1�RYʤ(v5B _-��-O�g����@�9b%�wg�+  �d�[��g�΃$�����'�y��*+��2�>zfZ3�:G:-����&8���#K^H\���]�»f9�?�`�]9 ��� )4BB��cFs�Y��u��GfUWOWwWwg���|ޯ����|���ROW���<� `8}�����p]�-��b�ӟV�Z����rXQ�g�  �^�j�3.s ��	��C�/򤤟�   ��(�   �g\��qJ:���8�1Bm��_�� <G҈�S۹�  ���?׌��s �RmwW��=����8�?��F�    ���   0|�����[���3�XG ZBҤ��8�  �����7EI�q ï|�u������JJY   �=�7   ���$�w�!>L���V���ښu` �%MH*H�   �v�}\R�8��ut��u���n�I��:   ���   �I��u��wVY[�Z-��@q$�H���4�  �/i��a~0�^�0������;�!1�   q�     ����F�� �X����Ɔu`����:� p,�L��n���d�8�$ɉ�K�O^s�@���|�۞�⸮�.�s|_n�|O����>?9�LJ���%7���=V�ۻ��t��=��rLc���N�VS�\�$5�u5�/4����wj�x,�^*���8~��/5�w�+WRNRJҶ��m C�	�w�9.܁#�_I�I��   w   `8�G�߰��b����J\ n�U�J��ګ� ��tQ<���K����r;E��8��DB����}�	�q���r�qqۉ����S_�X������hk�U���<n��jV���f�r�q�z�h_��qt���N��V*I����j6jH���j��j�|�f���ڧ��_RQҁ�]I\��A�)���pE��|�u    ��;   0�^!�}�!n�SSPq����R ��R{R��g&�K��z^�>�A�X�+�J�L6������TJ�����N��ssy=����@��R����l�0I�`�)ͷ�uՏ�����4�ە���'���}��@�rY�rY��=����#)#)��4��m �����Ύ�\�:Jhq���~Hҿ�   ��Qp   ���D��:�VwV/��# ��4�viT�﷋��t�P�%�����y&Ӟ|����=�}|�T�fO��N1=��7��0 Lbɤ�L��h�j6���o��e5U��o?>U�ot
�����㣣%�r��9GG�׸�r��%�.�oK���0��׮Qp��q�>$��%=o   ����   �_��r�?��l�_�� ���4���c��b�����X:���ȍ�y2��Ȉ��t�q���dڟ�J���dK����{ @w9��x6��"�M��K��Ǎ���t�NI�V*����W�s�88P}�}�L�G�%$MJ*Iڗ�� �U���<�u��J$�<O�Z�:
�-#�$�E|;   w   `p�N�OY��``��۫�J:|�aN�i��S�=� 8��*�ɴ���l������d�v���L�]<�|K���u���� @��i�����������|�vR���;y��������;�����Zu��WRNRJҖ$*� �Eyy�:B荌�hkk�:��Mj�?��u    ���;   0��'��=Ĺ0���v?�9��M�@(���j�9cj{4�TP?u;�s�i� �p8���/��k4+��S��OO�otn��]���T��U�s߬T��'<�����%�� Χ��b!�2�w��/I����b   ����   �_���Lp����>g�@Ҹ8Y4b���\�d��I��%u
� ��� �R>_�߬VU?�����z~X.Bu$�HJHږ��?���~wr�=HJ�CI���0�   ��f	   �7I���!08\�U���Zͦ������:��N= |�x\��⣣'�Ǐ�\��s�l���y�zl� ���
��{����ލ�{��Z����[�TR��GG=��<8ORAҁ��܇������j��r	�(�E���5��#���    8?
�   �`II�=�<�A:���8�1B���gC[��������~{���T�ν_(ȟ����*62"��1^>/�u�� `�xw�`f�?�^*���q�����Ɔ*���"����}u}]����	n�H���4�r_���i�TY]Urq�:IhQp�}�YI�����   �|X�   ˇ%=b��E����җ�# &\I9I��p�XL��X�6>.|��8�k��s�vI���u'�� @d_Tv^��#�wwU��Vu{��xg�侶�ݾ�����Z����Ӎi�;b�;�[���)���p|I �U�j�Y    �w   `p�7�~�:O&���Z{�A	���S������(����������r
&&?.���+>:j  tQ,�T,�T05u�ϩ�﫶�uS齶���Ύ��B|}gG��Mն���9*���:Ls�b��e��ƹ.ܧ'$�_�{��    �;
�   �`��o�����֪�t��3�1���IUt����2�՟��?1�x6��P�?1��Ȉ�lV~��`rRN��d  ��♌♌��<�Y������ޞ�����V*������ummmimu�=A�TR��\w �*++�B�s]x ?-�O$}�:   �;c�   �4g��m�϶����YcGbDCRҘ�1���Mߤ������(   '\ߗ_( qF    IDAT�/�z�3��V�Z^^����j���Ƿ�ݓǵӏwvT����`Qp�3�u��%����K�(   b�  ���FI�o��E��~�k���s՞���v���~��)� ��������]W���>�Y.��ݏK���v1~{�=5~kK�R�2<0 ����B�s]x@�Iz���X   p{�  �p�H����(��m��v@�C.�4�h����S?%/���  �@��ǕN�u��u����&
��LM������j;;����ꥒ�����v������Gp�GG����B�����.�'��/I��   �lQZ�   �oJZ���Ƣ��(�cX9�F$e;��b�e/S�[��:  @WA���%mllhssS�V�+_7�N+�N+1;{��Z�Z������ޞj�%���wvT��QugG�RI�z�+� ܬ��L��68ׅ.�$���WHb{    �(�   ��vI��u>�nU]_W�T��t����v�:�����.ɉR�  ;�qT(��dt��uU������������w=������n������������R�Ύ�������h�!90<����c�Y�%���*��u��%�O��Z   p+
�   @8%$��$�:_&���:�<c躌���5��X�u�S����  ��dR.\���vvv���">2��Ȉssw<�qp�Zg�{}{�=��~}�dJ|���Sr �*kk�Bmdd��;��g$�����   �f�  �p�����C`80��V�>k蚸�S�� �~臬#   ��뺚����Ȉ���U�׭#ݳX:�X:����m�i�j'%�Zg
|mkK��]U77U��7�8��R^Y��j###��ذ����K�=I���V#   @�Pp   ��m���u&����k_�� tEJҘ���G��4��W[�   �L&�.hyyY����q���<����B��5������4��榪[[�u׶�T��}-U
�w�@t��%�O�~�:   �(�   ᒐ���vW]亮��u�Pi�j:�|�:�@\���)� !0��wZG   �x<���y���jeeE�f�:R�ŒI�fg�7~{[��U��T=~���~~wWj���8���Z���XG	%:���+�����     �(�   �����J��z��^P�^���7�u5��+5=���v��T�޶�e"�J��-�b  ���訒ɤ�^��J�b't�3�U��L�om�ڹն�T��Tu{[���>�nh�˪����嬣�wt�/����:Iѻr   !
�   @x<)�ǬC`���w��g��� ܞ���?>.o|\~>//��76&?����k��G��o����7~�a`[�o~�b)�� ���}_KKKZ__��֖u���x���)SS�=������*��nn����~~cC�j���%��
��9/��k$���>h    w    ,\I��Y�pI���B��k_�����ӊ�r�r9���r9�s9Ţ�\N�Ą� ���b��fffnY�///���ۯ����ۭ#   �s]W���J�RZ^^V�Ѱ�4T�S�o�����Ύ*kk��������Ύ���nl��d 0�]umMz�1����bg���K�cI/��    @�   ��Jz�u
�:|�y�R�TJ��q���	��S��ޯcJ�Ӛ��Q<~�i�����F�������&�   �122�D"��ׯ����:N���i��i%fg5����~2~kK��MU66T�ظ1	~cC�Z� 9®��j!����IK�7���   0F�   �����X��pb��f�rY��u�@���/䏏��?1!?��76�.���r�����8���*
�=��_��{��K_��   n�y��������8�8��z��.������~r_��Pu}�|D�WV�#���Co��j�   ��   ���$z�	�nV�rEj��c �\�k���

�Ţ�\��.��[��433s�-����>%
��+^a   ��Q�PP:�ֵk�T�׭#��٬�٬�.��z��@յ�v�}mM��m�vv�e���ըT���Pe��m�k!z�7$�GI\e   ��   ��Q��)z�����\�� #�+����{Xd�YMOO�uݻ�	��  �(�J顇ҵk�tpp`(�N+y�¹��uUVWOJ��j�ω�������}��zPp�=6&�%��    @TQp   �LI�%�nw��5e
�C+�N����-vrR��o�x�f>�?�����v�!�R/ZG   �X,���mnnj}}]-v�Z�[��������V����8�F��Z�$ot�:J�PpG�m��l   �"
�   ���MҸu7�nvt��u�'otTA� obB~>/ob�]^��;�o�x�����{�(���g{�(�\�Wbr�:  �����J&��v����u�S��h�������j������I����ݞ"��
�gH��r]WM.�@o}XҟI*Y   ���;   `��Hz�u�t:m!Tʗ/[G�m��מ�^,�/�����bQ��YG�t:���Y�b�{���K�z�(�33��Z�   (�TJ.\еk�txxh!��b�����j5U77O
��UU�������(���8Z*���<��u��qG�dR�Q0ܦ%����   Dw   ��2�>d�@����֖�8Lycc���z�s�
�r9�x&������}}�ѕ+]N3833�   R<����׵��i��<SS
���|�V*��)����T��kk����9�𩮮ZG�t:M����%�����:   %�  ���uIs�!�L�:Bh1���\߿i�_,*��8yn���߫X,�����%��c��  p��Q�XT2������u$8/����*}��-�5+����WN�߫j5��Kye�:Bhe2���Y���s%����I�g   "��;   �_OJ�!��
�7Dy�u7ųY��JLM�/N��^�(ot�:�@H&�����������V�7���   0�FFF��^��J�bC�%�畜���V�����M��ӏ�����;���%����X   ���;   �?Ǔ^�9}�8�M�6����f�wJ��Ԕ�bQ��I�SS�%���Z.���Ԕ�y�U��6�T�:  �P�}_KKKZ]]��ΎuD������5r��������U�~����'��1*�o��;�콒����Y   ��b   �?�T�+�C :��\׵��o�e�
:�`r��LMɥ��u�XLSSS�f�]�����m  ��u5==�d2���U5�M�H�$��7:��ŋ
ff"[po�˪��k��>K�=����A   �(��   �Ǽ�n���Z��*���1L���Mʾ�U���$%�>�}_sss
���_7�����u  �����H$t��U�j5�8�M��I���������/x�����9   ��Ǹ+   �?~G:s�e�g�buCyyY�F�:���7��^�z%��(��Q:�օ�^n��V�'kRp  �D"�.��$B'�N+ῗ��U���J��# �>$i�:   0�(�   ��NI�:��B��+W�#�r\W�������5??/����X"ѓ�;�  z&�i~~^�|�:
p?�S�+++�Bid�y"01!��!   �aG�   譌�߲�hb���ׯ[G0�OL���q��u]��̨X,�q������=��a�w  ��rG�bQ���=�`�WA��Lp?�`��Iz�u   `�qF
   �!i�:��E���t��㟡~�}_KKK��{E�����u  �H�f�ZXXP<��D�����ù/r%�+I|�   z��;   �;����C ���~Cey�:��$��H�RZZZRЧ�y,���ʊZ��u  �HH&��p႒ɤuD\P,ZG0���q����3�!   �aE�   ��\`�)Vm�V+��Lp�\.����b���g�'��&  �Q<���r��uDX05e�L�\V�T��:��4o   F�  ���QI���hc������f�j�Tbv�:��rG333�����8}}�(�%����   ��8����M~�$)����`*��%�N����%�/�!   �aD�   �1I�0��-�S��Ubz�:�P:�b9::j��n*e�aqt��u  �H�ؽ��x6�X"a�L��o��u]%�I��wH�N�   ����   t�oH*X� (��U���#�
���x�u������L҃�	���2w   3�TJKKK
"����/�#�a�����!�[���   tw   �������! ��c�O8K��ZG:�tZKKK�/��y���V�r�:  @������%.�F_SS��Pp?���~�:   0L(�   ��H�]I�эP�d��-�ss��J.�����\����7>n����O[G   �<�u5??���1�(����u3����/��OKz�:   0,�Wc  ���^i8�����uSLp��q455���i9�cG��OLXG0UYYQ�T��  y�?+OF�x��	"�����f!�8��	$}�:   0,(�   �Q��s�!�c����<��Z������1L%ff�#�X,�����M��y�����U�   �����b16�C��Ţu3��5�c�w���%}�u   `Pp   ��7%����Hcq����*5��1�8���ۻ��}---��)����~�:   N�d2ZXXP<���!LMYG0��[��i���}HR�:   0�(�   ��u�0�q-����#�������u���J����$?�����1�   |��.\��D"aC�����w�~���[G
��YI�   :
�   ��q$}X�l��aq����b�T0=ma`���jaaA�X�:�m�A���uSLp  �x<���E���XG��q�Ţu
3Lp�CR�H�c�!   �AF	   x0?&�5�!�cq������W>���̌Ǳ�rWɹ9���^�j�:   �ຮ����筣`�$&'�#��Pp�CR��i   d�  �����s�!�����v��l�T�	���qMMM�8@� ����L�����1   p�bQ�.$����}���[G�< ľY�wZ�    w   ���I��Y(��U">�����O���rO/�KR�_��   �����\��I<8�.J�*�oA�!�[��   � �,   p�����C �C�]j���g�T05ea �b1����x�'�K���h   ��f5??�X,f.ʿ�V66�j6�c�
��r��~�:   0�(�   ����[� ng�����f�����c����ZZZR*���r_�ss���~�s�   pN�TJ����<�:
X"��[��j���1B��;��%q   �G�  �{����j��d2i�\u}�:���ԔǱ�j�dRKKK����^)���֖�ׯ[�   �9A���%%	�(P�Ą�x�:��J��w�X,S�1�;IK��u   `�Pp   �MZүZ� ��UR%�܃�i���N�����X,f���㊳c�J_��u   ܃x<���E~w��q���u
3Q߱�,�[��%}�u   `�Pp   ���K���M��k�'�SS�B+��i~~^�;�E���Qp  <��j~~^�l�:
P09i�L�w�;w G҇%��   ���c%   菇$��u�<�ɤus��/�&��~���	MOO�q�(]�~����(�  $�q4;;�|>o&����Xw
�OH�1�   ����   �߇$%�C ��������399��nc������V}o�:   �S�XT�X����G��^������R)��y����u   `Pp   ��풾�:p^Q_�k�Z�nnZ�0�OMYG�q4==���q�(=�wIͦJ���u
   <�|>�)~��9%"\p���g�d2������   � ��   ܝ#郝{ ���b��uS��5k5�f�lV�d�:F(8����Y�r�;+}�u�P���g�#   ����ivvV��)ܙ����}5���c�J�=`����ǬC    aG�   ����j��y��'UVW�#�
"<��4�u5??����(=卍���c���  0�٬����,c����	9�;R]_��*�t�:p/<I�   �]t�   �'-�}�!�{���,�Fy�ݱX,�����,r3�]���W�88��  �.�d2������d�='W|�w꺛�_��bQ��C�[$�M�   @�Qp   ������C ��	�R%���Op���Z\\T2����7ܥV����?o   ]�J�����x<n!
��T�֬#�
��0�>$�or   �mPp   noQ�?��+�X�MDx����Z\\T�Q�*��#�Ba�3���   �.
�@����}�:
B(���Q���Ř��uQҏY�    �;   p{�%):�142��usՈ/��]�r�%����Ba��;  �Љ�E��;/��#~���(�c�����u    �(�   g{��wX� �ܥJ�'�SS��.�JiiiI�x4wvN.-)Ƃ����%����c   �����H$�� D��	�f(�ߌ�;ظ�_�   �Q4W}  �;s$�f�8Q/��j5�vw�c��%����X��t:���9�nt��w\W�G��g?k�V����|F����:	�ЬV�,��8<T��P�VS��H��(�ժ�ڏ���j6�j6U�ߗ$��U5+IR��P�z�}l��V�����-��8u왙�e5;�{�׫�[���Rr���X2y��n<.�E?���i����ǎ���L5�%�r=O���M$��b'@�29��~�sL,��G��@�� @�b1-..����:�|_@��Q�ྱ!�Z���K��;�K������    aB�   ��Hz�u�~e:������y#*(�#���F�x��������X�ZU��@��C�K%5��ԬT�88h�v\N��T��W�V;)�7�u�K%�����u������s�<H���ˉ�o��;���i�(�����(�H�M$�d�&��ǩ�b�̍�FF��DB��_�	�������]�zU|ψ����{Z�VSmgG�ؘu�P���<_�Ŏ�   �M(�   7$��u�AD}Q/��t������r��F�x�:B(�|�S��Ъ�����q9��@�����>nt�;>��y���;M:�ph��j�˒��ϭ0�T�]v��>�&�%�e2�w^s��vi��Z|dD�tZ�ų���##r=�G)��뺚����������jF�g����������g����6I��   �w   �f�TҢu�AD��^Y[��`*��{&����,��S2/}�u�P8�tI��U�o�ӬTT/���RI�RI�����O�~r���t�J�s1E7
���+����ApR�?���Y�FFn�?~��g�4��!I�����U^]��b�����ŋ�1B#�NSpǠ�MI��ݭ)  �S8k   ܐ����!���d�#����B�:B�e2����q�(�����76����us۟��������f����j;;�mo��;���wvn*�����c�ԬVU�ظ�Ϗg27M����3�s9�cc�����˝�;\h�r]W���v���Y~�݂{���X*��6�c��J��H�#�    @Pp   n�%I��!��	�/�OMYG�l6�����y�K���[�0���S��_��-%�����Ǐwwo<��8:�N��������=����Tx����W��7:z��W,��Az �����,%���E޷S{����Q���"�%U��    �(�   m%��u�"_p�ܴ�`*Q,ZG���QMOOSn����^F�]��SOI����<�V������[[�nl����������������mȋF    IDATm���-5�֑���-����7⽱1���������	y������
�%�=L������U*���ςܙ�~���h��1/�]�~�:   `��;   ���|�@7D}A/�w��������'��WXG��֖��yF����:
B����.�������.�oo����PukK��U����2�z����9'�ƒɓһ��˛������

����z^����8��NO����q�G^��Lp�Y�>`��G��J��IN   @�   I����:���ɋp��U���m��Ba(�\N����1���}��x\�z�:���O~��{��vvT��T�S\������yRd?��Y�YG�si���]�r�c㣣���v�PhO������+>6��Xl���bH@j�܏o��Q��^��T���� �#�N[G �%+���~�:   `��;    }P+A
Q�VU�ܔZ-�f��I�]w<��K&�y�Q����j����?�����f���ꪪ�몬���'���4�f�j ��wwU����s���8���ML((������bQ~�(b���XǓ�%J�Q�G��ެ�T�ّ76f%(�c����ߒ��u   �
w   D��Hz�:�-Q_̫F|{�X���U���'��_�����.��/����x&cwЬVU]_o�66T�vM�S����mm��lZG��ЬVU�~]����x\<�mO�?�
J��ʟ�PP(�<�����Z��J��u�X|dD�DB�r�:�������}���$����e   �B�   Q���!�n�|�}s�:�)�
��l����)��W����us�z];O=��o��(�լ�T]]UyeE����_WumM��$������  �ꥒ��'�ǒISS�{��`jJ��)�[bfFn�15p��I�܇�_(����&���J_�h#�~NC���,�/��    (�   �~\�#�!�n�����֖uS�2EsddD333r�:�@}ի$ǑZ-�(�?�I
�=ԬTN&�]�z2q�������u Z��#>�����ǜ����Sbv�d�_((����}L�(9.��Z-���Y�AQ.�G|'��(�c9�~]���    (�   �R���u�ۢ��W����	�lddD��������)����^��bn����0�껻:�vM�k�T�~�=��3��������uD @ȝ����S����337��OM)��>�8(��Y���sG����z�������G��b��Q]_��Q?'������]��c   �7�
   ��-i�:�mQ_̋��`����4��.ɾ��%UVWu��J=��u�PjV�����:�zU���U>��N	 �c�J��S�]WA���쬒�����̍I��|c 9����9J�C,��
�Q?'���k�>*�-�   )�  EyI��:��T�:��(Op�g2r	��-�Nknn�r{�����Z����:F(l}��.��K%�;S؏oGW��//KM�� !�l�����ʊv?�[^v}_~��.��͝���J.,(F��'���Љr����O��91��%}���3�   �w   D��%�Z� z!�ӪZ-U���S����r���Q���OZG��O|Bs��}�1z�qp�.�w��/��ެV�# �3�j��������u|������Y��J-,�/Ò뺚��ӕ+Wtxxh]4ȿ?���Z��K�d2��^���'�b   �
�   ��I�:�+Q.��J%5k5�fuA?�JQnXTrqQG�.YG1W����8<TlP���Z������e]�rRb?.��ww� Zխ��E�_��-��A�����J��+ٹ%��P~Z��j~~^�/_��ёutI0��wC�^W}gG�ؘus����<�"|nCmN�?��A�    @�Pp  @�����u�W�ɤu3Qߖ{��ɤ���)��H��.�Y�i���J�o}�u�;��J'h�{N�=�.�_��F �f���g���3������%fg�z�!�zHɹ��4��i9��:�\���.]��r�l]�&�g2���[G1Q]_��ޑJ���E�^��I%�    @?Pp  @�|����:�KQގ���e����[G�'APn��k_��?�c����񏇢�^��R��^���ի:�|YG�/�|�*%v  B�Y��\x���S7�K&oL|_\TjiIɥ%����Z��tɽR�X�A��b��闼�:F(��i
�f����w[   ���;   ���$ŬC ���p���	�Ţu�s�}_���'��rO>)�u�j6�����˿��{���~|;x�Y>�ld7  ��ё�~ZO?}�k�lV��~�a%fgO&�'����B�XL���t�j��u< bB��=g�De}�:BhD��"��%���U�    @�Qp  @T�I�7[� z-�LZG0S��wb�:¹��q���+�D��GG�~��Q������^��������.]��K::�]���+WT/�S8  QU/�T���U���oz������pAɅ�.\�Fi!I��Lr����q� ��n�Rp?A����~I?b   �5V�  �"ɱ�Z&���`&�����Ŵ�� ����D��ORp����'��^/�t��s:xi��=��^���  ΩY��v�?1��C���=����*዗��x��K�.��hX��}��f����B��;"��ޭ�Y�    @/Qp  @|���X� z�u]%	�f����fC?��u]���)y�a�{�ku���[�����k�{�����)�.���N���I @�T76T����SO�x�u���U�ᇕ�p����r�X�'� ����._��&2� �w&��H�R��~�$����   �w   D�/Z �!�L�q��QA��a_�wGsss,4}�k�z����us���k�|�S:�z�]f�����++jQb  a�l���]��͏}����ܜ�/�o�<��ŋJ��H�]�[�ɤ���t���Z-�8�G����j���H���~Yҗ��    �B�   �^g�(��[���{{�1̄y!�q��̰�l$�Ji��/��g>c�\�Z��ǭc   ܿfSG�/���em����<K��\\T��e\�V��Eycc�aS:���̌�]�f�����n$/^m5�mo���b.���9�ڃ}�i   �
�   f�����K���ie�OLXG����)e�Y��6��7Pp  b��C�������я�<���Q��G�y�1�{L�����&�lV�FC+++�Qp�S<�Smk�:����&w1���^-��A   �^��  �a�}�^n�H�77�#�
�E�g���T.���ycox�^��߶�  �>+_�������O���9�PP�Sv�<��2�?��',�����hh}}�:
�AP(D�ྱ��ŋ�1�%�I�@?��~E�7[   z��;   �U\���C ��E�Z��a�����5���Pȼ�%�'&�;    Ҫ���Z_��_���s�Ą2�?���W���T��/��H����	5mE�0=���	�_��a"��E�Ey�"뿕�fIi   �6
�   V?,�a�@?Ey�J�a+��������p�^�:�}���I   BՍm��_��ޝx\#O<��7�Qcox�ҏ=&�u�Sژ��T�����u�C09i�L�w�;F��+��b   �6
�   F���X� �-���Q.�;N�
��tZ����1�"c_���  p.�z]��^��^/������{��5��7j��oV|t�:b_MOO�^�����:
�"L���6
7�=��Ϭ�    �D�   ��'$�[� �-ʋx�ܽ\N��Yǐ$%	����q�(x����z9��V�i   �����?�S�����<���*~۷i�-o�����z�q����^P�R���;��f(��E��"�E�   C&��	  `�����u�B������!�P�y����亜j#o|\����  �׬մ�������w�S��-z��Veu�:VϹ����y!��g�E�fj�B!ʻ"�^#�ۭC    �Ī3   ��OJ��X��"^�'������({��[�j   C�^*�����>��w�+�}����%�H=��5??�X,f�ፍɍGs���GG�1���q��Y��_�Ķ�   �  0LI�XI���L4+��c����jnn��0���XG   �j5Z��?��~�����i>��u��	�@sssr����8�#[�2�]R�w8D�}��wX�    ���;   ��?��aQ��^�޶�`�z����4��"}񢂩)�   V��6?�1}���[_}��T�~�:QO�R)��p�)���	�fj���B�s���)�   �  0,��@dEu����p�~rrR�l���q�G�o~�u
   �V����~T�]ߥ����ժu���f�*��1p� ��#~~�XTϏ_'�oY�    ���;   ��O��툸�.�ՙ�n��|^���&����[�#    "���.}�#��w�v>�)�8]��D��	�[[�B!��ǀS�/��  `Pp  �0HJz�u�ZT�/������Q���'�T,���  �9�|Y_����������q�jrrR###�1p��E�aP�ذ�
Q=?��2I�   <��u    ��%i�:`-��j�'��	�2���g"����T_�����r��6?�1�(x@�Ȉ⩔�x�����J��x\����f���ё$�~t�f�&I���~x�f�n�  DR��������O��_�Ee_�r�D]333�˗/��sl�Q.�onZG
�$�$����u   �~Qp  ��KI�I��5���y�u���=���<����u�n����V
�!�}�gg���VffF��I����y�cw}��Ͻ��j-�$�j��mc��`�mC�6�� `[� �2�0�$3����0���p29�$�2L�	�<,�L���q ����^��k_�>Twu�{�E�W���:G�dI%}�������/Q((����W��)��)��/�	+KKZ������ssZ����쬖''�t옖��ұcZ��k  @Z=vL��ַj��߬]oyKS��X�}_��㚘�P��	��XG0S��.�����,�U�>g   �.
�   �v����荒��̴s2],Ӯ]�J�v�;���j���Q��yʌ�������u�^s�F�=��2N�N+L��7>~��U���x�����¡C�}�1�>���T�\nSZ  �+��}�SZx�a��)h�T�����u��!�y�m**���S��V�^�Gv�	���#�/�w   t)V�  ����c�./ޭMMYG0�΂�����x�^�
��t�~�:J��b1�o�AśoV��땻�:�_w��.���R�_���_���Z�\���G5��i��I��E��  ��L�z�o�͟����w[�ٱD"���Q9r�:�Ӽ0T�ͪ�����z]ՙ�����i\<�Mb�;   �w   t�wI�tW�jU5���a�Ж�R��*��]wQpo� ���Ӟ�ҭ��p�*=�z���)�o�r��i�K^�q��ѣ:����C��Ci��A���8  p��Ç�Лޤ�~�w�{ֳ���X__�599i�iQ��d�]�ʧO;_pO����N�a1�   ]��;   �U$��!�N��t��쬓ێ�Վ	����*��H����u�&���ct�Xi��4���n�]�k����ֱ�e�Ɣ�5/{�$iejJ�����}�:��ojuz�8!  �$չ9=��w�)��J��ggǊŢ*��fff��8+���[�0Q>}Z�׻]=F\�͒���    �VQp  @��eIc�!�N��t���%�p`��ϟN�5<<��׀��S����V����u2cc~�s5|��ٿ_��;hlEr`@{^�)�s��7�����&��=իU�  �Z�\��տRuqQ#�|�u�R�\��Ғu'��d�NU����`��cd�|X�  Ѕ(�  ���g�$�N�*;^p�Z8Y=�k||\���5`�p�:���Y��
��>U��W�^�b���e�����Sn�>����Z�����{��Wt���V�\��  �4z��[^j�������yӡC����f�9Q�O�d�ӧ�#�s�pϔ�����    �VPp  @7z����!�N�rt�p��-�=�e�X,���q��ߒ�Gg(��Eܯ �o�v�s���w��{�X��Y�lV{_�R�}�KU^\�ѯ]���ou�[�R�R��  ڬQ��я~T�rY#�z�u�9��jbbB�Z�:�S\.�W(�3�����;   �w   t_���C ����T�'��٬�0l��z����qEQ���Fg��v��\Nչ9�(#=<�}�߯=/y��{�Z�qN��蚗�L׼�eZ��ב�~U��E�z�!�h  ��=�;�#?��+^a�fG�(����>�F�a�a�h���=F\��$�H��k   �,
�   �6o�t�u�Ӹ:���p��U醆���yr����?��_��uS��k����u<���H~,f	Z��~�����������:��/�����U�� ��F��G�R��[�ّT*���A�<y�:�3"��SS��%	���z�n�4�F�  �E�k   �ē�/�C ���Bruf�:��VL���r���M^t���w[G0��M>����E���_�﹇r{���ޭ[��n�����;?�q�~��yֱ  @�5�U=�h��ǭ��X�PP�ug��i���][YQme�:�)���\��\   ���w   t�_�t�u��Zpwy��x�'�'�I���4�9���o�]A6����u��z�st�/��F��GI����P��G��G����:����jkk��  @�Ԗ����ާg�ɟ(��q�����������
�=j�DyjJ�]��c�J�RZZZ��t��[ҽ�!   ��`�;   ���e �T.���*ss�1̄�BӞ+���S�u�*�u�u���|_c/x�^������4z���w���ݺ��]?��/��w�[�R�:  h��c���>�z�leG|��������c�5���nRqx�YLp.�nI϶   lw   t�WHz�u�S�Xp��ΪQ�Y�0�MyJ(�}�u��	3������/}I/��AO{�u$4Y��_7=�����t��>��޽֑  @�?��&�����c�\�>Q�>3w���)��\<Nl���)�   @ǣ�  �n�A� @'sq�:;k�T�I��CCCL6s\��X:m���Tj����/��y��CC֑�b�(�u<�������Wv��H  �Ɏ�ٟi�ߴ��c�dR###�1z��ܫ���̹x�؂���T�   ��Pp  @7x����!�N�bA����m3&�
���7!��E*�y�u��	������^���݊g�֑�f��k�=���������շ{�u$  �,�����Tun�:Ɏ�r9��y�=��{��i��(�W�K��   ��Pp  @7��Z�:�e��p�r��}};z�T*����&%B�+�}�u���P�=��^������_�B�:�m�?�Y=�#Qfl�:  h���I=���Y�h���!�{l'�N�t����%g�x�آ_���   �h�  ��n�t�u����q��{荒��̄���m���05>>.oρޒ߿_�n�	����/�+>�y���)�p�����y�����}N���*�D @כ�����/}�:Ǝy����Q�ah�'EM���[U(�Sp�.��A�   ���׀   @���x�
\���*�ܷ��}���+�51���H(��u�-)�t��������Uzh�::\,�t�ޠ���E����s��0  zɁO|�'�TA���1'OZo�0�������̌ԇ�zL    IDAThX�0E�ؔ7IbR    :GK   ���Hz�:���8u�	*33�̄�¶�wxxX�D��i�+��:¦$K%����?�c�n��:�L<��m�����g4��gY�  �T�������u��H&����{<O�N�f�JE����(�����~�   ��Pp  @'��$�i���E����m.����+��59zEᮻ��f�0�Ϳ�Kz�_���{�&pcG
7ܠ{>�)��ۿ�;   ЕN~�˚���c4E>��Z����nW�v��ce�6����u   �RX	  @���:�@7pu�{��{��E�x<�!J���X2��^`�����O�T���
�����}������K�����4 @�i4t����$M�n[���̸��D�؂~I�   \
�6   �T���t����KK�1�lu
],����|ʛ���}�YG�@�H��w�[�~�����g=����=�� �u~XS_��u���}_ccc��b�Qz�vN�k�O[G0��2`�+)�   <+�   �DiIo�t�*���L����?22�(b�
W���d��1$I#��������6�g<C/���U���݊�; ��q��_�z�:FSDQ���a�=��	�.�z'���!�MÒ�d   x2V  Љ�!ik�M�a..ڕ���#����b������A/��P/~�i�0���?����~O��,p����u�g>��7X�  ��|�N���e�i�٬
Oo&�'��~���a�}@�g   8_`    x_�;�C ���E��ܜu3��+��6��d2�R���D�5���Ӊ�����t=��U�����g�_{����?���G��?�鞙
�S<O���.��y
2�s_��"����l��<n��L�;F}}jl3j}uU�J��ժ��˗����Ը�k�����瞻\^�ZM��e��PuaA�T=���%5j�m���p���Hw�}���n688���U-_��	lN�p��B��:�m���
I_�   �E�   ��%�t�*o������q>�i||��"���ݦh`@婩�����io~�����\�\
��z��ަ�3��o��Z�������>�ɤbɤb����>�R��K"!?����ףH^ɏ��G�bg�K&��bɤ�)H�%�?�5���cv���r|�R9W�_ZR��X/�k�Xߨ�U]^V�ZU}mM�rY��5�VVT[ZRuiI���WWU]XPmy����T1 Zm��?���������Q���<��������q�ҶEŢu3�܃ PE*�wb ����(�  ��Pp  @�y�u ��Ppw�f'Ѝ��)�D���t�:�g֖�K��j�G?��-������~�s���~V��o�����i���(Z/����TJA*%�l9�LQ=�J)�ɜ�?�T��l|��:���V�����ᗗU]\T}ee��_[YQua��}g����������_0� ��؟�y��%)C�������jp�ж}}��P�K���ʎܥ�]�(�[�_��%}�:    Qp  @g�Wҭ�!�n�L&�#����(���c�N�ې��t�}m)���ɟ�s>�!��b��LFw��oi�����ߩցE?�d�뗾���K%E���)<�1���(���s�Hn�=�����6��g�W��U[X��ku~~��kezZ�z�	" �b������J��m�iR��t��)�(�����Zsp'�z���ҒbH�R�����t�J��   �D�   ��_Z �����Y�f�6�=�N���6�h���oVr�.�<�DK�ߋ�t�;ޡ�|�%���u<���7�����k���Q�0�W��)�f�f7
�a.w��~�%�f�..����Ri[�ۨV7J��'���T��UuvV�UgfT��Uev���@7k4t��7]��X'i���-//kii�:JW
'�������]<^4�+$]'�1�     w   t��Kz�u���`���+�c��FGGۘ=��Tz�Ku�S�j�S��y��i�9�i�s�P����g>�o��o����}��٬���KNS?{��D�h`@�6�)�����BA��ɁOvvR|uaA�)�O��������˧OK�F�� ��䗿���z��X�:JS�������V��Q�N��zIezZ�]��c�q�x���Hz�u   ��;   :ůk��)�-J$����	�����ollLA�G}4���_����4��W�����+��i�@'��@��A���O��|E���m���
��(��W��+*d��ql�٩�Q��Ծ}W}|�\ޘ�^��Y�?;����*�:����zI~zZ��5��6�) wU��5�侮�u��:{2��Ç��t��������LQp����>$�u   ��Uo   t�QIX� ��kv��U�VV�c����b����[���cc��z�����<��?�sz֯��baؔ������b��P^,&?��?֧��7a��o{����5:v��V'�Q���⃃Wp��^|?}z}���*gJ�k�N�r�}���ևzԩ���+�KR:�V�X�����"��#��Pp�� t����H���A   �6
�   ���t+��\��.]���L&Ub"6Z`��/�q���}���w�lR*`�/��-�_�����/����g�9rD�J�����ߘ5��e�MN�2=�^�?[�?{����ɓ�-/�!8�]����+�=xbe�T���V>�{����T)�[G ��/K�-Ik�A   �.
�   ����F�@�
�@a.�_Ief�:���I��|���証�&
�2p�=:�����wM�I������_��d��Xl��~��~������H$�w�^=��Ze�2�&��RJ��+��{��Ֆ��v��&'U>uJk'N�=S�/�:��	�pOuqQ���=9���<���jbbB�Z�:NW��.h.Xs���H$�# ݬ��u�?4�   �Qp  ���K�t+�\.����'�>22�(������_�r������&�E���P�Z�=�������"{��}��@{���ѣG���h�#b�R��)�o�eS_[[/�OM]X�?qBk�N�|fR|�^ocr��N��=Yp��(�4<<��G�ZG�
.�+�ܙ��دI����u   ���;   ���: ��\\�sy�{�������f�Fi���W�Z���/����3s��酟��2��-L���y��ϻ�Qj�ŬSn����ɓ'5��W :��+�{���w_�1�jUk�Ni��������Z=s}��q�?�z�������~�[�Z*��jqqQsss�Q:^��ȏ"'�Qpw��dO�t����   7Qp  �����AR ���b�����sQihh�0\�ڷO��P����M=~���O���������й<O~�+�?�k�ۇ$=����b������� ��xA��Ȉ##�}Lezz��~���z���W��ۘ����ǵz����QZfxxX���Z[[����<OQ���'���]muU���<v$�y�h�!
�   0�۫I   �t� t;�*����Dg&�{����1��o�����w��׿.��W|�ೞ�~�
S�6%�	�[/�G����*�J�}_����Q �)�BAa����o���������ǎi�����ǵz��V�U�I�h���~W#=\p�}_ccc���P�*��]:Zp��ON���Y�0��13��t���   ���   +O�t�u�۹�X����L�}ppP�D�8\���������_��e3��^𻿫X<��dh	��(�o�ϟ�N�}ӊŢ|��	GU �K����Z������W�v�V���ѣZ;vl���v����r������?j��c�T<W�T�ɓ'��t����\S��V��;���$�_�[��   �=�F  ��$1z�!K�.ܣbQ�LF��ag���N�����%�Q������W,��a[<O^�?;�=�֯����P�<�=#����}?~\�F�: �	2Oy��Oy�%���k���.e����`B5�h�ᇭ#�E�P��⢖����t����Е�i�f(�M�:I�R���P   `��;   ,Hz�u��R)�mW����`&Q,jdd�:d2���#�����>=�#��%��xA�1}��;S��.����}=z��; \F��*��*s��W_[��#Zy≍��#Z}�	��<I���z�*��
��������8�Z�f�#�Ţu3e
� v.!��~�:   ��J   ,�O+@�6�����z�l��ص�*��
C��P��~��}����]w߭���<�MY���¾Q^���R;��t���>���Qr�m��q���V�k���z��>����������'$���j4���#���o��� ��Ȉ�9b�#9=���]�(�M�+�>.�j   �`U   �J�%�@�p�����lZRq����y�����)��뎏}�u;��Fyݏ�/(��w�����Ȉ�;f z�EJ]s�R�\s�}�J����Oh��!-OL�<9i����9Qp���g�r9���YG�8�������̸v�h�QI?/�O��   ��  �n��4l��M����ZG0H��}���9�0�s��5��B�<�wn�y���(���=%�˩�h�����Q ���a��޽J��{�}��e-OLh��!-<��C��/�;�kT�Y>x�:B[kyyY�J�:JG��E�f\���0���<�w   ��c   h�wY zI*����VUGf����X�:
�d2�ݻwK��VR����x���x|��~f������M���U��u��I�( �X*���nR�M7]xG���cǴ<1qA�}��AgO��f+����}����СC�Q:J,�V,Wmm�:J�U���#�J&�܁�M��$}�:   �@�   ��<Iϴ�׶[.;Xp��XG6���K�����Z9|���%xaxa���WNT�Y�BA�ZMSSS�Q  ��}%�ǕW��;/��:7�>�}bBˇ�����ѣj�jF�q%�R��ԉ��TJ�bQ�O����Q�|^�'�c�]uiI��5��u�DB����1�^�^I�`   n��  �vz�u ��$�I�m����PR��u
�0E�������g�Q��޽Zy�	�WW���g�:T����J%�j5�8x t� �S��[���n�W*Z}�	�LLh�l~bB+����d��T[^VyfFQ�`��J��������	�y�����>�=>2bÄk�!�6�YIC�؎   -G�   �2 �~�@�qm�Υ��'�p��w؊�bڵk����CI^(�g��N�Pun� ]x����ϿD�S�@�CCC�T*Z\\�� �&?�ڷO�}�T|�}�S��|�\�h��Ǵt� ��6*�<�\���<���jbbB�F�:NG��y�f��S��u��D��!���A   ��(�  �]�+ɭ&.��-��ly�rZ_1:��;�x��]�v)���?���U%��ډR��Ƅ��E�b�x\�3Ev/��Ȏ��<Occc:t�V]�	 z\T*)*����ܾz��z���ǵ��c��P�\6Jڻ�&'���F�m�H$T*�499i�#�ܫx2�v>��-�>*�j   ���;   �!��F�@/rm�Ε�{\R�I�Qp�����M��	s9��N�Tu~���v(�(�����Tv�����A��k׮]���P�R�� h��Ȉ##*�qǹ�u�9r�����Zz�q�>�F��v�O���`�X,jqqQ����Q̹\pwi7�'s��&��^)�ϭ�   ��Qp  @;���1�@/J$����EY_RAғgESp����A�r�-}�J����ϫ|�j�eϓE��0��<I%�z�  ��Wr�n%w�^�⍛땊V&&�|�}T�h�Ǵz��h����FFFt��A��_���u3���v�h�_w   �w   ��;� ���<�&Q���T[]���rY]��z�Tjw8���_�bq��K��ܳG��e���U[\ly������<�ɧ� �)�kllLO<�u @��P��W���Uz�K6n�--i���/?��}Tˏ=f�a�����Z,�"�J%�tx��$E���̸0,�r\:n��~I�H��u   �.
�   h�[%=�:Ћ⎕6�ss�Z..)s�����vJ$j�s�R)%S)5�UU��U[\\/]���E�bg�쉄b����C]�~�LF����� �p�tZ�[nQ��[���hh��1-���Z~�1-��?��׿n�T�#�+
ZXXв�'?��u3.Op����{%��:   z�~   h��Ir����k�t�/�{���/L�S��I��V�b1�������>��
�PP�VSmeE����K��F��F�z�7���XL~��ϛ���bM�t������jqq�:
 ��x�ccJ��I/z�$�{�y��}�8��'��522���^�[G1��K���]�:���/H�5I�E  ����  �V�Kz�u�W%	�m���9I�e�s9�����kttTa�޼XLA&#e.�gA�^�<ϩ]*��y����QMLL�\.[� t����)��'�c����XG�Qi``@����QLxA���OOx���)WB�h����J��    �M��   \譒��!�^��"]//�F�.]�=s��@���q����\�t�N��Sn��b����ƚ�� �=��y�uS��B��ܱ����u�rY��e�&\x���   -��   Z���^�ڢt�G����JmJ�����X,Z� p�D"���a� �.���Z��u3�J�:B�8�K��'����u3���&R��u��]+��   �M�  �*wK��:��\+�W��#�DVRx��D���bAhdd�:�K��r��r�1  ]̋�w��)&�_ �"8�K��ܥ���J\;vy�u    �&
�   h�wX z�k�t�,����6�����gttT�X�:��VE�1  ],���'���h4�#t�b��D"a����~�fzuW��q��`�e�ƬC   ��Pp  @+�~P@���k��<I�3_�&*�Z�.+�J���1 \�����m�_  .�r�=��g���<���Q�`�Lef�:�	׎�FI�l   ���;   Z�]�X= Z̵)T��y�M�'i��x�b��Q�D"�'P ]!�L�ȿ �m���:�?��Б��s�-�|�:��^�Y�;�Y[  ��(�  ��<Io����)T�F��cCI�-<�	�h&B�g``�� `[������}vު���: ���x<.ߧ������C   ���i   ��rI{�C .p��V]XP�^���4y���Y��@���a���N�Y�^�y�FGG)�  ���r������y�����c�M�r�}f�:�	��{�u    �VB   �l�b p�S��4����zE�ض�h�d2���~� �!�"p� `������Pp��T*�\.g�-b��0��a��	�[�� c/���:   zw   4�.I/��"�JYGh��ܜu���I�j�8��ϴ14��y��me ��P(P� lImi�:�>O]��Аb��u���<��Nq���|I�  ��A�   ��I�u�.m��+����A���h���řb	t5��4<<̉* ��i4T]X�Na&��g���b�������j���1LPp����"�   ��  �,���Z� \�R��&�%$���}Q���(pX<W��&���H$T(�c  �@yjJ�r�:���/7%��)��Χ���j�]�*33�LPpڪ(��!   �(�  �Y^!i�u�%.-�U�|��'i�K���@3��q###L|zH�TbG �U�=j���6oxxX�����N�{`x�v�t��o�   ����G(   �No� �&�JYGh�n/��I
���Ӷ�$�|��}��x����!� �G����fEQ��;>Eܫ���]4vC=    IDAT��Z�   @���  �f�t�u�5.-�u�@Rv�R�@�b1�J%� Z �N����: ���^p�ZG�*�b��w�	.�Wff�#�p���!|I�b   ݏ�;   ���"��K|�W��1ڦ�����|T(4+
600�X,f@���v� ���9b�ܷ��<[�h���{�	
7H�@   v��;   ���� ׸�8׭����νsy��E���=-�"8!
 p����Q���N�,�J)��Y�h	�O"w���H$�# .��S�!   ��(�  `��t�u�5�T�:B�4*U���clYLR�',��,p�����(� �ӨV���c�1̄ehh�'w�
��������XG0�ڐ����u    t7
�   �)R\�>խƲj·���؁t:�L&c@���R�d �a�T�\��a&>8h�k�b��|oᅡ����[���w�̽�ƬC   �{Qp  �N�%��:�"�
���y�[IJ7�y<�W����ع��!� �(��)�[�  t����:�������Z>���rp�ߌ�ֺ��w���&&��!   н(�  `'�,��V��.���\7��%5c�� ��׃[£=(���<�''� �o���:���޽��^/�4:Zp��˪-/[�h;����Ԝä   pw   �ă� W��8�m���fU��|�I�XG `���ϩ�	 �+s}�{r��]/�L*��Y�h*W�T�����v�7L�t�u   t'
�   خ�$=�:�*��*]Tp�%5s�?*��lpI��(���S� �Ԩմ���1LQpo���A�zhw1��ڎ�� so�   ��D�   ��v� ��\*�w����f.���b���<OE~v �e2%�I�  c�?��j++�1�x������1zB=�C�����w��^!��_�   �6
�   ؎P��Z� \����n)���2M~Έ�2���� $�� ����:������ ���3��|��r��{��Tff�#�]���],!�u�!   �}(�  `;^%�w�6]ȥŹJ���%yM~�0�o�3��1��Y�t�i� �y���={�#���4<<l�)\��^qp�{<��S� ���:    ���   �o� �.�HXGh��u��Ji}Q�E�B��,��*C� :'� ���=��u
S�k����sR���٬u����������lI7Y�   @w��  �����! ׹Tp��	�֧��BH1[T� ����sj� �9��:7g�T�O��Г�~�����&\:�t�7[   @w��   ��VI���9�0�h����>I�=7ܱ�tڝ� 6-��[G  �����#���F�=)î�%�O&�;:���	�C�р��:��0*   zw   l�� �3�Xk++j�j�1.+�z��e�O)[��v ���߯ �c  �l������LF��1�=�P((�򂸫S�]-��r�pC�~�:   �w   lų%��3�\�<U����pE9I^�?��xh�x<�L&c@�<O��� �Y��f��]��27�(y����6��U*��c숫�z����u��K&�� �{�u    t
�   ؊_� `�+����u�ˊ$�Z��A&����:����|>/�� 8c��U���R�y*�Z-��*�j���
-�KR�Ç	�܁��RIlY	  �M��  �͊$��u �\)�wr)��K�!�elR,S6�����A��	 p����e�\���#8app�:¶�:�]����Z���h@�Kz�:   �w   l�+�d�c��0W]X��pII��ƴRT,���+�٬|�C< ���� �f��;��$�Lv�ItA.g�w �^o    ݁�O   l����\'Np������9��Ci�f�R)��>= `�:7��G��a*�d����R�$��cl������z���C   ��Qp  �f�%��:�s\)�u������
mxt�d2�B=�M�9<� \1��H��uS}�x�<v8j�(�T��ϯ.�;q�@��r�"o�   ����   lƃ�X :DE�Y��m�}I��|=*��J�fLo����]9a �y����us�g>�:�s�Ŭcl���;���t��h}�L   ��hD   `�^k �9.-�u�����A�	����Ͷ� � �����: �Eժ����c���z�u�������[B��-.K��nIwX�   @g��  ���V�m�! ��ҶʕZt$e��z�q5�l֙� 4O.���  h���}O��y���(R��7[�pR>�����>y�~�r��w�#��:    :����  �o����Ң\'Mpϩ���Ƌ�6����lG:�V�1  -p�k_��`.s�M��:��<�S�T���i��)p�ĿN&�..K���J�3�   �v�   p5�� �B�,�5�..Z����Ғj�k2�W�ŔJ���@/�<O�L;�$ ���o|�:���3�i�i}}}J���16-�﷎`�2;k��9�t���WX�   @�bT   ��NI�Y� p!W媋�R�nC��jK�������[d�Yy^;� �K�٬f,6�}�kk����Q�����F��ڙ���S]Z�j5�VWU/�ըTT_]U�V[���8�=��j\�}au~�ү���z�r��jU���n�|_�M���Ӓnf��HlL���w�O$��E���|��'���XL�TJ^*�Lʏ��G��dR��� 6k��?�ڱc�1�eo��:��u��A���j��^.���*ߑ�K�;�Ҁ.�FIa   ���;   ��M� \̕E����-�������%(�2�٬u ],�J)U�U�(���yՖ�U[YY�,.���������UՖ�T]\\����������WW;�=\/����%�dRA_�z	>�T,�T�ͮ��I�����s��׷~�d6���z��׾f���Sp� �DB}}}Z8sBS's��.���9r|Ir�XЅ^"� i�:   :w   \N(駭C �X<��J���,��GŢ���[A�d2i@�<O}}}������&iT���ϫ�������/.RH�`��%Ֆ���\�t���{,�Q������\N��K��)��W�Iu]c����:����7���s���Z\\T�Ѱ�rEA��g���)���6܁�Jz���d   ���;   .��hXȕE�N([�����n��S�pu�lVSX�P6���ޡ�kk��Ϊ:7�����+����Ϊ<=��쬪�����ʊult��e��-~�����lVA.���� �߯h`@a>��XTX,**��L�7�|�{�:����>�:Έ�H�lVsss�Q���	��9��C��+�Ҁ.�ZQp  �%Pp  ���: �Kse�{͸���fz���bp�L�:��L&��T�լ����ښ*�O�<5����*33�3������(���4�����M����{�TRp� l��bq�v��M3��k�#Pp�,�RI���=���{'h'
�@G�]�.IOX  @g��  �KIH��:�KseQ�b�ؚ�݇f��qe��+�ri��V�<O�L��'�v�z}��>=��S�T��^/��>�q��}��%�@���������W|��)��
���B���RI��!Ň���b�6��ө�|�:��X*��ӟn�	�P�|^����Q.+�Y��n���{�0������u �%�^�Ǭ�   ��Pp  ���J�a��J��r��/)k��Z�f	\B:��ǤS M�N�)�?Y�����*�:��SZ=yr����e��̌��i�j���?������(VbhHQ������
K���Ţ<�o_��|�����a.w�m��=;�������:v��O.�8�0�Hhyy�:�K�yQp  ��p�   ���  ./�[Gh���kg$YΈ^dǕ��i� zH&��9���5�MN�|��N�\/�NNjmrRk�N�|�ʧO�Q�ZGp�z}����.�	�E������z48��X�z�DA����?���p	�XL�|^SSS�Q.)���/4�Q�ε	�w��=C�S%��:   :w   <Y��Y� py�Lp7Zl������q9��Q�V,S"����u���׵65���ǵv��N�\�z�V���䤓E.��ju��~��K>Ə"Ň��W|tT���.A��Ϛ��.I��ޱ�Ţfff:r���
�IU,=�:�@G{��Y�   @��  �'{���u ��ʂ�����K��K���
��:���d���^[^�(���8�ճ׏_/�ON2y���e�>��Ç/y��^T~O���tޒ����	��##J]s�u\����ɓ'��\R��9Ypw��?W��]�բ�  ��t��8   X�y�  �̕���|�_3&)��W��q)�t'�t�5�LFSSS�1�z]�'Oj��Q�=�գG�r�V�\���Z'����Zx�-<���w�����e�3��]J�ޭ��݊%m�L���a򺝦p��p������V�R��r� ������v�\��r<�b�Jz���Y  @g��  ��$�*t8�����N��.1��F�@+$	���z���ת..n�W���c����U��� HZ?	��1�;vɻ��A����(�'��Ur�n%FG��b-�t�o��5��e�w�eWqv���,�٬u��U�������Q�ƅ�i@xP�  pw   ��%��! \�rՅ��h�kv��vI
���KHM��<�S2����RS��:?�QZ_��$v �E��I�''5��p��^(>4�>�}|\�k�Q��k�SbtT�m���w��r'��a,�L���϶��M��r:}����u����u3��yE��u���;T����Iz���  @G��  ���: ��s��^[\l�kf%m�^�<^,� ������k��O ��J��^.k��!�>|Qy}��	5�����ѨV7~G�~���K��ܳG�k�U�k�ڷO�}��T�}���U��J�s�+?��c`<�S�X�)�1G'�KRev֩�;'�]aD�]��n   �(�  �qI�[� pu.L������Q����w4����x ��J�.��:?���t��F9s��-OLH�z�C@��--i�G���#��vm�Sg.ɽ{���$�����_��A��S|��#`r�����T�T��l.�W��#���Ӏ�zQp  �(�  ���J�C �:&�W��z�2�]���~��@�*��N5�u���[Y��?�C-:��C��|�ꫫ�� �I�Je���4u��dRɽ{�ڷO�T[^�	�A<�W��;�c`�Nq?q�u�wg�p<�?-��8�  �q�  p�+� ��0���.J���;iz�tf�;�$Lp�m��ꕊ����emM�3�������5����g�N��8����Nw�����H��D��L��.˒l˒�<�|���T���}�d��̋d�T���IR�7��U7sS�Ln���)O%�;q2�܉�+o���"%R�A �z��}_ �H �s��~��
��ϏZ�������2 p'�ZM�o��ŷ�6%1��Snd�tl��ࠦ��3�=[���`Lkv�t�X1�H�ݒ>-����   �,
�   ����N�`c�L�j�XpO��vI�����	�@�\�t )��
uE+��FC
7|���q
� �Ty�9��I���ww�rM���E�  �y�   I�&���Ѐ\Y��k�{Ҧ�KLp��\�����Ⱦ�����bB  zo��J����	�ss�#Ċsk U�"������\   �w   H�WM �9�,��Up�W���KR@��6ꀻV����{�l�Ⱦ������1 �ґ#*NL���mJ�w�X���*L@�>nm
� �k���%���    0��;   �I:i:��qe1�C�ݗ���W�:&���(���"u�u���
�uE�vl/?x�2����y  �m��ϛ��J���5��Mǈ]{~�t�X�rM���E�  �i��    0��Z�yHW��qLpO��vI�����a�[�VS��-�>��ٳjMM���k�]��|^����  l��sϙ���1�=	�J�t#Z�Mpw�`�WD�	  �i�  �WM �y�]�==~R��KLpǭ2��r��� �,
C��_W���K�ׯ�^h_��=���  ������Q�1�����f��c(;0`:��ZMQ&�ǥX,�� `k�Jz�t   �C�  �m�$=b:��se�T��I��.1����r�d��_+����P͙UϜQ������H���n�  ����ϛ��.I�wW�Ԛ�5!6�\S,�    s(�  ���Zd %\�6E���jώ�K*���;����X�+�6 ֋���gΨy�j"����B� ��?�Y��E���
��h������#Ć�k �����)  @�Qp  pۯ� `k\�6.-Iaس㗕�a&��f�\�t ;6��;�ƕ+�-��001a:  wT<p@}��o:�(��hxx�h���	��$ܨ�'M�   �I^�  @o�Hz�t [�B����سc{��{v����ey٬�H�,�= �֜�R���j��lJ�ؘ�a8  �v����聡�!���M&].�7ggMG�M�w �-_3    fPp  p��&�+�@ʸ0m����Oo4	C�H���Q��y5�]���t�M��yOP �N��������4h�|8�T���i�&�Kn� ,���    0#���   譯� `�\X��������ד#wOvh�t$w }�fSճg{��Y������  ���x@��q�1�#����<3K�.OpoQp�|�>a:   �G�  �M}��6���r9�z���Г���m+(��f�L��Ӂ�	�ΝS�l���me
� �����K�#��� Ѐ��y��	�T.\W,�5�   ?
�   n�I�! l���z5�'G��-ّ<�lV�L�t ��Zno�MG�&� �(������c��FFF������o�kw���z�t    ���3u   ���  �ǅ��v
�EIi���w�,�͚� `��v[���u:���Xy�>�  ��࣏*;<l:z,�˩����陌����_7:�������  �xQp  pON��C ��R�E�=��%&��V܁t��H��Z��tEit�t  n�祗LG@LFFF��n00`�uMkQp�_3    ��  ���$��bX����n��+i@�7�}�t �иrEa�f:F���� �0^���g�51)
*�˱�n�т�k�]X�+�    ^�  ��U� l�q�./��ez�$e��LG@�Pp��������]E� �4#�<#�T2121�=�Tb�$[-�����qap`�OI�g:   �C�  �-I/�`�\(�w���v���b׎�{�.�cm܁d�:�/]2��(� �f��/������e
�X_��	�R�$w �<I�t   ć�;  �[>#i�� �/�^���];V���KR�R!nB�H��Ԕ�v�t��˖J��� ������x�t�w��{gq�t��PpR�WM   @|(�  �嫦 �&�o�/)m���i�䣗(���Zj]�n:F��.x �e��?//�5���+����;��4�݅�j�垒�	+  �#(�  ��� ؾL&c�B\X�+l��r���LW��LF�B܄�;�\��i)�L��<;�  b��/�� C2�����b{=�'��Tpg�;�zYI_2   ��  ���%�c:���f��dRU�޲v����H��ʑ����Ph�M(����j�Κ��SLp $A���?���0hhhH��rv���?��y�bc���_1    ��  ���� `g\�2���԰���U���C���?��    IDAT*r ؚ���VOo�$߁� ��}��`��y��t���j�6�.\[�I��   �=VJ  ����@ʹ0e�[���]9J����1��� �Q��w�y٬�  �y٬�����H����X^'�K�>p���Ұ�4��X�"�i�!   �{�  �0$�� vƅE�n���x+����6
�@���u:�c����Mu �d��g�2	���T.�{�:^���M~��Я�   �ޣ�  ��_���
`�:](��u�w܌r;�L�9�b�j� ����b:ddd$��	�Ӹ�ε��MG���#����    �=
�   nx�t  ;��"\k��@R�;Qb�4	B�H���T�Z5#� &�����c����)�˱����������nziQ(LG �G$�k:   z��;  ��IϚ`�ྱ>Ii�3�7��$�+��%
�  �F_~Y�X�ĭ���z�>ܭ����!�t    �W�   ��yI�! ����¶֓T�^��Qp��(�	Ej9Tp�)�  L�d���_6�	T�T��~O_#p��ީV�(2#.\[�   �Qp  ��WL �.L��,-m�gKJ�I��� ��jUQ�e:  �|���7	�y�{����Ga��w�K
�U�4b:   z'�k�   ؜ϛ �;\X�����/C6��G"G��i����Oi�i6MG  8j��WLG@��t�+W��ήǤ��# �x�^6   �C�  �n�J:d:��pan��
���F�]v`�t$w Y\)��2� `@P�h��L�@�e�Y������A��t��y�b����1_4    �C�  �n_1 @�����f����&0�7��$G�VS�n��+
�  �~�K���;344Գc�Lp�^�<*�E>+�7   ���  ��^4 @��>�=
Cu��-��/���8�����EQD�H���.�f�f�t ��F�l�\.���H�r�ݡ��.� 2$�1�!   ��  �U���� �����Ғ��BoYR��qb�0 ���#�,o�w @�*'N�t���H������傻K�ym��8��   ��  ������ ���	�-�LFR_����/��	�1�0Lp�[-������� �۾�~�t����<����.���m��8���  ,E�  �^_6 @w
v߳ҩն�3I~��Ď��XK��# �s��s����~ �9��A�<���H���߃2z�g�-�����^ۯ�zH�^�!   �}�  ��Y� t����3�ݖ��R1	��tLG �����lИ�3 ���_��<��w�}���]?f&���h���P����k��2�^6   �G�  �N�I7@wپ ��b�0���M��Lp�(��EѶv�Acv�t �C����H�R��|��W�L�O��C�^�w�8v4  �w   ;}�t  �g�ʝjuK����xd���5Pp���뒣�6��MG  8b��I�2)544��c��]��N��ҳZ��   �Pp  ��� �>�'��[(�g$�{%v�N�ÝQp���W�h--)l�L�  8b�W�t�X�R���]=f�����Eۡ����� GHz�t   tw   ��Iz�t �g��V��E�uB�4	D�0�Ղ{cv�t �#���y�Y�1�b��i``���tv�{����4#Lp����    �.��    X��$��*
�#�T{qq�ϵm����y؁�;`VX���`w @\����<�o�F�v��qW�;S�)�����    ��t    t݋� ��'�o�H��}w�d)�c�s�fS���6��LG�+2���e�Y��2�//����+�y���ok�K%yA�L6+�PPf�go�����-�(Z���Y\���_�����ӑ�h�9�Z��V��Q�|#g������QX�)l��?�Z��X%���W�b:,P(T(T�׻r<��{vd�t����X�I{$M�  ���  `�gM ���å�M=���&ܱ��7����te��+�# ��\N~_�����r����������BA^���_�>��+��W(0��&a����T�h�S��������ZM�jU�jU����U���:ժڋ��ϻ���u�UE������'�Pq|�tXbppPW���	�����ఌ�/J���   @�Pp  �˸��M� �}��)�͚��S�ju��d$�z%vܱ
�9����˗MG@��~eT*
*eW>n�:�￥���SJ�o�F�n	�M���o�h��������:��˓恘��Ϳi:,R�T499�0w|�`e��Rpg�;`�E�  ��  ���� ,��t��&&�$����l�b:��j)�"e2��ĭS���`��ŋ�#`�2e���RnxX��e��)�k�G�������y�S���\N�]��۵kK?�ᭅ��Y5�_WkzZ���պ~]͙�ffV��:��.`��'�������x����>�����X.߀N�����Yd:   v��;  �]>o: �ޠ�������X_Ej����� $N)l4L�0�	���J��ݻ\T޳g��Ȉ���˟W�칡!
�芌�);8��ࠊ���E��쬚��j_��\���QsjJ��5�^UsfFQ����H�L��o�������`w
�Lp�w�j{$=(闦�   `�(�  �##�i�! �F�P0���Z����Mm�&`�;��j�(�1[-)M�0�	��V'l��Wn�.eW���޽��ݻM�6tc���h�ϫ95��q횚SSj�|��u��e��v�]_��J�����ee�Y�Z����])��0DpܗE�  �
�  ��a�! ��oQ��\(�����䱍W(ȳ��/�o�� [��#�i4T�~�t�T��[���ޭ��=���{�*72��
�.P00p�rs�n�53���+jMM�~��/�q���W��y�����1�F7���7�a:,V�T455��c}}�x�"o�q���w�z�����C   `�(�  ��K� �����S�!�	.O���(����Y�tI�"�1�+�Qn�.�Ɩ?��S���J�=��3�H�L,��gϺ�	�M5�\Q��U5�\Q}� ߼�k��,O*/�ױ��]y�Ns�QpW&#�TR{q�;�Rĕ����� �	-oz��B  �x�  ���  z�`y	�S������e+��`�Y@��f�tc�Ϟ5��LF�ݻ�߷O�����7�:?:ʮ+@x�����*������̌j/�~��.���~�W�*�tbLe2����}��1����r*�J�np�a#A?w�1��^A�3���A   �3�  ��'�� z���R��1�0!��7	F��������3��2��ܮ]�����R~ttu{~t�;`�����x�۾��j\���J��R|�]����j��Hl�������_4��J�]�/w)Qzt6���(�NxI�  R��;  �^��Í��ŷ;-�f$��;���t$X��TE�d2�� �p��~���;��r*�u�
���Qؿ���e��#0,�N�uך�o�ͩv��j~����?�����߷a�k_��7�a:���/�����N�����X�s�   `�(�  ؁�u��l_|����$/�(�su��E���
���(��VK
C�1�IK����?*���o��{�*����@����+�?��m�[-��(��;�ڹs��;��^7�6���������ۦc�1�穿�_����>���Nka����R��m�%�$阤]��L  ��Qp  �çM �[�/��iJX9�&�.�c�(�����i4�x����Ri��~s����r{����Q�ߣH�+WT��CUϞU��YUϝS��Y5''̈́5(��:����~��LG��*�ʎ
�.����2��8���iy0��m:   ���;  @��H��t ���w_�ݿs�α9�F�t�a�e:�1�g�(�yz}��US��A�TqbBŉ	�&&��5 �H&�¾}*�ۧ����[�juy����k��-�9����~�������}���|��Q�R��\.��6o^ty���Ғ�� �y�B�wn�(�  �w  ������Q �����:܋�2�F�wl��;���׳c}}*8��]w�|��J��p�]*:$�	� ,�J�;vL}ǎ��xgiI�?\.�����+�K��(2�vg��zJG�w�۽�t@����������e���[�z�gl��d��f9�����    �
�   ����  z/�˙��S�uPK1�0���p؜Z�f:������;��� ��¾}��Z��^:t�i� ��\^��ޞ���������ϜQ{n�Pҍ���ա��w���LGVn��8\p��a�6�|��;`�#��K�`:   ���;  @�}�t  �g}�}�o ����|
��@��Q�ٴ�� 	\.�_{�M=�/�U��P��A�Tqbb�c|\N����8�ʉ�<ޜ�V��-����N����vN�PR)�T���_�]_��<�wC��r�m��=���ۋ��#����������t   lw  �t�/�� z�����&��0�]���~���j��;��т{kiIsgά~��<�GG����Tb/<�������r##ʍ�h��GW������������xs��!���]�/�,�P��k;Q�T499��sy��z;�����l V}N�  R��;  @�}QR�t �g{���;ܱ�ZM����c v�"E��F\��/����ݿ��*NL0� R����w������Ǣ0T����;�h����;j����J�k�����_P�}��4:���
�[�v��n�u6 ��1    �G�   ݞ3 @<�٬�=��؄��ʇ
�؄j��pX.*�L�0��/~!Ix�!��5� ��Sq|\��q����Wo\��\x?}Z�3gT�xQ͙�gg6��?�)74��ؘJG���{4p��r�v��-ۖ�fU*��|>�;\pwe����� ��t���L  ��Qp  H��M ��-�������h6�j��
.� ����vI�Z)�'&' �J~lL��1�<���(@��\p�
yA������X�EQp  H%�t    l�I�M� ��N��H�z���J����wlV�V3�Z�阎`D��h���$I��q�i   �k``@�Lf�?�\�2�������:��|�t    lw  ��z�t  �y�TX�*
�կ�|sqb���0���թ� ���	��o���ʟ/Lp  ��}_�����s�ft&��Г��~�   ���  �^�1 @|l�,��XiץiA��H�EG&���:�����_�$�TRnd�p  ��T*[��x�Rp��:���t��   �:
�   ����  �c�d��O3r���;:��l6�l6M� �����?��$�t��    =���'��ڲ���ێ�f�u6 k���    �:
�   �4!�� �c�d�v�����:Quu�۷��4=��(MG�]��u]�IRq|�p  ���<O�[�A�/�t��G:��R���s6_g��gM   �ֹ�   ��L /�'KuW]4��&�c�o��@w�Xp�������  �k��r�GI�-
C����=g�u6 kz�t    lw  �tz�t  �y�-\��:#�
�ف��2�jU��� #\,��������m0	  @o��ey���]�!����a6_g��QIGL�   ��Pp  H�'L /��N��p��{'�./�c{�0Tu� ����(u�G?Z�:O�  X��<�m�<pt��$u8��:�u}�t    l�k�   �t�t ��<oKS�Ҧ�Rpwmz�$[�"����� +�Vp����՘�]��	�  �v�[8w���^\4��(�Nz�t    l��	   {� )c:��ؾ�֩�$9Zpg�;�aaaAQ���Ǳ���?��[����e(	  @<���6=@���A6��t �{�t    lw  �����  �e}�}iIyI�� 0���n�Uu`�x nQ�c:Bl�0ԅ���[�  ���y*or2�_*�8Mr�(��~����K�0   �G�   }�4 @��٬�=�^Z����.O���,,,�� �ǡ����Ǫ��|�@&#���   �Կ��]�q�C����7    �G�   ]vI��t ���j*�a���ؙ��yE�qtׇ�����I���4   ����Wf�{�MNz��wۯ�Xw  ���  �.ϋ�p�sl�*���M�0����8��:���ժ��U\�i$l�u�/��Ǽ|�P  �xy��Ri�}䂾>go lSp`��M   ��Q�  H�O�  ~�/���u��	(�c���MG ��H��ʫ��17w�c� �K6|N���;�Ʌ	�� ��#Z�)   )@�   ]5 @�l/��].�;��9vn~~^a�� e��ɟ����   ���߯�&��}}1�I����=g��6 �ʈAR   �A�   =r�6@�l�*U��%N�lbj��0��t������Wu��Q�c   ���T*m�<GoJ�T��#����� l��   �9�  ��	I�! ���R�lVrt����st�st�����=(����w�i6o{<l��  0�o��]-�3���4    �C�   =>c:  3l�*U�Ė�����U��T��M� ���韮�xD�  8�����z�.-���s6_k��㒘:  ��  ��q� �a�T� 8\�6��lS�l���~��>X�{Lp  ��f��o��Z�h��S�[������ lJNҧL�   ��(�  �� G�:U���_�����Ip边�9�ah:�~��*r�O�d��E�v�I   ��o��r�T�)I�Da�N�j:FOQp����    �w  �t�W��! �a�[__��w&��[�0�����@�Y\p������}o��G��"n�  �٨���1%Iۯ�d�YyU	�aO�   ��q�  �L� fc���<�J%�L;�izzZ��[�ؾS���:����w  ��b�(�����O��jA�� ���$�{�;  �%(�  �Ó� 0'�˙��u�RI�穵�h:�1�nu��h6�Zr�� ����������w6|^�jŐ   92����Lx�Yہ�56� �iÒ�1   wF�   1 �96.��X@va"�z\���133c:�jK���韪1;����  \t�����y{ہ�5�|�t f=k:    ;  @���I�Ӭ.�;0l=.ou��XZZR�^7H/�Q����6�ܐ�;  pP__ߺ7:�<�݅�A�� �,vN  H8
�   ���$�t ��r9���P(���;ժ�4������S܁��x�]*��?��>�pS����  H��TZ�����v&��v����4    wfߪ  �}�2 �Y�Mp�y��6܁����W��2H''�����ݦ��N  ����3�����Ё�����'��?�  R��;  @�=b:  �l.��\�syz'�"MMM����m�/���z��M?�����4   ɵ^��+�{��Y.$��z�-���  @��yF  �.�M `�M�|�W�X\�څ��O�Co��ͩ�l����e�_~��[z>w  �\.�|>��LF����S����s�Hz�t    �ϮU   ����t f�Tp��T4����#Lq�Ǧ���}M��Ɩ~�����   �Mq�o�I�%mvܳ�z�m{�t    �ϞU   ;=c:  � 0�k>�`:0l=>w���ܜ���@�XRp��H��ַ��s� ������;��Z�@��	�(�    IDAT� $�0    �c�  �^O� �����N��/�<�=Xg:�-Lq�&���#t�����u�ԩ-�\k~�i   ҡX,*�������;���=�w ��I��t   ���;  @�}�t  ��2Q�P(��Xy���D��0��6??�w`l(�Ga�_~����Y&�  �y����鞫wvܳ�z�{�t    ���;  @r�0�y�,�ݶ�w�M�詫W��� �����ǚ{��m�lka��i   ���r�ܽ]�IQd:FO1��

�   	E�   ����  ��e����;����Ҙ��<y���p��Ғ(�����{kiI��ַ���m��   ���~�0Th��`�\o�c��   ��Qp  H�'L �6Lp�<O���]��z=^����)9�199����{@7�����o}K���m�|gq��i   ҧP(���{B�����N�f:BOA`:�dxXt�   �7i   �u�t  �`C��X,��X��傻��T8�W�ͦfvPz\������z�?���	�   ��>��w�݆	� V�$3   ���  �\�M `��yVL����d�B靸�@3����n�M� -������N���c��_�R  ��*}�|�c���(����   �v�  �� �n�! �g��vI*�1���;��0u��5�1�dKi����K�W;>NkfF��.$  H��_��A=���n�@	 ]��    �w  �dzT��V ;bC�=����w��Pp�����:����L&#y�\�i4������+l6�^X�ʱ   �*���r�wx�{���G&���	�   p�t��   ��1� $��mkMo��.��O��Y�/_VĄf`]��Mq�[�����];^sj�k�  H���cx����_�����yP�:   $w  �d���  ���	��ܗ�bN�>�aH���V`]i*�_?uJ���v�����   �n�����N�f:BO�p�@�$�o:   nE�   �>a: �d�a�m݂���w�w�4==�F�a:�Hi)�������O��]=.�  �R��L&#����m����7    ���  �<%Iw� Ҿ]r>�W������wB�&EQ�˗/+�"�Q��IK�����5���]?nkf���  H��T($�}�n�`��_s�u��   �[Qp  H�G%�����O�*�aҙ��`���@\j���_�n:�8�un�J�����Ʒ�ݓc7��{r\  ��)���RIZ���ۯۤ����;a:    nE�   y3 @r�}�T���:KK1&I��	pH���I5�1�DIz�=�t���ծ�{r���TO�  �6��32����0�����~�@�= �;_   ��;  @�|�t  ɑ�iRw,�[����0�IE�.^��(�LG#��_~�ۚz�����;  ��R�����v�ћ�ۖ_�I�57 ]��r�   	A�   y2 @r�y�T6���b��[]߉���H�F��k׮��$����˵_�Bo����5���==>  @Zx�����v�X4��&�p;,  $H�G  �'/���ve2A�V�e:�5�<M�N��%��LpG�LOO�\.���@b'�7��o~SQ��uW����   iR.�U��8z���;�Qp߾ ���$)�ϯ�vpC��R�ӑ�|c=�"'L   �G��b  ����fEjy��Zn,�*
*
��.�*���r�ӫ|�_-_g�Yy��D�Z-�+E�z�.I�t:j6���j�������V�iaa�Y^p_Z�)I���0�.]��ÇW�W%�����O�t�R�_����������  @�W&���Np���$���r��*�����o�\*�n�6\(��n
�t:j�۷\���z����E���kiiIQu�wl�æ   �#��  $�I�`�r��J���h���k�w��r��b�V4���iaaAsss����������477�v��͸���Ŷ�/�މ�ۛ#���.]������<����i�Ip������_c{�������z]��Eu���K���j��+
C�u:
�UE���KK��m����v[�g�FC�7_F����d|_�:��bQ�lV^.'�PP���J˻"��;����LFA�,�X�W((��_*}���@�) ���q]�su���;����fy��J����!��Q�T�u�v�|ߗ�����T*>?��k�7_���������f��$e$qw  @��  �.�M@�y����!�ݻW�������e�$���ڳg���ٳ�����t��U���hfff��6M�I�b�f�:پPz'LpG-..jjjJ�v�20��	)�_?uJ?��ߋ�5�/�|�h���Ya���쬚ׯ�9=���Z��j�Ϊ15����G%����YZR�������岂����~e+���
�����GvhH��Aeؽ �5�(�w���NGQ����v'Y&�����X�^1��kddd�cϞ=ڽ{wjw��<O���\��KKK�����̌&''u��U]�~}u7Q`��%����    ��  �4��t	�@{�������E�RQ&�1-�rY���ÇWk6����ֵk�t��]�tI���S�LZ��M�].��:��w��5
������	i�I�qk�������R�^��u/_���$)
C�ffԸzU��I5o|�vM�+WԜ�Rsz�����j˓�gf���A�����j�=;<���!�FF�۵K�ݻ�۵K^�S> H���.*�jW��ZZp��w�Lc�=��ittT���Ӿ}��{��M]��I�\V�\�����c�v[��Ӻz��._���/j~~�`J��IQp  H�t6%   씑t��H�R����Q���illL{�����[�r��ŝ�~X�T�Vu��MNN�ҥK�x�bj��Zp/nb��咚��ߐ�.]���7܅�U&�Fa����h����_�ޣ�{{~^�T;~��~�W��95������bc�9��椳g7|n00�\x_)��w�Vn���Sᮻ��} �*�b����ZMZg���r]�\.�9���<�3+qn�ٻw�mׅ/]��K�.��ի��.c>%�L�    w  �$9*i�t$K>���Ą&&&��~U*ӑR�T*�2��nkrrRgϞչs�499�(��\[Z��f��"���ʣ8��t:�x�&&&X0��2٬�z�_�k]�����N
�Q��ڹsZ:sF�>P��2{�ɉVh�ϫ=?����4�*�o�
��}�yll�?6&߱� �ts}�{'�݄�M�{����y�������W��H���u�K�.��ٳ:{��f����	�   �,�M	   ;=b: �addD��������O��� X�x��O�V�����:����}---���*�w��������N����sx�ң^��ʕ+3��g���������?0���+W6~R�q��O�V��-�|��=��l�HkvV��Y-������Ua���SqbB��U�� @�����3Il/�'�ׄ�����5>>�g�yF�jU�Ν�|��gϪ�l���4    ˒s�  ���� t��!:tH�p�5��X,��ѣ:z����y]�zUgϞ��ӧ555e4[��6k3���ZI����H���9��y������*c��ޙw����M���2kMpoLNj�7�?�|S�o��N�j lpc
�ҩS�}���T:xPŉ	��U:tH��	'&�s� 0�oh�tcl�~c��������w��5a�J���;�cǎ)C]�xQ|���{�=-,,��3�$I�n:  ���ה   ��:���=�ܣ#G�(�˙���LF�����?���y����z뭷499{�4܋�غ������;RdrrRA�R����&��y�����7Sm�����f~�U�{o���0�n
�M-�:��5����{U��P�������*=��ࠁ�  ��)�[+��n��ittTG�ս�޻�kh���y:p��8�g�yF333z뭷���o'j�O�\Fҧ$}�t   ץ�)  `��M@oy������رc��Sd``@Ǐ����533�S�N�ԩS������m-�۾@z'LE�\�|YA���p�g��ުV����U�P$�"��w����mW��q��f_}����{��|���>��W}�ޫ�訡�  ���`L�^7����vs���ѣLjO���a=���zꩧt��e���{:u�ew7�w   ��ה   �Ӱ�}�C�7FGG����{�Q>�7;0<<��\�?���]��7�|S���=\�K[�=�ɨP(l��w 5�(�ŋu��An΂2�/y����^�n�~��u}��� 6v��>���XP����{�w�}˟�Sq|�`J @�����I���a���ܳ=��uxxX=����>&��\&���ؘ�����OZ�ϟ�o��3g�(���c�e  �HWS  �^'���!,���t��ꡇҞ={L�A�޽[�>��>��O�̙3z�7t��yEQ���I[�=�����׮VcH�L>��H�N��?�PLݟK�vx�\le�������~�k�h��i��Wo���V��	|��?����2�� 6���)'����lP��~׏w��=���:p��2�װ��y�����Ą��N�:��^{M��Ӧ����q   X�  H���;��ٳ:�������n1<;;�7�xCo����]*p��H�ىT�O �o�$j�Z:����ǻ^ �&��J1�]����t�?���� �53���}OS�����
�'Oj��1� �T~�L��Rݺ~;<<���_>��v6����z�!=��C����/�K����j�ۦ�a�J�n�  ��jJ   ����}A��������5<<l:��O?�'�|R�O����s]�|yGǴ��n���,t"����j�}3�5 i�e����5���?ԛ�����U ��������=�<��o|C�O~�t4 @�d|_�BA�ެY�{��u7��t��w�ĉ�b*�ў={���~VO=���x����kZ\\4�W�tD�{��   �,]M	   {��a
�J%=���:~�8�yp��V��ONN��^�;Ｃ0���[�LpҫV��l��y=މ����~�/�EO_���f_}U����ܮ]|�UyDC�>�<�5 ��b��?IӶ�����n�\N<��>��Oj``���f�BA'O�ԉ't��i���?�իWM���w   ��Ք   ��=�`�u��q=����+#~{���/���{L�����x��Z�M�|���}_�|~S��T�=N�\�&o �liiI.\����)��J��?���Y?�g��g��3ͩ)M�ٟi���L��w�F�W����J�� LɖJ
ff�6$f�(��u7��`+n�r��%��'?�|�(�LG��}R�wL�   pYz�   �: i�tll���:y�&&&(�a�*��>����G�믿��^{M�ZmßKS�}+�{�/�މ�"(,�����/ꮻ���EX���zr�����G��+�Ʈ. �X|�m�~�m}�/���|�K�C�]�L� �,(����+�o��U�m���ȈN�<�{�W��Ő
���/����)���?ջﾻ��>�M   p]z�   �:a: �l߾}z�'4>>n:
,P,��c��ĉ��/~����j4�>?M��&�w,_ ��	���.]����1J�J/&����?���?P��t�� z������G����j�k_Ӂ_�u�c b���Krm?����o�wx�?00�GyD<� �vtŮ]��/|AO<�~����7ߤ�l�L   p]z�   ���� Xۮ]��裏��ѣ���B�lV'O���?��_}ݢ��ڒ����xLp�e��������O���x�2A��ݝ�������D��@X��¿������#��[���K�# b�LpwMd�|����X�}�Q��虁�}����'?�I��G?�{ｧ(�L���I�KZ:   z��;  �y���[������=��CQ=���t��I=���z������L�fs��k-�%Ua�����;a�;l����?�P�  kd�ٮ�O}�;�����"&�Vi����o~S������{�i� `9�XTV�'ɥwu�(�y�D__�N�<��z(U��^���������)���ݓ������M  pw   ���0!*���z�)��0�P(�����?�W_}U�����0T��-��m)���w�wتZ������a/�U�ÿ����ٻ��8����OU7@c%A�$���H��(J�$j�D��,ْ'V<��ؙ$g�8v$'���M�Q6*���ڞ��3�=�NNb'�8�sm�VdǋƖ-J�@�;[�F7����H���4��~����spD��>�����~��?��SEJ��z����ڿ_�>�	�o�� *U4�#�J�囯��hT��պ馛�m�6��b��z��t��}�;���ӧmG�w   k�є   �\��5�C�]UU����z�p�\Āu�x\w�y��mۦ�|�;WL��Lo�4��`�E(������K������sc�Y?����ɟh��?_�D �j��i����?�#Ϳ��q  %��%���n�y�\NN@�Ö́1FMMM��_��/��lZ�d�}�Quuu�[������lG���v   �0c�  �]k%��V��hӦM��>�]�vQă�̛7O�x�;t��)��^]]=�Ǉy�{���v��FGGu��1e�Y�Q�9�m�'���{����ہ�ɧ�z�7S}����( �p/������)�TJ����ZZZ(��w�����Oh��݊���k�f�   �;  �]�l�ŋ��Gս���E����^}�U?~\����Lj��+��h�\&�#�٬�;�t:m;
0k���>64�o}��:���W	�;/�ӫ��[��mG Y��	�aSI��������K�x��F�s�N=��ڲe�Ǳ)���   fQ�   B��eV__��o�]�ׯ�(�1F===���W[[�.\h;�[̸�^AGg��;�"������jkkScc��8��ʹ�>|������h���%^6�W?�qm��C5mm��  ����*I�$c5MyUc�N�>���ny�g;P���z�}��ڸq���o����v��Y.�FR�  �  ��v��pG�6m��?N��5>>��Ǐ�������b4U4:���+i��LE.\���S�N����v`ƜhTr;}z��W�����r; IR��O���o��x& ��\<�w�	rAR�J���~�={�r;���M�}�{u�w��*�{IX�J�`;  @XQp  ���u477�]�z����O��hxxX���שS�d���a��w����_nLpG����̙3����D!S�_�����}������!��H�߯����ڎ (�H]ݥ_�l���ꐂ���<x�W�"��r]W۷o��?�+V؎&[m   ���`  �7kl�d��jǎ����Dl�����g�jppP+W�T�eZ˭��zfO0�"���-&�#���d�l�2��!0�Xlқ��|^/�ٟi�_���� &p���½{_��v �]~�zL҈�(e��a�t��	e�Y�Q��kjj�#�<��^{M��/�����v   ��b�;  �=K$5�Q�Z[[����G�w�܎�6::�����ֶY���|&�"��ʉr�9�+����ѣ	SA6��L����k��?ڟi ���r�ڷ�v @D/,��uM�
�\NG�ё#G(���9���7�}�{�֬a�R�m�    �(�  �ö�%ຮv�ڥ���=jmm�(c�zzz��+�hxx���ϸ�Э��!2ÿ+�]�&���� �r&(��߿_���:���[H h���]���� �9�|7��܃2����_��������(@����顇�<0�]6Q���   �w   {��Pi�s?��h�    IDAT�sڵk�\����l6���̙3e[3�(6�t�ɘo��^vA���n�:uJ�|�v`R�Op7���������?h��?k߉?�s�  s���o�ZR��f�|~��'N���K���� V�_�^�=�����lG�D��&  ��0{  ��ѦM�t�wθhTc�N�>���A�^���{f:�]b�;�7ittTmmm�_V��b�=�߯{�i����-'D����F_]�+Wڎ ���U7��$��J��{:��ѣG��qF�\. z饗��/��<ۑ*E��U��X�  :��  ��m� �����׽��K����Ȉ��߯�����3�}��.w�-r��^�uuww�c;p'Q�O~�������̞1:��/�N ���
�aፍَ��uww����ہ˸���;w��GUss��8���  ,��  `�Z��n���z�'�a��Q _�<OG��ѣGK6��	�3s�q o:���;�l6k;
 ������O5��c;������$n����\��T��6������t��A�8q�	��$/^�����\;)�km   ��� (�O��K{{{c��Ǘ8�s���3,I�H$��  ��^}�պ�~���l�*�q�}�v�v�mr]�����ק���Y�F�E.X3�}f��L-����ѣZ�h��`U&���ӧ566��+4��K�#��s�4�ӟ�q�V�Q  ��D�rc1yn�S�=�	�TJ]]]�𽋻�.[�L���7�!djkkw���A��  T*�q���|��u��ncL.�N���d?����Pp��|�3���������ht��yˍ1K�i�Ԩ7vȫr'b�qFFF.Z�1�n��I  J���0��bڳg�֯_o;
(cccz�״j�*͛7�h���|Sn�GFˍ�;0=��t��jɒ%��>̖1F���:����f��V��b���w 0���R�=r�#o5Qyx>�e���['O����6��mٲE---��W�����q������|���s  �߿دQ2���8�������4d�9�8��uO����D"?�����?��tY� (*
��L&WJz��ݒ6KZ�8Nc*���$�u/�q�8�[�ρ>  �r��9�i޼yz�����b;
H�穫�K���Z�lل�3��f���߶�.�78K������5��9���N�u��Y�]�s*N�@����jկ��� �Y���|��
I�����t��1���[�Y[[�{�1}��_Չ'l�	����ێ   .c�q��!YTR��&�q�K��y�\ו1F�TJ���9c̐���^�􂤿��'_��@�(��Ѕ2�c��q��Ƙ����� @p���؎8���ڻw����mG���[���jooW4:�����{���P�uwwkhhH�/f�D>�Woo����&�z|��2'P���Xw��[[mG ̂{��H��0��y'�ɨ��K����2 �"��Gы/���������Ȉ��Ƹ> @ c�$�\��,�QI�uvv�c�$��uIE��(��@2���u�_�<�m�VH��]1Ev  *Ooo����8�n���ܹ�ɭ@�R)���Z�f�����^#���ya.��55�# ���d���k���Z�`��v� &288���n���O���%K�VW����"1F�/���?l;	 `"W�?������&���ѣ�v10w��j���jii�?��?+��>sg�Qoo��.]j;
  (��[/|�)����䘤��~���>��?��ܭ���?�4�N��1�~I�$�80  \�ΰ0�HD{������mG*R6�Ձ�j�*͛7o�ϯ�eY;�A&��g�����500�h޼y���Y�d2:w������u\W�+Vh�С2$P����_)�@@]]p˅v�͖}���n�<y�Ap@�lܸQ����������!�={��;  ��Z�:���I��d2��t�q�����?�Ї>t�r��	�q�u����H��1枑��E��   ����mG���Z=��Cjkk��h�穫�KmmmZ�dɌ�;�	�&�A�	�����y�;wN���Z�hѬw�@8������G3z^|�*
� �����M^6+w�� �\}�:�K�ĉ���.�@-Y�D?��?�/}�K�����zzzlG   �����ydd�����!c̿������Ǿf;\Pp/�g�}vw.��ϒn7�0�  HzcZ$1���ܬ�~X��Ͷ� �q��i�r9-_����ȳ-��y��K�(�L&��_]���jmmUUUX�%�����ק���k6;)�W�.A* a�O�5������lG ����#�\I��Ow���x���G���fT ���ԤG}T_��u��I�q|����v  `�1�Q����ݟL&G%}�����>򑏼`;[���^d�>���l��v�\.�`;  �s�α�������C�����r�����ؘ֬Y#�u�|l,��1���<���m@�)�J���I,��+c400���^�����ujW�*^( �7��Pp� r'8���T��{٬d�T�@����r:|�0�a jjj��#���_��^{�5�q|��;  �J����\no2�Lc���~�#���l�$܋ �HD������p.�[V�C  Nl�:�M�6iϞ=�.�����!8p@k׮��$:��������ࠚ���p�BE���
3c������۫l6;�ף����C�  ��j������ƹ�R���d2:t�PQ޷��H$��{����Y����l�񥾾>�  �58��\.��d2�'������G"��Է"�J�ttt�$��u�[�1�y  @0Pp��Ν;u뭷�����^{�5�_�^���>f����;�R�XtRss�ZZZ(���1F�TJ===E-��W��\W򼢽&��J���##���َ ���$�0�g2%9��N�u�С9��8�Ѯ]�����o~�����N�5::���  `:�%}�����;::^���SO=�o�C�1g�����d2y�q��9�s�v  0lc�V;w���ݻ)�>��fu�����N�u
�C�(����ק#G��ܹs��r�#��<�S����t�ԩ�Otc1մ��5����5��ێ ������r;m)��R)8p�r;�3[�nս���N�`�  (�1&�8�m��|/�L���'?�qۙ�(,��s�H$j:<����8�U  ��6�orG��v�v��a;
�	�r98p@�ׯW��)es)��3�ݍ-��.����T__�0i������_������%]+�z�2'O�t �1��j���ڎ ��0Op/v�}hhHG���I�/mܸQ�HD����ȿ��twwk�ʕ�c  ��Y��':::�/�u�<�J=�H$�{�|(�O�3��L|dd����o��1U  ��������8���m߾�v S���:x�֭[���7����b�~�0Op�0��fxxX��Ê��jiiQ]]����ؘ���488X�m��W��;�)�Z *��~`; `�&*�G�Ɩ�^��8�```@G��4������F���|��7�����mG   �8N�1������cGG�?����b"��@4
�H$�����~���  (�\.�t:m;�u��jϞ=ڴi��( 
p��v�Z544���jN[Ԇ��>�v� �+�N+�N+����I���SUUX�.�1F�TJ)����V�}M �k��A���	˒  ��{v��J?�Q�s9���:z�h�nR07���z�G�����f���X��  �ǉJz����d2�w��ÿB�}b�o$T�D"M&�����z$��r;  (����П�w]W��?�v `<���Ç5444���Rq�~�[]m;����u��y>|XǏ���P�ߧ���ؘ���u��!�:u�J�]zc�; ��)��+�S  f R[;��˜Æ|�����Rnhٲez���|N�Pp  �t�������������H$��v
���'?��������^�K  ��z{{mG��u]�ݻW�֭��,x��#G�̹X�xڏ˅ ��FFFt��)>|X===�N~�����߯cǎ���K�ϟ��%:w �6�ӟڎ  �w�	�a��l�x.���OǏ��T[[�~�������o;  �Lc�������dr�1�^��EHJ&����ٙr]���  �L���讻�҆lG0����ѣ��.iŘ�T�Woo�������Eٽ����u��	:tHgϞ����X�D��U��j;�
��� ����2r
�sVp��U��@����顇R$�}+&�J���|  *ZL�G���7�L&�v?u���g����ٹ_��1���  ����o��6]{�c (�q�ӟ�T�TjV���\p���@���Ʈ(����Rv/��K�O����o�/�۷ێ ��������w ����>�YQn*Ȋ+���u�Y5�<oN�_   
q�������7��cS(�u&��d2�e��^2�l��  �GX�/���[�c��1 I4U>��O~������(Z	��o���ؘzzz��եÇ�̙3��y���1F�LF�ϟ����Qj�\�Ν�# � ッ=y�v @��<�=?�	�TJG��	�0k֬�=��#�qlG�����v  ��,s]���d�ˉD"��CWp��������^Io7Ƅ�7  �&���n�I7�p�� ���6����z�嗕N�~��	�6�N4*'�Ӎ�J���400�S�N����:~��Ο?�L&����\N���:}��:��G����[###��;��k�ҋ� J#�ӟڎ  (�d�#����f��
FFFt��a��@�ڸq����ʒ;w  PN:�o���������y�-7�K��Ă���0�첝  �����e�c��|�Ͷc (�H$r���lV/������:UOr��ra����b�# (2c�FFF422"Ir]W555���U<Wmm�����l6�t:���Qe2�U����65lެ��~f;
�
���O����c  
0Y�]z���g��������Q:t�r;P�6oެ��Q������U__��   ���y����W\׽����ہʡ�o&�$uvv�NCC���  ����!eg��kP�[�N��v�� �,}�}ҙLF/�����ǧ}~���   �<�S:�����u�ĉK��Ϟ=���~��i�+hc����488���n?~\TWW�Ξ=�����*�_�z���# � ï�f; �@N,6�n>�>U�+�v.���Ç+���v�ܩm۶َQV� �MƘ��������Yʡ������7��cL��Q  _
Ӷ��-�޽{C�=%P�&�D<22����gںu�ޯ��dJ����*� ��1F�LF����UUU�����GUU�b�؄7�A>�W.�S.�S6���ؘ2���٬�1����{���g�-�� S9|X���L� ���ʭ���}�?��O!<���ÇC5��t�w(�J����v����  l3�D%��d2�����[~�����L�R���������y��$��  ���^MMMz�;��ۂ���������<�k��f�Ǆy�{���v >q�,><<|���QUU��hT�H�-Ÿ�0��O�q1���/^�j�<�>������ڎ��GG�9yR�+V؎ (�����^@i��ѣJ��eH�O\��<������ٳgm�)����   .j<�L&?��O���0�Pq���?�|������yޝ��   \����#�\MM�~�a��q�Q ��t7��={V���Z�r�_��� �2�(��4��u]��{��~q��q.�a���y�ޘ�xqں�y���h�����(s�� �"}�0w ��Z��FU�/�_��rS~�ĉ�>��F�z衇����J�R����訲٬b1fm  _�J��d2��+V�}��G+jK�����S���5Ǐ?-�N�Y   �V�'�]�����v͛7�v %TU@I��ѣ:wn��
��U�"�ն# � ��i||�Ҕ�L&�L&���Q���hddD�t����,ً�v�
-ܻ�v b��a�  r'ٝ���S��w��Yuww�1 ?����#�<������  �jw?~��3�<��v�b���{2��p6�����Y   &288h;B�8���{�j��嶣 (����s���	o��h�s�� eՇ?�Hm�� *�ȡC�#  
�NR܌��.�O�L2����_�N�*s ~5�|���o���\�
Î�   ������:;;�v�b	��Jc��L&�&�9cLaM   *��s�Nmذ�v %�n�'<�����5vU�ݛfK�J�Rp��R�ڪe�{�� *�0w ��$ܥ7J�*?A�}ttTǎ+ ��b�
�޽�v�����  `2�1插��׌1����H$����aI���  0���!�JbŊ���m� P�No�(���g?��<ϻ��0Op�� �g��߯�u�l� p�S��� P��vg���������9r�9 �hǎZ�~��%3�Υ   >sOgg������E`��d�������㬶�  `:�lV�L�v��khh�}��W��Mx�LJ�t貉��$[Z��T� ���b������ ̍19r�v
 @���I�-c�r��|�믿��]� �r{��QKK��%���o;  @!�9�����>��u�DJ&��*����lg  (DOO��E�D���*�ێ�LfSp��3g��̙3�$��3R�D(?@E���k��O�c ��ÇmG   RS3��y�@���w��ʝ �����C)V��D��  �&���˅�u��8;�L~Rҟ*�� @x���َPtw�u�-Zd;�2�m�]�:�T*�w @EZ��cZ��wَ �2'Oڎ  (@�'��R)�>}�r A��ܬ��O��؎RT����#   ̄+�O;;;?e;�L�8����o%=b;  �LU�D��[�j��Ͷc (�ht������W^Q[>_�D��Rp�����W��	����`���r�QE���,4��x��rE�q9Ѩ��jE&(�9��܉v�2F���|:�N��a٬򙌼�Qy���������-ҟ~G� �a���������);6���.�Q L{{�n��}��߷�h���d����>  �lƘ_K&�k�|��lg)T 
��7�L~�q�;lg  ��Jڮ���Uw���2 ��2�]�2���64H�#S�T�A� *��jSg�^��G5��َS��U��AU����mlT�����^�pkk��q��'*�������f�O����������S�7>�����������0��

� a��.�Ց#G4~ٍz P�]�v����:Y!�y=�S*�R��  ������R���D��x�?�N$5����:���v  �٪�	�HD{��s�@0��~��Vέ��}�"$

� P�"�}�9���S�{�E�qǭ�Vռy�-X��y�T5o��,P�¯c--�͟��y�mn�㺶#��[S#����t�3�R�}|p�ү�}}���eϟW��W�CC��� �R��J�	��[�fg �亮��>��_��2���8E���K�  �1f[}}��D"�1�H��͙��D�����5IKmg  ���
)�q�jii��%ź��<��̑#rΜ)���C� B������N��?��/|�v_pkjT�d�b���Y�HՋ�QboiQ�BY=�`A`&���\�a�^6�lo�r�����)�ݭl_��Ν�عs�vw+s挼���|:�\���  vLUpw�F�=_�4e�t�̎�S ���z�}����W�b;JQ�������v  ��ZU__,�H\�H$l���o��=�\c6�= i��,   sU	�U�Vi˖-�c ��u]9�S��F�=��"�>+�r�y� �Lq PYܪ*�y�)5nۦC��{ʧӶ#��[U�Xk��/׫-z����g=yV���j��T��6����9wNcgϾY|?}Z�S��9uJ�
�ɬ�FO��� >�����*��^]-s�}RHv�PZ�֭ӦM���~�Q�l`��=0 ϟ4�    IDAT �B-jhh8�o߾k>�����3_�;::Z��쫒���  P###�#�I<׽��[�r+��)���K/�y�9_�Rq_�ǜ�*�  e���{հe��tt���߶gvG��f�R�,[v��,Q��E�8!��MM�ojR���~=�Nk��IeN��Tz��1v挼��X�̩Sj��r �&�Ko\|���p��el� PA��N�>}:��Jl  `�Yh�9��ѱ񩧞궝�j�+�'�z�uf���  *B:�V6��c���=�ܣx<n;
 ����>z�w�=xPΫ����h��� ��T�d�6�ۧ�o[G�{N�c�lGz'U�ҥ�]���{�e�Y�Ln,f;"(��~����̹so��/�އT�/�?����:e; `��y<�]�7�Lr# �V,���߯/|��<�v�Y�  �X�;��j"�X�H$|u��
���g�T�1f��,   ���mٷmۦիWێ���Op�$Ǒ��w+�o�4<\���ʁ n�o�]�v�V�/���oJ��J�3D�(�/]���v���U�t��k��s
�庪Y�D5K�H;wJ��lV߽�.y���p�d(���9Ӽg�����hj�w��S �P�-ҍ7ި�}�{���Z*��  ������~������7[�����矏����:���v  �b
����F�z뭶c ����%��Q�;�)����4��# ������r��J�߯��G���?){�|Q׉-X�x{��֮U��]�ի_�JѦ������������ڎb��ɓ�#  ������e�QR�#s���1 �Ѝ7ި��.uwwێ2+� @j�f�'��b
�/
��7�L��8�
�Y   �-���ў={TUUe;
 (Y�]���:��X��I��4ݔ7 @�4lڤ�M������4��K�я4r���Ξ�)`��؂�]��2{�ڵ�66��O _�M7Qp �Z
�f�f�\�PZ��������y��w  P������c�:�c�M�/
�������8�m�   (��!���3#�6m�
.d ��uݒ���w�NΑ#R�7��D���v ����7nT�ƍZ��c�$/�U��Ie{{�e2�g22��HM�"���SͲe���ZW�֭�#X���<O*�{o ��Mw�z࿃���m��N $-Z��۷륗^�e����5::�Z�� @�qgugg狒v��b���L&�_c̍�s   �����3��u��ێ�GJ9�]�Lc������/�t��� (��)�ޮx{��(@Yխ_�F�;������Sl��I  �p��y=���]w�p�>�2��[t�ȑ@^K��  *�M��SO��f�7�wvv���o3  @�q�����6Us!�eJ=�]�̭�ʬ��ͽ"�  ����(�j��Ve{{mG  La���+�)O��ko�Y��v
 !�F�g�9N�{���ێ   P2��<�L&�63X+�wvv��1����>  @��R)�fd���Z�n�� |�w9�̣�JQ뛍��SUe;  ��}�
� �o���icu��l�b���v
 !�|�rmܸ�v��  ��~����m-n����g��n�����  �-H�X,����v >�n�&蘅e*��tS�    �,]j;�U���
9�b���v�T_o;�������mǘ���A�   J��?��?����e?�N$����/H��{m  �r3�(�NێQ�]�v�� �R�����KZ���k���َ   �{��mG  L���{�.����\{�� B���F�v�cF(� ��pc�ط�D�/����^__��ǩ+��   6�R)y�g;FA����m�6�1 �P$R�K�Ѩ�(�e�Pp  �Vu[��V�lG  L�'��;�ʴs Le˖-jmm��`��ö#   ��1&^WW���1e=�-�b���_����k  ���w�qG�K� ����u�̚5e_��"\  �XK��V�َ  �B�Mp_�^&仧 ��qt��ێQ0
�   L�Y�o߾�+�e+��۷�Ƙw�k=   ?
ȅ�+V����v >�vf�y�|�di�R`�;  ����Ϸ�*&�������i�U����۽�v
 �²e˴v�Z�1
222b;  @YcޑL&�c��+KS�駟^���?[��   �$�Jَ0-�u5@�Y�ݡ�M�7�Y�\
�   Ӫjn��8Xɘ� �7��A�)f��^jl� ����oĎ�� @H�Igg��r,T��kc�[[[���8�R�  �7A��u�V-X��v >fk��$���jj��_4�+' e   ls"E�q�1��� ��VWO��@������i; L���Q;v�cZ�lV�\�v  �r�Hz!�H��^�¾}��$iq��  ���a��TSS�]�vَ��N˩���g�������   �s+��Y�ڎ  ��t� Lp7��*UUَ ���TWWg;ƴ�0�
  �،1������z߾}�4�<X�5   �,�Jَ0��;w�&�� ��9�]��m�I��[�0Wn�M�   
5]q�����< @�}�{K��5��N S��b���mǘw  VƘ;;;�]�5J�Rx��=���R�>  @���؎0�x<��[�ڎ  l���{���f�+�S�  &�wy��l�v
 ��inb��ws�-��؎ �ڲe�mǘw  fƘ��H$�K��%;���$Ɓ �P�s���nP,�@ X/�K27�(��؎1kLp  (\$�;�y���#  ��VUM�u�/��ʴ��N q]��S����3  @�U744|�T/^��B2����8ח�  �į���:mٲ�v ��a�W$"o��)fm��n   xS�'�K�Sp _+������y7���v ��i�&555َ1)&� ��3��L&�.�k�����k��Q��  c�����馛�l	� �����.�\���j;ƬPp  (w
� �kA-�/Z$�Ze; ̈뺺馛lǘ�  $I�D"�\�-��u6����p�}  ���=ϳ�-�y�f�1 ���蒬�ʻ��)f��;  @�(�Sp ?s���Lr̔��V���k��F��ϷcB~��  ��buuu_.������g�y��[���   A�ש�v�R$�@@���.�l�.�d��3��}  �`N��J�Qp _+���y[�̊�S �����]�vَ1���a�   |�q�[���/�k���H$����Q��  :?��q�F�1 ��
�r��ﶝbƘ�  P8'��e�\�v �
9�����C�P�֭Ӽy�l�x�QnN  ���D"Q��E;�nhh�s�q��z   A��m	���:��U���Ef�V���1f��;  ���=h9��q�  S(d�����.X �|�� 0'��hǎ�c�w  �79�SWWW�ߋ�zE9�~��Wc�[��  �~ۖ0�i��Ͷc _��2�w�N1#�  f �wy�� �)m��ٹ��� *¦M���mǸB:��1�v   �p]��~z]Q^�/����X�  P)�6�}�֭��b�c _�%��n���Ō���  
��]�ʉ	� �o�*���ˬ_o; E$�֭[mǸ��y�f��c   ��1Ʃ��y��5�c뎎���1ۊ  ����i�.q]W۶������XLf�.�)
�w  �y�ݣ� ��VUM���$3�]'��� �����UU���r�ێ�   �9���������u�|4�8���k   T"?Mp��k���`;� ���Ls�mR@��Lp  ��-��ێ  �JP&��b2�^k; UMM�6n�h;�R���   ��D>=�טӱugg�KZ0�   ��Oܯ��:� �o'�KRC��Ȃ ��    8B^p���N  �B!�}q6��k��j�) �访�z_��f�;  ��tvv>9���;>c�����   �ltt�vIҊ+�p�B�1 ��.L��qG 
PLp  @��� ��	�wו�}�� PMMMZ�z����iGg   ?1�$�1�>D��;;;;$����   ��/ܷm�f;� s|^�1�ˬZe;ƴ
��  �7�\�v�x� �V��i�gSV��m� ��ٲe���0�  `Ru���4�'Ϫ�����ǌ1�>�E  � ��؎�x<�) ���wI27�d;´()  ��fmG����.J vnUմ��}6�\{�� PZ+W�T�On����+   �����?��gu��ĉ��f�   @c|Qp߼y�\.��� |1۶���ڎ1%
�   �{�]��� �)�~�{]] v���pG�7o�C�422b;  ��Ŏ;���g�T0Ƹ����l  �t:-��f���= ��	�v찝bJ�  
gr9��r(������n6o�0�  ��/C���  05�u%�H�������%��?p�f��  ?��Z�l����m� p�(�K2�vَ0%JJ   ��w��#��ܪ�ic�l��H=���Z�r�����  ����럞�f\pw��f�  ���C�}˖-�# � �)�/Y"�|���b�;  @ἰOp�# �Z�w+gT�/�ij��2 Xq��ڎ@�  �01�̨�>������E  !�����Y��j (7s�M�#L�)�   �3!/��5l� ~V�H6
' Bf��ժ��[c��  P�ڎ��'g򄙵�]�7g�   �FGG���q�FE"� T��Lp�$s�uR,f;Ƅ��	  P8/���*
� �s~-����0�@ȸ���7Z�066fu}  ��p]�c3z|���'>q���'  !��6X]@ep'PwUW�X��1)n:  (X�'�GjkmG  L���*�qe?��n���h� T����[]��5A  � Y����@�.�7�t�.  @��<���РE�Y[@�T���m��r��  P���a���� �V�.m�>�b֭+� �����?���=�S.�7�  ��>���{2�\)��Y'  ��6��
�����l�$��؎�VLp  (��<�C^pw��~ pI���:K=�Y���+���]�����t���   ��B'}Z�Ww��.j   Ae��n{+F �#�wE�27�N�Lp  (L>���<�1�b�; ��/'��]+�e����lذ����  
�H�d!,�(���g  �L&ceݦ�&-\���� *O ����#�E��  �.74d;�UnM�v� _+t�{9Ϫx=r---�?���m�  �w�i��d�$1.  `l�7l��B* �	���a�TSc;�(�  f|p�v����mG  L�w��q���\��o���	�   3R��3ϼo�2���E  *cccV�]�n��uT�����\{��W��  P�w�  �(t�{٬_/��n� �kÆ�֦�  03�|���{̔G����/ic�  ���	����Z�pa�� ?2[�ڎp
�   �a�;w �;�Mp7kזi% �y��i���V���.  @�m��Q�Ԕ�|>�;*��i   �"�͖}�U�V�}M �-��u�⮏J宏�   ���А�VE��lG  L�O����L[�� �����|  p��y�y�LYpw�狛   (��e��L{���8���   ����n; `nUUA�+�؀+$w�K� *���ٸ.  P��Oz���Oz��%E�  �\���E"-[���k�ߙlG�����  �n���v�b�Ͷ#  �Qh��,z WX�l�b�X��+��   �-�L��싓�GFF�Ki�   T6cL��˗/W��$�"s���+s�5�#\⫋�   >6��m;�UQ
� �{~��ݬ��  �亮��P�  f�q�ߙ�k���y�4q   *[&��1��k��r |m�"i�<�)���N   ٞ����� �Wh���cZZdJ�
 ��kf�  f��}a��>��EƘ���  P�l�Ģ� ��w�G��   �l���� �i�e�6�9a ���kf���  �Rc>��3K&�ڄ����'K	  �r����u���F5s &d6l�A���/  �-�S��y�)��� ��c|
� 0���F�+�ΞLp  ��|>�щ>?a���Hi�   T�l6[�����T��i��Y�Nr'<�-+�\�  ��^��lǰ*��d; `N��KzV%�Y���+ @��\����1�  `N&쬿�*"��cV�>  @e�d2e]oٲee] ��Z��_��  �.��k;�uU���\?�ľx1� `
mmme]�	�   s�����Ǯ��[�z�p��a  �Y*w�}ɒ%e] ���`�7�  ���==�#X�����؎ ����e.n@�,-�Гr��  Pa�'N<��O^�	c�{ʓ  �2�sJC}}�ʶ�pq��n�]6~(��    ���E�lG  ���{)Ϫ
� 0���:566�m�\.W��   *��y?��&:��Y�,   ���ro� \*����n;�?Lw  𹱳gmG����  0
9�/�YǑY��T� ����r���a�	  �l9����GމD�YҼ�%  �@�܆��; ��Af�|�(�  L/s��VUSV���z�?�TSco} �r^C�<O���e[  ��߷o���8�nhh����  �<���V���~�L�  (���-� P '��1%��ti�^ *J������   @%�<�������1���  �<��PUU��e- �TI[��U����  0��ٳ�#X�� �aq��Y���� $---��be[/�˕m-  �
���s����2  �H�:��x�b�6��P�*��.�w�[�  ���)��k;�UՋێ  (��	��� ��hI�gRp  ��+:엮�c\I��  ��VkkkY��J`-��Q�1   0��s2�g;�U5� 0�����4����y�g~�_���g8�C%Q�J�(y�^�k;~�N$@�dÈ8FbA ���ȉ8�"F� ��I��țc�s���]kq��cuߢ$��x��9���]��!Q��ǐ쪧����%9�~�$�ͮ���{6�Y������������� �FY�m���?��M��������?�L �JUܯ��J�h�N'��Ү ��J!�,���#Y�}۶��-}��ڶm[ek�� pu�������ƹ���=�f�H  �2*Y�ʩ�x*���N�Hx�w��  1���֭��vS� `��q�_ʮJ�EM�6���n�; ��˲��.��~���� h�*
�N'�n�Z�: mR\�c� ����c�����o_�8��G���pe%u4(]������<m�˖ML$Y�Pp�,[�n�N�y�����; �H��|��~Kۦ� �P��[�l��D7Q kǎtk;>���WW�䣏Ɖݻ�����#�#��\}� \�Tw�.Ϲ�Qǎ+}�*� ��[��`2"�(������̧� �ULp��HE`|��!��������r �ǙW^��_�b�s��18s&u����e��#�Uɲ(��fԯ
�z۶m���n�; ��˲l�(�N�e�dD�����~6�I�  �Pńw�+0?�qcD�"af�; �������~�|��Q������ �Id������~]���Ꞛ	�  W�(��?�����F��'#"��_O�	 �5Lp���"{����Upk��c���N���Q������� �I
������; @��ÿ�
��a  ڤ���[���@Q��0���o�HPpOr���<���ś��{���������7�� ��X�u��wU6o�+��-[�T���; �hLLL�?�
�H� �U�</��;�N��ϗ�@[[�D�Y�	� c���;��o�F�z��Q���t�1}���c p���K~���6������|t:����U��#m    IDATq�3 �8(�ⶈ�
�EQ�9 ��pX�����E�$`�+��w��r���_���;�:
� 37�����I�],,T�&@t:��������R�)��  ��>"�ܕ��  #R��M&� )��,	w Jv��ߎg~�W�ہu�p�-�# p�RLpWp�r���r?  ��("":����7�{�� �zeOh�b���Dw9�ño~3^��"����Q�Qph�u<�>�{̛Yp��e�; �hdY6���~cgÆ?�: @��=�A��JQ��Vlz��33կk�;@�߽;^���2�� u�afo�5u .W���وnw��0V����� 0:6l��N�e?�: @����E+�Ql�R��&����={�_�u�v��̘��J#�U�'pU���V� , �q211qO'˲;S h���
�@U�Zp��[�_�w��Z;u*��G�(��˩� �A��q�� ��;@}lڴ��5Lp �;;��K ��
�@k(���������GS� jbn.��\�: �i=;&#�U������
�G� F�(�[;�N��A  ڢ�ͫ����� �x���ƒ{�qc���c� �s����8����c 6��O�� ���qR�HwT�	\�*�)� �N�e;:EQ] 0"����ן������R� ��6�S�^��� 4�`q1�����:�pswޙ: %�J133�W?U�_Sp ����H0� ���޼ڰaC���Q�,��ͥN @���S��:�:�p�wܑ: W`=��tGž0�U�)�a!w ����D�ǽ F��ͫ�7� >J�}4Lph�ށq�K_Jh�ک���\���H)� �ԆNDL�N �&�m�Ƃ{1;[��
� �����Q�q��	� �e���wS�\����y^�� ���NDtS�  h����&�Ukc�=�w �c���x�k_Kh��֭�ݺ5u �D��¾0�Us� �Q�:Y�# 0"eAMp��ڂ�%nD�Zf�;@k���"_[Kh��;�L���t7%�"��p��.��r/  �,�&:EQT{W ��Lpڦ���݊3��P@y�K�# -1w��# p�.� �HwS��#<8p��"�ʽt �D���:Y�.; ����y5mRP�<�SG(G�'b��h�Ճc���S� ZbV���F��R�C� -U�=6w ���Lp ������>�G���^T�~��r�v8��C�# -2w睩# p�.q�?Ҋ�=a���|��; �He�2 ��7�܁��vS~r�����w��8��#�# -�ML��Ν�c p�.q�?�q��F��{l��K HD� `��޼*{��G�u�{Vu���+�Xz��)�����'�3=�: %Qp�w �fѐ ��7�&�,dD{7�
og
� ����[�v�d�@Kl���� �
���Wp�w �fQp !܁���#����2�� ����3�# -2�kW� \w��)���; �h�� � eO� ���n�Wy"�	� ���쳩# -b�;@�]j��HwS<80&� 4K�, ��)����;P�<�̱����T��܁�ɲ�۹3u
 Jd�;@�L�<�D�
 `�:�z� ��+{���>��w�����Xٷ/u�%6�|sLnܘ: W���~��;@��� �,R   \Pk� p���%&���x�=�# p�*-�+L�D�tF F�(
w �Q*{�J��Zk��խ���μ�b�@���# p����_�N�}��^� ��Ȳ,:�-+  $Pv���P��(�Yr����� c��K/�� ��§>�: W���#��W��>@��}��w ��2� `�܁6j���n� cfI��lr2�v�J��t�	�#�	h�@
�  ��� �9ZY2j���*�޻m�ĉ�=�:�sw�����1 �Z���c�wCO FB� �Y:Y����  �FٛW��	����?S #K/��:�"��d� ���f�c�-ܗH��!R
�  #UtZ9�  �N�S������������B����^z)u�E��A��y�"�� 0Z�  ���S���k�{O�'b(�4֙�_Nh��O:u F�"��q_ ������  F�w �*{�{+K�@�q�{V����&�Pog_y%u�%fv��ޚ: #`�;@�(� 4K�, �1S�����j��p>�|�fe�����i���G����Ė�~6u F�b��#�E�'0e�cSp -w �*{�j��B&@D'���vz@#�}�5����l��=u F��	���)� #P�=6w ��Rp ��7�z�^��p>m���-/W��r$@#�}�����ޱ#>���1 ��"{%e�d����!R  ͢� 0B�N��܁Z7����ʗ���� ���믧� �Ď_����"���P(e\5� �E� `�&&&J}}�%��6��HPp7�����ٓ:���6����c 0By��þ0�U+{�T�� ƍ�; �)�mTE-*hg)&���!��P��wo�@��w�nL�Φ��eOpϜ�	p�� �E� `�܁�j�����	 h�ޡC18s&u�᦯�>n�;'u F�B܋0�����Pp hw ����,����a��������y���H2��E �b���SG Z���O�33�: �v�	�]���pU��~�{ܝ�
 �(�t 0Be�#Lq�h�ww �ᬂ;p���sq�_�K�c P���$e�dN��*����� 0Z
�  #�eYdYV������>���i�{�8Q����@}��ۗ:�`37�w���: e��>Ii�'���J��� FK� `��>�P�H�U�S��� ��Xy����������ߊ����Q (ɅNj+m�Ğ0�U9}�t�k�} `��t 0beOhPpRhS�=;y��EMph��7�Lh�lb"��w�.�v�L�2)�4�	�  ͣ� 0b&�mԖ�{����U�n���(k�NŠ��n@�t:q�o�Fl��gS'�d�Op��#K���
�  ͣ� 0beo`Uq�"�G��F�8~<ͺ-y@ `\��z+u�a��ɸ�������ϥ�@.Tp/u����+�� �<
�  #�eY��o�;�Bk&��<�f�$�p���ۗ:� ����ݸ�����Q �J��#">�b
�  �3�:  @�LN����ٳ��yt:�U�SE+�{�'������qa�;�^���?�[�n�5u *t�	�^�|pE���byy��u� F��� �*{+�sS܁$Z1�=Q�=�"ͺ \�w�R�,n��_�������0��Sp����,�	� W��{j
�  �e�; ���=�="�ĉ�y�������pSSS�c\����4+�4��}�# 5���[���Oc�O�T�( �P��^�X�T�4����+Y��{�  u�� 0bU܏;��~{�� |�`0H��>�d�]@�y���O����뮋���ߏ~�"3�`|]�!���ǎ��@+������V� ��Pp ��
� UK�U[�lq1�̙4������G�硫���wĎ���㺟����0��쏔>��{w_c�ƲWh��� 0Z
�  #V���;�B�������6��1z��� ������/�����??�c�� P'�&�GDv�X
� �E� ��� F���S�N�p8�	G�jz��s�p����c5�@��d��pCl�瞘�ԧb�g>�;"�RG���T�㽂�m�U�@;���XZZ�d-w ��Rp ����?b�yǏ��۷���9�A�jK�r"���P?
�7���+u(M656��ƍ1�eK�\w]D��: M�p�{8��;v,���f��n%�  �w ��jBñc�܁J��B�)��=�����Ŭɠ  �u�	�
� �s���Mw ��2� `Ī��Q�@DDQ1��M����G�-_4�� �q2�ܳN'fv�H ���s�_DE�'λ> �W彴�� �w ��j��;�S�: 4RG�"ّ#)�����^p����: pA�{�}��K��|�nU�K3� `�� F�����Ç#7��XS���I�7��9V�I!���nJ ���w�_�nIv�`��4�`0�#^�+� ���; ��UUp_[[3��\S�Y�{f�;@#N����r�Im����  j�?�k��(��ˑ#G*U��A �q�� 0bUn`t3�Xc���%]�w�f���&� \�yb�t����*Wh��_�� 0Z
�  #6==]�Z��l-����O��8y2iw�f��|�� p	�y�F*�-9{6bq����{h�N�w �Sp �*�UO� hb�={����o���; �%�kk���wK2f\TQ�ܕ� FO� `Ī,��={6M�*TE���1.K�o_��;W�ÇSGHn�RG  ���<����3�O .�ĉ���*[���V� ��Pp ����J׫r@D���`�����P?��GSGHjbÆ���O ��>z�?����m�'pQ�t=w ��Sp �*'�GD0��X�&��z�8��h�C c��D�IM_w]�  ���k�$W�ǏG���be�FPp h>w ��z���}�*]�Iܳ�^��+���1&�4�ژܻ
�  �4��?��$�$y��)V���(�͊�#� FO� `Ī.�/..�ɓ'+]ok*kg/��:BDD�;g�^p�Qp ���^��)���ѣGcyy��5� FO� `Ī.�G��T�Q�_y%u�����w0��<��N�N��	�  ���Sڒ]���Q�V���̦��+_ ��� F���F�S��,w�J��0u��9|8�.'\(���کSy�:FR�۷��  P��Ovf�ٳǎ�Z���Lp	�  ��� P����J�ۿ�&*͖�y#J�u�����n ��Z]�Jh�w �K��)m)wH2�O >duu5>\��
�  ��� P��7���a�߿��5��ր�v��˩#���@�>�:Br�k�M ����""�@Y�)� u��oF��t������ h;w ���԰ϴ�B�?5�ߏ�7R�x�	� �7XZJ!��͛SG  ���#�����S� ��T��Lp =w �����F���@��}�{��5*��P&�GLnڔ: @��(�'����>����(��7lؐd] �6Sp (A����ӧ��ѣ�����OpϞ}6u�Qp���Op������s  ���k�:�N�^{-u�Z8p�@,//'Y[� `�� J�j#��W_M�.0~j=�}0��R�����_ DD���b�IM�� �.���k�8�޽�:T��ڳgO��� FO� �333I�}�W�(�$k�%����c�W����^�b�;@����Iw �u��Vp"۷/u
���<���h1;;�lm ��Rp (A�I���q���$k�gP��v��ө#|La�;@�ΞM!�Ʌ��  ��C새��Fy_�pj1@�߿?�����?77�lm ��Rp (A�	�i�`��ZK���Zd/��:�ǘ�P��J�IMmޜ: @#���^�+�7ވ��S� H&���T��  �L� ���EQ$[��������S|��;@��SG  h�s������0��{S� H"��x�גf���M�> @)� � �F���R>|8�������g�I���]�ay��:BR��#  4¹���v��9�So��V�^�OMM���d�� �J� ���"|�W������{���^J��Lp����r�IM$<�
 �I�:Np��x������M`<�I�����t�� �J� ���"|��c8&� �_��z�ɞz*�����c�;@�WVRGH���  ��{���{�}8��� e�����3 (��; @	ROp��z��k�%� ��:Mq�}4u�Rp���O�̦�RG  h�|m-��r�sϥ� P��_~9�O�4� �
�  %H=�="���Ou)�g�E��T$����5�7-� ֧X[��~r<q"�C�R� �L� Pw ���ͥ����S�N���\m
�?�:�E�{i�	��0u��� �'_[�~�a�;0.�9G�MC� �$
�  %�������������
������][�x��).*7���ƽ��MM��  �����gO��j� �{�RG��z�� �F
�  %ٰaC���/F��c -6�(���g��le%i�KRp��q/�w� ֥��c0��WR� (���Z���˩cDD=Nu h#w ��ԡྼ�{��Mh����s˲GM��z
� �7��n7u �F��Q�O��sϥ� P�={���t�0� �,
�  %�ˆֳ�>�:�rIo$:�o�[��� pi���3� �e�	���١C�S ��g�I�}7nL ��� JR���[o�G�Mh���;>�l�ˡ�� y�:ARY�V1 �z��db�dO>�:@)�~��Z�����K ��ܵ  (I]
�O=�T�@�%��~�tdy+�� ��,K� )c �OS
�����N�N0rO�������  ZI� �$u*����+����:�R�� ���|��CE���{%
�A���&&RGHʿU  ��kJ�=�3 `�N�8���K�CLp (��; @I괡��y<��өc -UE��P���#�T��U�Mp�=ww �K��<����^x!�^/u��y�'�[�� ʡ� P�:�#"�{��7e��8k��G�XY�tͫ�4P�^p��[ pI�^/�A�"�}6u
��X^^��_~9u�����n��: @+)� ��n�~��?�|�@KU� M�G硇�[o�&��S��d�I)� \Z��k�5~����a� W�駟�a���6lؐ: @k)� �d�ƍ�#|�SO=y����P�ܳg��8y���F�i7����Opw� �%�z�țv�����M<�\�~?���
�  �Qp (I�KKK��/���P�ߏ�(�_�(��o��ΈyEͦ�a�>��0� ���8�=""}4�����~����z�c|��; @y� J�iӦ����G���@�E�
n�fO>q�P�딡�7�����L�I�� pqy��j�E�⋋���B� W���ǓO>�:�y�q� @[(� �dzz:���R������x���S� Zhuu���<�(w�)���ĘO].-��  Pk������G"�_O<�D-��G(� �I� �Dsss�#��c�=Vɤe`��K���=�xd�S�e2��:c^p_;u*u �Z[YY���{�g�Ff�	�0�^/�z��1.H� �<
�  %���M�Ξ=�>�l�@˔Zp���o������RG �"�}���; �ŭ��4�����"krI;�?�x�U����B�  ��� P��Np����~P�MA�y�A�y^�kg�>q�x)�]�B����� .fee%���./G|4���J�5�� Pw ��yckee%�y��1��)���� ��Oo���WWSG �":
�#  �V�������#"{���9��k �M�6��  �Z
�  %���O���XYYIh�2n8d��nd�O��u���z�# p�5~8�
��[ P��{��m(����%w�;}�t#�4-,,��  �Z
�  %��������x��S� Zd��3g�ӂ��C�jmŗ���>Q�c  �ҹ!!m9�-{≈���1 .h���1SǸ�,�j?�
 ��� JԄ��?�|;v,u�%F]p�|�k-�|n�;@�M6�{��� KK�c  �ҹ�{���8Ɉ��y��) ���ߎ�_=u�K�v�155�: @k)�*��    IDAT ��	�<���Lh�<�c0�����?�k�@+�1h��1���z�p�  �SE��{h�U��{�D�ߟ:��4����\�  ��� P��Mؔi@3�j�{��{#�b$�Um9����}�{DD�С�  j���E���D�
��y���<O�}M:ux�ƍ�#  ���; @�65h
��ݻc8����(
���OG�w�����io ��d�>��eU� �cVVV��qѲ�{��Nt^z)u
���X]]��~8u�u3� �\
�  %��������1�������SO������N*_[��W�:�05b�;@�M)�G����  j�����6�=""����6����y�G>�PQݙ� P.w ��5i��������1���_����7�q��Ճ�;@�u�mK!��ÇSG  �������ʂ��rd��~���;v�X<��3�c\�&�� �D
�  %kR����Ƿ����1��+�"�Wx�7;|8:�����C��Pk��11;�:FR�C�RG  ��~�kkk��|�Ƃ{Dd�<��|�D���o~�W54%w �r)� �laa!u����oĞ={R� n�J��E��q�p8�@5`�;@�u��6u��z��  P+��(��JQD���ݓ����C|�z��ͩ#  ���; @ɚVp������+++�c v%ܳ��l߾ч����;@�M�y�}��k'N�� P-�����ĉ�<�x���Y\\�Gy$u�+�� P���  ڮ�������w�?�3?�:
�P�~?���,����٩Sѹ���S���z�# p	�m�RGH��޽�y���1��G���[o����,/G1���LL�����B��v[Lnڔ:& 5��! E['���裑���σ@E���\Ѱ�:Pp (��; @ɚ����/��w���rK�(@E�~?������ٟ�iD���ED��?@t�oO!��{c�O�D�pU�Ǐ��k����^���_�3���o�����n���;c��xl�ɟ��O~2��0\�q������e����yd�gQ��/F�sh��z饗b�޽�c\�n�6lH ��� J�����x����_���v��� ������{�䓑��b��Rp���;RGHne߾�`݆�˱�o_�ٳ'�_=ξWj_;y�_s�ĉ8��q��G#"bra!�������\,�؏�*: ����cPp��8t(�瞋¿{@����c��ݩc\�����  ZO� �d[�lI�-..��������/��4��:
���bt�4�)����M7����rC���bE�Ç���[��o_����o����E���җ,.ơ?��8�����7�ʯĵ��\t��J_��Ξ=��_�k��ߍ��#����w���>H��#  ���; @�6o�Y�EQ��\�g�}6n��ָ���SG���GQ�]�H뢈��0�<7��h8&7��l��SGHny���8��]٤�c��?~<z��Go��Xٿ?V�|����z+�5)�,��{~�7������������o�-�?h��Np_[K�$�����w_��K�N�4@�<���gϞ�1����|�  �g� �dSSS1==�^/u�+RE<���˿��1;;�:� EQD�ߏ����~=۽;��_�8U:�2���fn�!���(���Q��8?�����tb���c��bÍ7��1�cG��xc����m�".��G1D�С����
�y���W��������Q��k�[��SG`���yO�+��i9z4�G�ⳟM�h�S�N��ݻSǸj&� �O� ����-�GD,//�7�������Ob8�����ܳÇ�s�}	���P��dt��.VL%�<�����;x0N?��Ǿ��v?^~߱#�w��뮋�5�$MJ���X=z4V��#G~�����;t(�G���ᑕ7ߌ��?��~��b��zd�#0"������������?���(n�)u��<���?�-xXH� �|
�  XXX�w�y'u���o߾x��g�ӟ�t�(@���f�`����#��%���n�I�}�~?V�|3V�|�_�t�ѽ�ژ޾=�����_w�|�1�u�BpC���/������ñz�p�}��~�PWVR�L�ȗ���Ÿ�����t��� 0+�w��k������#~�W���	} ������ÇS��͛7��  �z
�  شiS�#�{����c۶m�� ���EQ|��Η�q�P�Ti|��8��馈�K���~?zD���~O���Ԗ-1�ukt�o��֭�߻۶Ew۶�ܼ9�6o��M�"�&52E���ԩX;y2�ǏG���X;y������ɓ�v�D����'#o��Ų��x�������-n ��ٳg����6�=""Μ����ٟM�h����9���lْ: @�)� T�-���a|��_�_��_�	7�u(�"��~L�7�k��T�����Jc즼4Ԇ�nJaly�~��쫯^�{�N'&7m��͛���M�br���n���7���BLm�7���������;SS������pi)�c����/.��̙w|���S������[������o�f�������z�k��=���Wc�ƍq�̙�I���zq�}�Eޢk��  ʧ� P�6Mrx�w������Z�(@C������t����'6o��"u�$��&8@�(��S���O�\�n�C��ɍcbf&�n7&fg�397F61�7F65�������N����+,O��E��|���~?��Lw��D1���׋�ߏ�ߏa��p��rE���w��һ���./��̙��\Q�^�|�+1s�q˯�j�( \�Mo��	��yǎXݿ?���SG�(�����c�k�6��������1  ZO� �[�nMa�^z�رcG���h�(@�z�ؼys|򓟌�+(����;@3L�xc��X��G~�D��8�:
c�������㎸����Q �g.0��(��.�O���w�/��R>����<��ño߾�1Fjaa!2'6 ��s�o �j�����o;<�:� kkkq�w���|L�̤��L��a�*@�m�馏M��,E{����U�� �t�	�kkcz*]��D69�n7n����q��ػwo��?Hc�Lo ���; @�l��N�>z�y��w�#i�K���k����LO'N���w�ڛ�����Oh���3���Wph�~�k�Ҟ�������������ǎ;'��ԩSq���G���6mڔ: �XhW�
 ��&''cvv6u��[ZZ���/r7������n�)Ξ=�1���+�4��Ν�# -���3�����c pΜ9s���(�������ϯ��zO�������_�r�[�`Ж-[RG  
�  i둅o��v|�{�K����ɸ�;"˲ܻ��'~����7u �fV���������J�u:�q>���z�#�,���n��1?�8�o}�[q����1J�y���  Ƃ�; @Eڼ���O�K/��:P#�N'��Θ����w�����Y�1��9��RG `6*�#���������c �EQ��������C���˙���;�3&''$���k����[���  0� *��#[���?��?��L��s뭷���܇~��M≙��jA���܁:��#q��S� �VVV"��~}���0�������;��Q; "���?�p��Sp ��+M ���y�{DD���|���N�s�7�w���1��<���� M2s��1�aC�@���/�%���&H�ܾŅ�u��"{97n��n���0@-<x0����GQ���*˲��kR�  
�  ���~?��ދ��۶m����?��Ξ=EQ�u�=_]M�u�:������1�Y޻7޹���1 ��K��������ٲeK�ر��4@ݜ>}:���p8L�t�����vS�  
�  ٶm[��X\\�{�7���RG*�����r��>����D�a��: �4�sg�@˼����)� 5��y�.q͞��~��:��p�c1���������86��6mڔ: ��Pp �����SG�̑#G���܍{6l��o�=�,����={62�h w`�V�z+N<�P� �Ǚ3g�(��~O1����:��v�m���Pr�.��a|��_�S�N��R�-[���  06� *2==����cTf�޽�{���1�
t��عsgLLL\�{Ϟ=33��'w��ظkW�@�?�'u ���ٳ����8Op_g�=˲��'>1V��0��<��~��q����Q*�
 ��(� Th܎.|�駕ܡ�&''c�Ν155���_^^�0���x�=�MN���̩���7�L��8s��%����9�W�aÆ)E_���c�޽��TN� �:
�  Ǎ�'�|2{��1�LNN�]w�3�9�}u�˂
� �љ���wݕ:�BG�/u >`ee%��%�/��+HSO��(�G���޽���_Q��o;^y��Q�ضm[�  cC� �B�Xp������O<�D��MLL\�4�^g|/E�++�# p��GSG Z��W�Q�c ��Lo��k��
N㛚��]�v)�C�<��C��Ϧ����; @uƷU  ����#���|��R� F����w����W��W;��:�py9u .��;P�ޡC���۩c �����T������n�;w+��@���0�N�3���  ��� P�q��PE|�[��c+�-Ε�����E��b\���x�@m��Kh����SG  "�A�z�u}o���k��Lp?gff&v�����#LT����{,u��bbb"u ���� P�q.�G�[r��׿{��I����W�:Y��Z����(�;vD��kR� Z�w�@� ����GDǹ�~��7lؠ���O��ݻS�Hn��ͩ#  �w �
mݺ5:�����y�����/��\�N�w�y�U��#":c\p��g�S�Jh��	� �p9�|u��$�v5�ϙ���]�vE��A"�*�?�x|��ߍ�(RGIn˖-�#  ���nW Tlbbb$�Ц��<x��xꩧRG�abb"v�����#y���L"b0�Wk��g�ӟNh!w�􊢈�gϮ���q��>��{D��̌�;4DQ�{��x衇RG���[���  0V�DD��aP����]�N�ژ:GjEQă>�~?~�~*u����b�Ν�aÆ����{7EW"b4����W�uv=@sm��Oh�ށ�# �������|��?�����^���Ʈ]���W_����B������O��R+7n��S� �	Ûa�)������H`���+�C���?kkk���_H������뮻bf�71#"��
����P��q��'&��c���:
�"+��GED���0��.��	��������VΝ���/��R;��{�߹��{N�`��o��rD�n��H�r ��k����?�w(RG���v���y�=��W�ݣ����M[���tb�g>�:�2y��'R� kgΜ����	�#.�GDLNN�Ν;cvvv�\��p_��W��/��  Ɖ�; @�^I���|����׾�� u{���q�=�D��-���k]ĻS�ǉ�;@3m�	���ۿ?u�����kkk��{�y��D	"�-��ڵ+6o�\�������O��O���_O���Eĩ�!  Ɖ�; @�Lx��W_}5��O�ı����͛c׮]199Y����R�*����۟�܁2�H`l]���(����r�4@V��s:�N�q��}���� .�������q��Ӌٗ:  ��Qp ��+1L��:�'O�L��������o�N��K���~���I��b��Q�ӟ�6��S[������;@:�������1����ae�����o�,�J_��s�dN�8�:J��M  `�(� To5"�Qg�O��?��?����c�[n��&��y�[ry��j� \�,���ϥN���![ )���E�2��8ܳ,:�n%KU5|x�Su/�k�  �W�  i��:@��z���?��x�WRG�V�t:q�wƵ�^[ݚ�)�R���0p������O�� ������# �������=�<�}bz:�©�7o�]�v���dek�8z���k_�Z��Q����  ƍ�; @�����0���x��G�(��q�u��n�}�ݱiӦJ�����w�����|e�*� ������L�F���2�$/���������4;;��sO���V�6��`0�o|���|�}���R�   �� �4e�NEQ��?_�җbuu5uh�������cÆ���MLD�S����wMph��-[b��S� Zd������R� +�� V����q.�O|dPAU�fضm[������������_L�i��p�0 @�� Ұv��x����ǎK��믏��+����e�LO���4��w�����?�:�&y���N0V�dz{D�p��=��JY�ŭ�����'��4%�*o��v|�_�#G����DG#b)u �q�*  �1���S��_���"p�:�N�~��q�7��rނ���;0����|���# -�z�`� cei����c=��#{8)lݺ5v���n7uh��(����/~�l_�J�K  `)� ��jD8��
����7����7#���q�1fff�{�-[�����5��~�(����X��dLmݚ:�"�RG �� V��T�|uu�i�#�I�|vv6��XXXH����W���x衇�O�:�� ���ޝ��y�����e��C�p'%n")���p;���i��@�<-��E���&���i� AQ�E�E�hN�i�x��h�v9�DQ7�E�9��̜}���Ő#�8$g9������`0�9���HQ�������(�  �hI��:D��;wN����c��l߾]�=��������*Y\�}�L �K����[�e@�ԙ� ]S*��;?��	�ZO�f�:r����c����)=�䓺t�u�$��:   ��(�  ���:@�MNN�����~�ӟZG")���СC:p����h��K�r��+�o�	� k{��?S*��� !(�@��J��\���?}
��T*��{������]e}	p]:uꔾ��P(X�I���   \��  �[.ZH�f���{NO?��|���~�g~Fccc�QV�Yeҗ����Lp�x�ݵK�~�W�c H����� �	�﫺�����-��ĉڱc�u 2J��������?��� ���$g�   ���;  ������ŋz��'u���(���S��;����8�t��_.T�}&�@�����:��h0� ��T*)��|
�єN���~>|X�l�:`��ŋ�����I��%�[�   pw   ;�$M�Xd:	���ק�ǏkϞ=�Q(�˭�y
� �8�ٟՎ����c H���"�@�J�M�|�����5� JFGG��c�ixx�:
�u�fS�>�,��v�Il8  ��  `笤��ª� ЩS��������tE*��Ν;��c�i``�:Κ�ksԓ��m�7� I���L�u 	Pg�& t����T*�����3��~�\.�cǎi���J��A������?�s}���Q��#�    ��  ����)�I5;;���˿ԫ���V�e蘁�?~\?�p�6�2�������L��d��ܩ��w�c H���u H�b��0�ܜ�^oS��I����ڱc��q���ZG:�Z�����SO=��*�@�=   `$k   �q�$��TA���������h���֑��I��ڽ{�v�ޭT*eg�R���U��UR�~UkC� �c߿����u�Ο�� Ƙ� �U,7}���	��RU===:|�������lZG�"C}��z��WUw�ƛ.�`   �U��  ���f�    IDATLm��BA�������O��D�c�=�={�Ĳ�.�s4���mc
� ��\N������ 6��; tN��R���]����a����[��ĉڱc�u`�
��������c����Y   p�  l��:�K.^���ׯ��_��}����ᮞ��۷O۶m���i��U������k5� �6�ݵK���ҹ��])�� ����u H�vLo����2i'��)��h�������`Ď�yz�w���o��<�8���w   3Lp  ���.�V�z��g�����$%�D*��Ν;���'��.I����>^�v'J�Lp�����/��o$n��Lp��)
m�����^p�mxxX'N�СC����cX���q}�[��o�A����ZZ�  �&�  �:k�U�������+=zT��˿����H�����u�����ZGi�m��������<
� �H{��U�$]�/�E
�z��NhLMYG �Dj4j4m����S	)�KKC$���422���iMNN*�f& �gffF���
Cz�]�   �2^�  غ))o�Ua��ŋ�ַ��7�|�	(��|>���ڻwo����ڦպ��BPK� ��_��?��(� X�Z�W*Y� ��i���0�Zm�Vep
_e�Y�۷O'O�����u`Y�Vӫ���	��q�:   �˘�  `_��2����o���_�%;vL�T�:U�T��[o����
� �7^�װ9Z��K�t<Mw�Lp�D��ۿ�t�.���(��� �QsfF��a� �(�b�-�q�F��)��b��7�|S�җ��%�ر�:�l6u��i�:uJ�f�:>q�:   ��(�  ػ 
�P,��3�護������������5�ZM��N�>��Ԟ؂�6GC-Mq�x��
}_A��t.g �!;�74t��~�����eN4�`��i<�u H�j��V����F[�WkYÉ��F�\���W��СC���H�]�y�Ο?��'O��P�(z�:   ��(�  �;o +��y=��s:u�~�~AG��莎���:}���}��U��$���㭫J^�]Z��N� �m��A=��o���Ϛy�i�8 "�13c �]��%ɯ��v��I��(�Mn������0�����\���G��_��FGG�!ɂ ��￯7�|S�J�:V�	�   ���j   >N[��������Ok�������y>|�:��l��ٳz��ո�$����:��������x��U�l�j �a��=���i�?�'��7T�x�:��jRp��	ð�������jS��0�ŋ��G��ѣ�җ�����M� Ї~�7�x��O�#�hiy   F��   ��w%��QSSSzꩧ�w�^}�_СC����V�:s�Μ9��6H�ZpOe2J�r
V�Z�iUI#���UA�f �E[>�y}������_��j��[G1��i� ��Je�d��ry�{f�
�j���m���.]�������^۷o�b:$I����￯��{�b{||`   �u�  �$ݔ��:�orrRO=���l٢�}�sz��ǕM��h�B��ӧO�ܹs�*�'��.-m����^Q�
�G�{�i����T�~�75��˚��wT<�aN �0� �gqq����ն^/N�^p_ˍA��p�P�n�jUgϞ��ӧ�4��r�:   ��h�   DÇ���BA���N�<�'N�s����c!�&''u��i]�tIA���'������0����Y��O�=^�l `$�ӣ�����뿮�ŋ����|S�>�6��dh0� ���}������S��	/��o��jn@پ}�~�gV'N�P&��P:���ܜΜ9�.��D	t��    ���  �K�U�X�j��S�N����:q℞x�	���Y�BA�K�.�w���&�*I.�g�����%���Sp H:vLCǎ������bQ�'O�x��*�/�z���ss�t	��=
���0l�5]��N�}usssz����[o�'�Љ'400��t�� t��5�>}Zm��]��u    �Qp  �����q����ٳ:{��v�ܩ�|�3z��G��嬣���������i�3���l��$��K�]~�b 1ّm��_��_����y����/�2>���K�������\�_�*C9 6eqq����.�'�ߥ�N�.��������'z衇����ȑ#J������(�����t��Y�pZ%b�&�u   �Qp  �&A$��̌^|�E����z��G���|F;w��}_�/_��������}2�F'I��z&�Z�U�X���J%� ��k�'4��+>ߘ�^*�_���ի�ML�z�����FI�CczZ�Y� �ت��j4m�nP����q�a���A���	MLLhhhHǏ�g?�Y�������� t��u�?^�.]R֑�^iiI   �(�  D�YI���,1�ͦΝ;�s��i�Νz���u��1�%|S�%��Ӻp�>����l�޶�IRQ�^G�]�*JP��	� �M�ݵK��vi�_\�y�Z]*�_����v�j
:��
��h��Pp�M���vi�{,W�����	ð#�n�rY�N�һﾫ��ĉ:x�Y���`nnN|�A[O�D$��:    (P  DE]Ҹ�c�A�~333z饗��+�h���:v�}�Q����{�|^/^ԇ~�����<��y]y��.I%�N �\��  H�����O����w=���߸��v���Ǔ�R�O��~͹9� [a�X,v��.�3�:��knAh||\����f�ڿ��=��G�Rv���k�/^T>�����8k    ��   $�yQpO� 499���I����:p���=�GyD�\�:��z#��L�H���(]�Qp tYvdDC##z챻��O��7n�~���͛�OM)��#�r۶�w���٣�={T�qCs/�h�Ts~�: �V�T��)x~�֑��A���:B�ts������/��#G��ȑ#:x���t�r`�Ţ���u��EMNNZ�A��c    �  �䬤��:�����M�L&������:x���9-MMM��ի�|���K&�V���;)������T��t� Q��бc:����A���ܜ�7n�9;��q��ǵkל�l��eGFԷo��[n�v��ء�}����]aO�t���b"( l���bǮ8�}N:�'PZ�h6��p�.\����>>|XЁԷ��2�ǝk�W�\���u$�	%�m   �  �����}_�/_��˗%I[�l��Çu��!=��CL��j���ׯ��իW=BSJ;5},
��$�%5$�}��	� �8I��.��掠�����SSjLM�9;����Z�����j-,����0��۸"�N�gtT=۶�w�N����w�N��޽<��w�n��yJ��#�t(q|4)���x��jK�.Op���{q�S���r�=�Jiǎڿ����Ϻpܹ&|��e5�H�����   (�  D�I� ��B����{O���r��~�a<xP�����ؘu�Dh�Z�����Ą�]����Y�ahkUQ�l��7Iˊ��	� ���U���1�����rٽ��/�o}|g�9?/�R�Rz�s9�lݪ��[�UntT�[?�Sn���	�=ccJe2mϐ۶M=��j-,���q�w ؘ��Ŏ��|R��	�P333���ѩS���߯������ڳg�FGG�#�^�����nܸ��W�jnn.�k�0��u    ,��  3�nJ�c��l6WLw��rڽ{���ݫ�{�j߾}�t�\�4�jUSSS�����䤦��c3��jYG蘍��Iq�a�w ��n��u���6h6�-.�9?���rY^�$�X�W*�/��*��ˏ��E���f���hI�rJ��);<������;�2����z,34���Q�mSf`�:�$i��-���u3�`c
�BG�����Nߋ�����j5}�����%�.��JE7n��͛7u�ƍH9A���   �%�  ��(��>�ͦ&&&411!I�d2ڵk���ݫ]�vi���ڲe����6�M���innny�X,Z�ڰ��7"��"U(�"i��i���;  ���۹S��;��s� �_.˯���j
j5y���z]~�.�\V�j)�����x�T�$y��B�_z�Se��^W�Z!���m��R)e����tvxXJ����W��G�f��U$�Y�}��W*�UvhH�>e���Rf``�Ǚ�!��`��a����y� ;�JE���z��7��������p6��Ν;�w�^�رC۶m��ؘ��JeyMxzzZ���*����y�:    �Pp  �����b�����T����FGG�k�.���illL�v����a���@�RI��󚙙Q>�������|�&��m�m=6:�]�ʒ�$�ږ��|6�  �T:�4��VI����C�L�A"nV �nY\\����j��׏�ͬ�D]���<�[u]x۶mڶm��o߾�6�ʍ�q�j����5;;���9���kvvV�z�:��u    ,��  -�Y@�A���y�j������l٢��amٲE###��GFF"9ݧ^��X,�P(,�/�J*
*
��n~[�7��g3�\{����z{"l�7�  ֫��{���
���ZG�X�<O�[��tJ�x�=���wj�v"O�A���Y��ή�|&���А�lٲ�622���!j˖-F��v{�I�PP�RQ�RY^��F���&����q�   XB�   Z�=�W�VU�Vu��ͻK�R��������߯��>���-��߯��^�r9�R)��i�r9IROOϪ�f��0��qѭVK�VK�z]�ZM�z}���?��j*�J=b:.���v[v``S?����%�+����  ���	����)��-..v����j�~�e�n������rA|5�\nյ�;?��rJ��J�R���$e�Ye2IR__�Z���@�F�!i�����u��P��\^�sm��5b
�0�SI�  �
�   ��:��93�������򦮓J���f]��$o��7Yp�K�%eڒ���rY��ۭc   DF߾}J��
��:�����y�: D^�Z\\����OpO��(��c�c��f��f��b�h�v�:    >q��E   X
�4!��0)��Y�7��}}J�2��B-�W^��Q  ��t.����|�: �B�\�����L�u��b�*�X   �'(�  D�i�  �#��T*���#�7����8�I  p/��;�#�jQp�5���vI
j��<Oe6y�^�%y����i    ���  =�X ��YG��n������w  �����a�w x�V��J�ҕ�rz�{��Lp�)uIg�C   ��  ��	 �%}�T;6K����~~�6�  �$�z��X��  �����0��yn�������:*�kn ��$�|  �
�   �sN��kh��o�eڰYZ��9�^�l   rr۷[G0��=" �W�*
]{>&�'W��� ���    X��;  @��޷ </���k�fik@�  ���w�T��  �V*���V�r�=��	�I_s�n��   `%
�   �Ĥ ��?M�]����N�>L�  �[��uS�����|~���狒t�'�7� ���    X��;  @41)�����m�H��L5&�  �-�e�uS�	 ��h4T��Du�'��k�&�Z��u �Q�t�:   V��  ML�  )��m�6N�۬K�K   w�q���w ��|>������Mx�=�C% ��I�u   �D�   ��+~]M ��{;���$��v��c�;  ��z�n��`��; ���}���?���3mJEI_s�.g�   �n�  �)��� �K�4�vo�Ʃ2N�  �n��a�2�f�fSA�_ �F,,,(��?���t��I_s�.��   �n�  ��u  �� ����1:�����s��O�  �n�T�'�>S�`�0���`��~�f�Q�i�{QD��ް   ��Qp  ���� DC��L��fi\�@Lp  X]�u� �R�T��u�v���R��5�I�gI^o�.I�C   �n�  ��u�  �!�n��,�J�����Gq	  `u�>���� +��y��uyz�$�~�Y��� ��9�c9  �9�  ��#I��! �K�ɝ�,�4v'�VKA���  l���)��'�ժjFEs�Z5yިH��ǍF�:�h8e    ���  mg� ���R����\�,)�ȕۋ)�   wK����� ����.I��ܳ8u/J<ϳ�  ް   ��Qp  ���� �����$�a��  �ݒ^�{�� @���eÿ=�'���i�r9����6 ��c�    Xw  �h�;�  �%y�{��O�tg^�ơ�W*�   "'��g�TP�[G �HXXXPڝ�8\p�8p�w �nJ��  ��Qp  ���%�! �J�[*�L�
LIQ��c�;  ��:u�O\��@Ahqq�4�_���p��B�=�% ��{�   po�  �mQ�� l%}í���Q��{�G�  DU��{�hXG  s����}�4�˧��PpO�@	 k��u    �w  ��{�:  [I/��;�iZ��u�����   "�S'��EH����0��u�oJ�ZG�0�o� 	g    �F�   �NZ `+���CC�v�hOq�JQN  `#�w� `�T*Eb-įV�#�Iz����� $_қ�!   po�  ��5�  l%}�{�7M�Zڭ�"&�  �-��XG0���� �����uInOp��0�(H�Z�5��h�F  pw  ��{WK�L ���ԲN�v��H��4w  �U��޺`�; ���e�#r�����#tw �NY   ����J  ����! �I��[7��.k��5�B�:  @����Q= :/*��%�g�{b%}��59i    �G�   ޲ ���$U:�,��w  �U8>�]Ao��Ϋ�j�Fhj��p�=��)����u    ܟ��   ��c�  �$��ޭ�`%IaW�i�(�  �-�����# ��(Mo�$��[�#��	�I_k�@yI�C   ��(�  ��KZ@�AI�*Ս	��K���%�  �b��u �f��R�dcY��k5�f��Vc%�km �u    <���   �1'�u 6�>U������*_�*�#   Dw� �usss�V�U��}�Mx�=�km ��    x0�W�  b�u  6�>U����-IQ���W�
=�:  @��2���?��V��b�N8��e��2�:*�km �U�    x0
�   ��w� �H�T�nO����m�  Xs��0�N  ]���F��>�Z��`*34d�����ྚb�;  @,Pp  ��W� ���M�t��[oQᗢV�  ��J��u�|��S|����u���.OpO����N�QLp�vVR�:   ��Ub  �xy_Ҝu ݗ�M�L���S�f��
�   �$�����!�|^AXǸ��p�=;8(�R�1:*�km ��-�    X
�   ��u  ݗ�	�J����S��)�^1Ju{   {�㥳t6k �"-,,X�X�W�XG0���I{���~^�   ����  /oX �}.l�Yl�F�VN�  `���;��b~~^��[�XU�p�=��!��8+���u   �w  �xy�: ��sa�-cPp��w
�   +��(|�f�	� \����܇��#t��$ �ꊤ)�   X
�   ��w�F@���1�<�B���;  �J����O�	� ����;\pO!�6�I X�I�    X;
�   �R�t�:��r��n�y�)�-
�   +�Op�� �>�]��r�:�����u����8�U�    X;
�   ��c�  ���@�'k8̺^�w  ���R�:��L�u �|>�c�    IDAT���9<�=kt�^7y�g��Y   ��Qp  ���� �.6ݬ&�K�S�)�  �Ԛ���`*���\ �
�@�|�:�yOp�B�-Lp�4)�u   �w  ��yYR�:��i�������eŜ�;  �JM��Y
� ,��%ɯV�#�ISp�LoX   ��Pp  ������! tO��R��1:�z��r�;w  ���1���I��~� �q��.I��܇��#t��$ ��5�    X
�   ��w� tW�7ެ'�KvS�)�  �!�ZX�Na*�w 	���a�� ��0��¿CLp��#�    X
�   ���u  ݕ�{&��$���V�(%|B?  �Z5��z�uS.�'N��=���K�X�鴤���˜��Z�   ��Pp  ��$E���I�d��l�.<g�y�k5�g  ���ĄusQ�� �i~~>��%ɯT�#���){���u6 wy�:    ֏�;  @<Ŵ	�)I�,��� Ijhi�{��
�g  ���ի���FG�# @[������k������tw�9�Y   ��Qp  ���X �=I�x��t0���_*<+  @�ԙஞ�[�# @[�iz����tO�R��u��K� 	 wy�:    ֏�;  @|�b @�$}�-��)��cC�ԔT��s2�  `I��5���$H�Պ��v��{f`�:BW$}����X�   ��Qp  ���$�! tG�����������]|6  ��9^pO�rΔ�annNA�%L��{��f:Ʌu6 ��Pw�z  �&Y�    ذ���%}�:��sa�TfpP��E�������wk[��;\��*�9��ŋ�\���������k5y�ʎ�(��)�}�r;wj��!=��#G4p�RY��  iB�S}r�:����Q� �6�fS��X���̸Pp�P��Y� �=�X   �ư  o���;�&Ke#��Z�4 )Յ��T��5����UU>�H��8����97'}��򯽶�X��G�i��9��c�4x��r۶u��  ���
/�Qp�$���
�����U�f��6�	����T ��u    lw  �x{A��Z� �y.Lp�YGX��T�ԍT�N��"h65�쳚��wUz���]��R��E�/^\������)�G�j��Q>�t.׶� tF�j�x��us��ۭ# @[��ucz3���Dsa��e3Z:	   1D�   �~$�)���p.����r{�{����J~���VK����>��?Scf�k��ZX��ɓZ<yr�s�LF�,�����#��o�>�2��e ,i�̨61��Ą�׮�z����ON*�}�x�zwﶎ  m1�����W*�̸Ppo4� t���   �q�  �,鬤/X�Y.ܣ6�]�|-�E;���a�;�d�'?��o|C��	�(����UWu|\��?���tO�������C�o�j��A&��&�ժj�ML�z��j׮-���5�ժu�H�ݵ�: lZ�ZU%�%q/��7+�k3�F�p�K�   �q�  ��5QpυͷL'�KRIҐ:;��g�;��Tt��_�����u�5	Z-U/_V������߷O�w�V�����{
 ,xŢjׯ�~�[��U�~]��Y�x�E�@�����\��`ƅ�<.� ���    �8
�   ������:��r���)a�����|���b�t^������=�''��l^,4?�X��^[�P���8xpi�����}�!�?�����Q*�2��i��/�W��~]'�tD���� `S�岪1?���{vp�:Bǹ��@�tU��   �8v�   ��I5I��9 t�ӥ���Z���N�����8�}�y]������Q:�15��Ԕ�|s��S��z��Q��/�zH������ջw��==F����fS��7U�yS�����z��{?��8�� ��0��̌u�M	=O����e"�6�.�g�n    �C�   ��ޑ���A t��(o���
��u�����R*աg :��w����G
��:����U�~]��׵��w=����C|���۷����2��"h�Ԝ�Q��5gg՜�S��ծ_W��5n�t���(I��(�k�u ذ���ؗ��R�:��lDO�k'�� H�^�   �͡�  ����;�hq� ^�(�%���)��v�jɯV#�{ ���w��K_��u�X��EϜQ�̙��R�ݹsi�������Sߞ=ʎ��A��4y}rRͩ���>n��YG�:��ۧT&c 6$�%���\��`*���.��P(�9�   �
�   ����?��s\�|�Ơ�]���C�n-.RpGl�<��.��1�/՘�VczZ:uꮇ3���۳G}{������={�۽[}{��g�V�� �%h�����̨q�9=��~fF��7)�'L���� `�����y�u�Ms}���.���EI7�C   `s(�  $�O$-H��3\8>9�MԆ�&�wb�YkqQ}��u��@{�Ο�G_��� ���x~��ʥK�\����������;ջk�zw�Vn���ڥt.��� �"h4Ԙ�Vsvv�F���SS˥�f>/��uTt���� `CZ���c����8�,
�^�   �ͣ�  ���J���:��pa�-;8(�R�/r$�KJ�������l�|^��U��M7q��j����:>~ϯɍ�-���,�S�:����[\\1u�9;���)5fg�
�1A�����쬂�� �r�=��)��c��\Xc�g�   `�(�  $ǏD�H,&��2ez{����Q�˓T�4����|E��� Ї��j��XG�:4�y5�y�?��_ӳu�z�mSn����m۔۱��cc��ܩL�����E5�y���՜�WkqQ͹���Ԛ�[z|aA��[GFL<h ֭V�����|��١!�]A�H����C   `�(�  $�S���:��pe�-;<���$%JJ���u׿�M-���ut@kqQ��EU/_���e��W�o��{��Գu��[�*76���Qe��ؠ X.�7�����j��.�����z>��������TJG�X� �u�I��^�l��+w�H �{KR�:   6��;  @r\�4.�u ����[vxX��Y�h�侵���(�#�Jg�����u�k5�&&T��x�צs�����r۶)�u�r	�w�6���.��g�VeGF��+@R���V� ����o߼���Z��j-,HahXֻg�3�B �Q,U�V�c������p�Ϫ�&W�� ��d    �A�   Y^w �\����Q��,iH�{a�wDU�h����^�u	�M5gf�\�D��Ȉ��ß�������(3<����ǕJu�W�n�MyŢ�Ri�7���K�u�'�"9����  ���fcp��z�\p�:Rp����@ ���   ��  ��9I��u ��J�=N����EI��t=
k���v�u8�+��ҍ�����ae���W������Ko�=�������L����P�hȯVz��RI��)����j�U��R	�RY��Z�_��/���zܯV��뷮���;��YXXH�$l��{�%��-�es�NY�   @{Pp  H�g$5%嬃 h/W6�⶙Z�Ԑ�ۆkQpGϞ��'���<����T*�Q��O��{{�޲Y����J��O�+�J)30 e2���)�[�-y��W���ߦ��Ye��J���b�y
��{f<O��O�I���˫T�>n6ܺ�ίV�*���� X*�7��+���W*)\�� �c��;��}_sss�1:�	����	�Q�ii.	   ��;  @��$�����A ���y�}_�L�:JG�qj]Z*n�G�4���?�)�� &�[Ep��A 8a�3���  k633#���ct����7o&w �~d    퓶   ��{�: ��pa�{6���-I�6\���І� �s�O�D��q�  $^ߞ=�m�f ֤^��P(X�舠�P�jY�0�w 1Jz�:   ڇ�;  @���u  ���\'�KRQ�fg������+Wt��'�c  ����~�: ���Ԕ�0�����'��uMf�\X_uQ҄u   �w  ��yCR�:��sb�{L���6;�.�:�s��7��g  '?��u X�B��Z�f�c�r;�g����ɬ��k��^�   ����  �<��W�C h?&L�y3�"i���Z���l��K/)���X�  �[�x�: <P������Q�R�:���Аu��pa}p��Z   @{Qp  H�g� h?6��\p��EI�9���;��������c  ���А�}�: <��ܜ�����^p����Z���8�"��   h/
�   ��I�u ���ʙ�A���}�ڔT���o-,�+
�!����Rcr�:  �������fS�|�:F�yܳJe��1:.��ߨ8�5--�   AX5  H�9Ig�C h/'&L�R�?� )���e�;,5����e  �l���# �MMM)7s^Y<�\p��|-f��X[���u    �w  ����u  ���&\&�Gb�Z*�owX���UA�n  ����/ZG ��*��T*�1��+��#������rempL��S�  �0�  ���Z �^ͦ��fc^p���6v&�G�FO����/[�  �)�?��Ç�c �=A����]����Ȉu����$��&�C   ��(�  $��f�C hW6ᒰ�J�HU�	�0������u
  ���W�: �����Z��u�����|�� �i�   	E�   �BI�X� �>�l�%�X솖&��wX�}��Ο�� �s��ʯXG �{j6�����1���{B�b�^�[G �~?�   �Π�  �lO[ �>��45� )X��SpG��&��O�S  ���ؘF>�� pOSSS
�����?����u��pempHQҫ�!   ��  ��)I�u ��h4�#tE�6U}I멬SpG����T�r�:  ���4[4 ��P(�RY�d1���e�f��s?܁�yUR�:   :��S  �d�Kz�:��pe.i��Ik�5����.
Z-}�?��u  �4��/[G �U�����i�]�W�
�X�L��b�^�[G �^�Z   @�Pp  H�g� h&��W^R����U��� {�?��W  ����/��u X��̌|߷��u^�d�T�bV�������Y�   @�Pp  H��� �=(�Ǘ'��֯e�;� �<}�gf  '����P�\�: ܥZ�j��פܓ��W�� G�+i�:   :��;  @�]�t�:��se�Tvd�:BG��Tt���et��3Ϩ19i  '���߲�  w	�PSS��)�Sp;O[   @gQp  p��� l�+�p١!�Jʯ��(��む��  :~\C�>j �2??�̺�j|��tZ��]��q ��g    �E�  �?� `�\لK��(��g�#�*�
���^P��5�  8��� ���lj~~�:�)�\��`&;4�T*e�+\9p�ǒ�X�   @gQp  pÏ$�C ��6�2	>� )��㭅�nE������  pR��O;�7�c �]����{��|��ܓ��i�� ��u    tw   7x�^�`s\ڄ�I��/�~3�)���
ﾫ��1  pҞ��me�}.�x*
�Tt�X�|��K�6���$�  8��;  �;�� `s\ڄK�����{��l��݌������:  NJe������u X��}MOO[ǈ�'�gGF�#t�K�#	V��u   tw   w�@R�:��si�ǁ�ռ���o��w;
ј���k�Y�  �I;��?Rߞ=�1 `���i��o#�B�:���Аu��qix�`/��.   'Pp  pǂ���C �8�6�\8��Ҹ�Ok-,t;
q��'�`��*  @'��Y=�;�c V(��*8\��4�'�Sp/�V  �
�   ny�: ���@��Y��

�T����f>o	�W�����c  ऽ_����﷎ ˂ �͛7�cDG�+�v�\Y��(�	�I���!   ��  ��I�u ��F�K��y����E�0����U�  8�glL��տ�� +LMM9s�Z�ժ�?\Z�qe]H����C   �;(�  ��#I?�`�ͦu���8���I��Px�Z�_�Y�AB�����#  �#���ND_�ZU�Px�:����vIʎ�XG�
�@�1�  �!�  ��7� l�+q=���J���/�-,XEAU>�H��c  ��m_����+�1 `Y�����9���n�re]H�P�_Y�   @�Pp  p�_Z �qLpO�-��HRc��v�>SLo ��z��t���: �033�V�e#r�R�:���Аu��qe]H����X�   @�Pp  pϻ��Z� �1�L�riz�m-I�Eg�;�%h44���1  pJ:�Ӊo|C��ۭ� ��j��^k��[\��`�gd�:BW�a�@���:    ���;  ���� `c\�4�P*����u%IMI�|�:
b����F @W�R:����F>�Y�$ �,ݼy�:Fd�~͔����ct�+C#���u    tw   7��u  ��f\*��CGd�Jʋ�;�g��#  ��TJG~������$ ����37�o�W(XG0��	zά�����s�!   �]�  ��i� �ϥ͸�C��wjI��q�:����ŷ޲� ��i��?Ԟ�~�:	 �P�V��&���E�f�##����<�X��    �>
�   n
%1��!�6�z�d����i�j5�����^R�y�1  H����N|������i V�@7o޴�yN�:=�^�[G �q߱   ���  ��Z �~NMpwh��Ӛ��&''�u��̳�ZG   ���������g �2==�ԍ��
��d:=���ؚ���   ��  �g%��{ĔKӦ\����j6��������j�̨x����޽Gɚ����Ե���{����(�JDWHtEtEV�K$�I\�$q�Zf���4���ƃ"D.�@BPP�.CF��={�V}���>�\�սg�ww���>O�ޯ�zUwW��φ=�]������c  0�R)���������: �dkkK����1��ڲ�`ƥ��Kkj������  �1Y�    0�I���W[�{NMpw��.Iը���?k���8  �Q<^����ɗ��:
 �RZZZ���Q�#�Ѱ�a&;1a�o(���a�    ��w   �}�: ��qi3.��&덂z�j9yaaAA'BҔ?�Y�  ����.������=�� bmiiI��[�H���]��ڋKkj� Y���   ��w   �}DRU��c���qi3ΥM�Ea(�ZUnrRAhqqQgΜ�����uU���  ���N����?�cʎ�Y��;���T����^�^pg�;����$��  pw   ��%}Zҫ�� ؝v�m�o��n_{�Sp����-U�U�;��	vg�s�SĴF  �Y��9�x�+u�U�r�wS ��y�VVV�c$Jgs�:���C?�(���߭   �w   <$
�@b���S�v�_�\���Ғ�Ţr��Q"$��#�XG   ����:�������|�K�T�: ���Ғ� ���(��-��\���y�u {���&   8��;   >*�&i�:��c��;n<&=-,,����F��Q�����1  H�TJ�S�4��h���4�i�[�U�,[' �g}}]�z�:F�7��vJ*��ؘu��i6�� ��'$qD!  ��X�  @KҟJ�A�  �Υ͸�А2�����_�s�M�F��r����)�DH�ړO�[_�� @�;��ŋ��>_��-�_����u4 �g�VK����1�V��]�VʡS�\���   �w   H�E�H�6�r���J喟_]]�qr<    IDAT��Ȉ�����I���#�  0uS����T�xѩ	� ���E�u�D��kod'&�#�U���% ��%}�:   lQp  �$�����Q�  �̵͸�Ą��l�D�6��a�T*�J��}N���<��u  �"���;Ev .[YYq�b�^rz����u��rmMH�OH�C   �w   HRKҧ%��:�;sm3εib�
���n������'O�1�.
m}���1�!���׼F��E�/_V�TR֩  {�V��9ϟW��y_�����9e������Z������v��ރ.�ؚ�kkj@�=d    �(�  `�E��=��E�R��u��pm��Z���cssS###wl�n���
�M��0����O��Տ#�WsvV�+WԸrE�������vA ����#�tI�3gTܞ�^8}ZC'O*ŉ5 pK�NG�1��ܴ�`Ƶ�܁�ؐ�)�   �G�   ;>"�.i�:���P��ihh�:J_�v\������>fiiI�bQ�\��wկ|�:Bl�x����8��j��%_�t��C�S�g�e����Z|o-,P|��MN>;���yΝ�ޞ=�4�� ��DQ����RtO�(RP�Y�0��P
�@b|BR�:   �Qp  �����)��w{  [�vۙ�{nr�:��Z��H�ô� T*�t��yg������?n!�:��Ѯ���5���j��Ͻ���5?����33jLO�93���̮.> ��i�S��iN�V�̙g�?w��������h4�c$^P�)r��V�~6Sp��   �  p��w �Z���لtm��Z��+h4�����fSkkk:z�h��!���	��N|��+����s������p�_��U*�q��W�\}�93��	� \:�W��ћ
�ӧ5|�҅�uD x�FC����1�_�ZG0�w 1�&�S�!   �  p��J*K����\ڐ�:��z�N�rׂ�ԝ�722����>�B5�����1�R:�W�Ȏ�kt|\���u�;��枝�>?��������dH �q�)�ӧ�;t�:" 8-C-,,(�"�(��x�ݵ5��Ӏ�CI�u   �w   \�#��^k��!�wl��F~�*�:��ǖJ%]�tI�L�S!�jO>i!&��T<��k�s��S�oz�Z�R�m~���{kaA��$��ؘ�N����^<sF�3g4t�ҹ�uD �m,,,���X�~�b��K��u:�\t$��X   @|Pp  ��> 
�@��Tpwm�؍:���~���ZXX�ٳg0�����b��?�'�n)��k��E_�x�}Q�[Yy��~C	���2H �R����S��qN�����:qBC�|���a  񳱱�-~7�)��QΡ5��Ҁ�����!   �  p��)iY�q�  n��n[G�T>�L���эȽn��j5��eMMMP"�U����������1�,�Nw˧'NH/y�M����Z���KKj--�����Ғ���j--�S.�`%75���G�?vL��'5t�x��~�
'O*䈔N[� �X����ʊu���qx�{vxX)�Nm��$��K��C    >(�  �F��?����A ܚk�r��	g���l_YYQ�XT�X<�D���������_ٱ1�=�����ĄF_��[�z�������Zw|�����͙�F�Sثt.��Ą�G�*䈆�U��i�y�s'N(3<l �ga�T*)C�(���a�Lv|�:B_���$���    ^(�  �V~G܁�rmS.;1!-/[�0���q�Q�T*��ŋ�d2�
q�Zj/,X�0w仾�:��t>����*�>}��t��g'�_����-Ɨˊ|���w�s9e���9�};vLCǎu�[G ���ҒS'���_�ZG0������W���	�w��  �x��  �[���I筃 ��k�r�m�^k?wI�t:ZXX�ٳg{�qԸrE����iM��e�)b+75����m��KR�n�[[�:	~g����ښ�jU���qb8���NV߹͍�+�]^ڹ��a)��� H���U�q�v�sy��ck-���	�a�    �
�   ���H�)� n�ڦ\αM�k��Pd��jZ__�a&������̍�7:W�����]'�K�'�����.o}�[~/�孬toWW�)��˒�^ Qr���MN*�}�����������䧦�ʲ� 8X�fSˎ�f�/.Opwm�ŵ�4 a"I�  ��a   ��>Qpbɵ��].��w�����U�E�(�5;k��!���M�PP��Y�vBD�+����P�RQ�\VgsS~�rݭW._}?t��F:�SvlL��1e�ƔWv|���������S� 1�J��"N�90Q��ڲ�a&;>n��(������[�   @�Pp  ��<&�IIϳ�z�mʹ\p�k5E���)�Q�T*��ŋ�2iv`�WV�#��z�K�#�F��G�(�Ȯ�H�ju��ժ:ժ�jUA����[[�������s���e�o��Qe����)�o�w�~�X�� �=[XXP�ӱ�1��JEr���Z\[K��   O�n  �N��[� p=�&��vl�u�H~����Ծ���}�������J�R=��h//[G0���s�k=�.4t℆N���[-���F�[�o4���
�M����Z���A�!�VSP�)�<ͦ�fSa�s�¢�^?��� J���$e�ƔR�XTfdD��Q���ǣ�ʎ�(]((]((7>�t�ؽ�X��ٝ�9u ี�5�j5�ϯT�#�rm�ŵ�4 AI�  �x��  �;�o��/Ii�  ����)׎;Qgs�
��l6����cǎ�(��[]��`j�E/R*���cW������Z��u��ͦ"ߗ���-�7����$IQ��.�G�����A������h(
��;�����Q�l�����l̎�*���W��Ȉt�����2����(3<�T*���X�y�ƤT���LF�bQ�\N�|^�!�r9&� p ����֬c8���i��kk-���	���C    �(�  �Nf%}N�ˬ� x�k�r�M�Q��ʭ���X,jl����������������+�   ��T*)�"�(N�/��[ka�;[�   ��b'   ��� \ϵM���uS��*���(o{�0�_�(t�{F��<�   �=��H�RI��[Gq��x�=�X��y�ӑ ��K��u   �w   ���%5�C x�k�S��2Ţu3�,�A�R��0{����r|z�$�>�9�   �{����F��~��k��
J���1�ʵa@B|Lݒ;   pK�  p7[���:�g�Vp���c�Ů��M�V������>'�x���Le�Ǖ?v�:   �o�jU����1���w�X\\K�}�   o�  �,41�⦜kGg_� ��U*���?/�/�լ#�*^�`   طv����E�Nry���k,.��1�(��!   o�  �$i�:��v��(��c�����;j�}eeE5��у t|��p�u   `_� �����0���$
�n�����K�    ;   v×��! t�a�N�c��\<>{�Am�GQ���y�w Ϗ��m���(�   ��(R�T����(�_�Z�0��w v�c    �G�   ���  ����\v|�:��R�hb?�/p�{������    ���ʊ���ug��B߷�a&���k�h@�����e   �G�   �����[� ��vlj����vDA �V;��o��Z\\<����r�����    �I�RQ�\���4oc�:����u�������Y   @2Pp  �^|�: �.�6�rn�^���y��_�V���~�_#t�b�e
�   ���Z----Y�p�_�XG0��)yQ��<� �|I�  �d��  ��x��� ��Vpwm��F��%ieeE����:���Fi
�   H��5??�0��8����̵5�������H�(I   �
w   �ł��Z� @��5=�}���S�&t���4K[   ��(�����N�c�:�Op�MLXG諶�'�1��    Hv  �W� ���{nr�:��~�&��ZG06�   ��Z^^V�^���m���<�\"�l6�# �*K�}�   H
�   ثJڰ�ε�{*�Svx�:��~n���m�J%EQԷ���KYG0P  @�mllhc���8q���)�.�c�܁���$Ǐ"  �^Pp  �^�%��u�u��%){�u3��|��jZ]]������VL��O�   1�h4���l7p���spm��54 ��e    �B�   ��� ��\�>�����`�S���k���3e0���^�YG    n��<���s:V����"���
w �Fң�!   �,�  �_���u�eN��2��7�.����:�c���{ka�:   p� 477� ���:_̝wpm��;�c    �C�   ���� ���9��&���ӣ(R�Tr򂊤�
�L5gg�#    ��y�y�u�B�y
\S����x.��1ӑ�^�   H
�   دߒ�N`��±��h�Z-�F�Ah~~�Ƀ1�v��ޘ���    \gqq���b�������$-Y�   @�Pp  �~-K��u�U�f�:B����.�n�{����yEQd���z�ݯV�/�    >���T�T�c�:������ 
�X   @2Qp  ��x�u �U.Np�;�	{-�o�����i�,�us�˗�#    �V�Z]]�����~mm��	�.��1�,�#�!   �L�  p/�@҂u�E.N�rq�ص:�T�T���n�:~�:������    ǵZ-.N���i]<��54 F~W�o   �D�   �"��߭C .rqs.w萔JY�0���$����Z�Z�����#R���
w   �}_sss
��:
v�	��pq��P�;�C    ���  @/<��B%�>j6���.��*;:j�L\
�����8Je2�>l���W���2   �a���Y�>�i�"N���-S((](X��;�/ 3%�u   $w   ܫg�]��G�nι8ilG�6��0��ܜ<ϳ�ICǎYG0�om�q�u   8&�"��ϫ�n[G�x1zm�o���4����e    �F�   ��n� �k\-����`&NwI
�@sssL*����#�   ����E��u��#?f���)75e���kh��uIY�   @�Qp  @/���5��K<�S�1���icR�
�R����ܜ�0���<w����   ����U*�؇8���W�TZ��u�EI��G   �
�   腎�Z� \��]���XI�lnJQd�&�VK�RIQ���p�usտ�k��   �Z__���}�M�u3���;�    �(�  �W~C�F��\<b��{��ȯլc�R�V��Ғug_�d�^�����)   0�j������c`�:�uS����u�5_���u   $w   ��W%=jp����ԔuSq>J}ssSkkk�1�4r���ba�ӟ��   ��l69�*�:���L�84 �"����m�    �  �K��: ��Xvu�؎8�%iuuU��,�Uvb�:���Gq��  ���y������u��'�:d��Z�� �U��~�   �  �K���N�G.Npwq3�ZI،_ZZ��֖u��w�usa���?�S�   0AhnnNAXG�=��E��š.����T�  ��@�   �Ԗ�A��+\ܤ�NN*�v��l�SGQ���'�}Z��~�����OXG   � 	�Psss�<�:
z��;w ��   08�m   ࠼M�5}��&]*�Vft�:��$Lp��%���yJ }D��k�_Usv�:   @E���w���r���)�.�c�]�Ѱ� ���l   ���;   z�	I�X� \��&{��!�f�m������Yu:�(N��-����Y�   � X\\T�^���r�����vIj�Z� ���u    
�   8,d}��&]�Ⴛ����N����Y��oe��<�yJ���1ba�U��>   ܃��EU*��$]4�kYG�R\X���   ,�  p��bt�ݓ��x��477�0���t>���?�:F,��V�����  ��ZYY���u�Z���E���G��ߕ�Y�   �`��  ��Б�;�!�A��&��w�VS��X�سV����yJ�l��/��=$E�u   $L�\����u�����k��Ąu���}Jz�:   w   ��J�C ���M���u;Q$?�����J��"J�f���#�F�����_Z�   @�T*-//[��I�k�^a�;���.[�   ���  ��2+�ϬC ���hXG0�u��.��ذ��o�ZM����1���^�T���s�~�u   $����U�W.[G0��ZJ�ղ� ���   0���  �Aba8@�n��ݔݑ�M�J����%�);6��K��c���׾��/~�:   b�Ӧܐ��{!��wW�΀>Z���   L�  p�>��$w ��M�����;�ؔ�����ښu��4��[G���w��:  @|E��JE�R���� �V�N�W�fS����0���Enb�:�	WO?��%��!   0���   0�BI����A�A�l6�#��ML(�N+
C�(&:���zbuuU�tZSSS�Q��K_��}�:FlT{L�<�C����Q   ����_��jO=���O�1=�������[>>=4��'T8sFc/x�F��|M���ʎ��9��j�ۚ��S��kK���Zz�\������'��_�  ��E�   ��%����u`�8;�*�RnrR^�l��� ������N�599ie`L~�*��+�<�(�1����|�K�Js�!  |��5._V�T{�)՟zJ�RI�Ä��VsfF͙m<��$)��j�4����}��*����=���쬂 ���>����)�.�c�����JZ�  ��E�   m]�H�Q� ��i�Z�̸\p�ئ���$Qr�L��ɗ�D�G�������'?�c��}�Q   z&���x�iշ���˗ո|Y~�v _/�}m~�K��җ4������_�ӯy�ƾ���$��433#������\]C���R��kg@��:    w   �ïIz���u`�A�N��\.g��o�Z�]�����N�5>>ne z��(���7�I���[��~�w_����U<{V�L�:  �텡��W��7�~Z��]���=Me�i$���>��O}J�^�2������^`�e�:��fgg)�;��ܴ�`��5&��˒��:   w   �×%=*�[�� ���l:Yp�:d�Lgc�[dI�5CQia�{�1%�{w�;�SO��-�1b%
C5��Ԝ����Ϯ~>�ͪx/]�ȥKy��4r�}*�:5P�� �d�U5�\Q��5�\Q�'T���S�	�?��Gѱ��^]�������r{�ӱ��>�<O~�n�L~j�:��F�aT�a    ���;   ���E��f��d!8Υ��v:
�ueFG����N�=�Jill�:N��:��K�Ըr�:J�E���v�l��g�ǻS�/]��s�������}�)˿M  ��rY�+WԜ���.2=���������'���Oh���s��&��o�Nt��577'����7�'��Evb�:��V�/�,�}�!   0�(�  �_> �%��W�Z�;<�]�n���.uK�RIgΜ�� ���i�;����=�UU{L�����CǏ�xႆ/^�ȥKW�w�T	  p{���n���g�}�rE~�j�@t�e��O��μ�u��?�T&cI��fgg�n����H�񂻫�W<�S�1�A�I\=  �G�   ��;��笃 ��Ղ����;:岊g�Z�8Qi~~���=:��߭��1L�����jo�+    IDAT//k�_���ى	_�x�[��N��R)��  �/�P�RI����+W�|�5��4���/�4����~����+��L�h'���Pnw\bOG�WO�su�8`���Y�   �(�  ���*�g$孃 ��գ���ܽߜߙ�~��Y[�I���@�s�Ԝ�����RQ�+_Q�+_���b�;���/^����tI�3g�ʲ, @����Z���McoNO�1=��������뫯�����լ\�!��!��{nj�:�	
�������   p;i   �%I��j� ��pu�.�������u������(�߃c�x�f��N�N�M՞xB�'����lVųg�+�o�Ӆ�QZ   IA���5E�����O?�V��(��%��׾�����Z/���Pfd��_{����E�ޠ_$~7C�����f��Z   �;(�  ����(�=��f]fdD��!�N�se�\�����ٳgU,��$����
�1�����u���R:vL�s�T<{V��g�E�s�T8sF�<��  ���5?�����o33�����jO<����O���v�����5w��^��\�H��R)e�NQ��.@�=)�O�C   ��  �o%�I�f� � py�>75�`q�:�	�J7Ahvv�I��P<^��{�jO>i�Ej//�����G�������/^��}��p��շ��� �-x���)���j�Jj�Jj\��������Qy�1}��o�s��kQnǭ���F��q�r9�&�> ��ۭ   �-�  `�m��k.o�妦�r�����ajnnNgΜ��Ȉu�D9�=�C�}��ժ��?���_G:��M|߹:uJiG-  ���KK���|�vnN�����z�uBl[��'4��:��;ԏr;n���a�Lnj�:�� =U���   pw   X���7K:cH:��[�>l���X�]�U���)��ѱW�B�>�(��� ��Zj-,h�_���tZ��'������N)�ey o��U*�97�l�}������ӱ��]z�WU���*�?����@333j��=n$[�騳�e�L��!�f��u`��[�Q  ����  �_һ$��8�x.�so҆���VSft�:J_�Lr?}����Ƭ�$B��QM}�wj����:
���Z��Z��6>����Je2*�:��ٳ:sF�ӧ5t���۬c�c  v������ו�WV�(���=O_��_�7��o*�N��y}����,�v�Rgc���!9����f���   @_Qp  ���J�YI�����-�<�]�Nq/:X>��H�R����|��)�㖢 PsnN͹�[ޟ���Zv/�:����ݷS�4t�ҹ\� �*h6�^\�z������E5K%���uD�I��_��G?��zUO��r;���Ю��p 
�@����y�   pw   Xٔ�AI��u �\>n��MZI���U<w�:������S�4>>n'�&_�RN�Tkq�:
ƯT�U�h�o����R��G�^-�_[|:qBCǎ)�e� \�ZW���ś�읍눈��w�SǾ�������t:�����y=J�A�Y_��`*?5e���C!��5�    p�L   ���%��zw.5���Q�|̶$u�BE�E�&&&���Z*�։�AM���Q0@�0T{yY��eU{�����9��ɓ����:qB���ɓ��� ؗ��P{iI�[Naw}B2��[]��C���^���܎�r��S�Ⴛ�C!�zDң�!   �&
�   ��w��L�wY���iT.O!�(�Kݒ���TrJ�wv�~@3�|�� ��W����y++�>��-����Zx/�<�����	��Ç�T����=a�}��%oeE������r����"�V���S��t�5��׉/��inn�r;v����y�O�sy�衷Z   ��(�  ��w`�\���Q:�W�h��s����Nr�����[��Gu��/�ڧ?m�ʯTT�TT{��[ޟ��?rD�c�4t���G�>[~�~?��R�L��@rD����G�׽��n�}eE���p������|FG��?�۟�<������J�A�|�����\^3zdF҇�C   �]�  `���Nr�u �\?n9?5��Ғuܯ����05��d�;9��?J��v:j-.��}R�-��:rDCǏ+w��
Ǐ+������S�������>�Uykkݷ�իﷶ'�����)���uT��?��=�[��fggp*�������Q�r9�f��ܳwH�I   ���  �8x��_�$Q��VEJ�R�QL�.��>��V�����=j%��_�B�������_[Gz'�^YQ{e�K���=ڝ�};t����G��Sp ���ݾ����)�_Sbo//+�׭�����cj�̨x��]�h44??O�{�r�=���܁{R���Y�   ��(�   �%�?H:iH�(��j�T,���py����!E��������� t��	�(�t浯����k����*��*�����𰆎Snj�[|?|���#G�o�+;1ѧ� F���Pgc�[T__W{eE��uy��j����]^=�:-�7���.��O��1�ZM�RI!�`��NG���^3�(���=���C   �m�  ��ߒ��� I�r����ڰ�QgkK��q�(�����0u��IgO7���/�
gΨ5?o����PczZ����c����9��ؘ���W'�g�Ʈ��WvlLyN� R�n˯V�NY�����W��?�VW���P��i�&+��.���R:}���ժEQ��ax������P ��;p<I��:   @�   q��J�I��A��i6�:t�u�Ç�#����)��F�RQ:}��ҷ)�8)����=���X'ϯV�W��zl�PP��!�V��!�&'�S�VnrR��I�''���辍�+1`!h6�)�孯���)sS�5�������:�:�ln*�}��@�WV��裚��o�龍�---� �66�#�rz(@��D`�~_Ҭu   ��;   �bC��J�	� @Ҹ<�*�h��W.�x�u�ت�j���י3g(�_��+_��w�[^�lpF�j���������d��)���+;1�����s;����n9~|\�B��&@�Ea�`kK�JE~�����(7����!E8�����M���u���% ����w��ʀ{Ib*   b��;   ��%���r�A�$i4�̸>�������u����ܹs�d2�qb!](��k_�g��6�( n#
y��ϧ��n*�gGG��ގ�<{;>~���ϧ���o�M��
�[[���Bzp�b��ǝJE�֖��-�� �h�/�BA����$ieeE���Ʃ0ڎ�;r����Zp�>#���!    ��;   �eF��$��:�$�V�:�����;�o��V����̌Ξ=�\�k�$��?�������ܴ����v[���9�6��>[�S��b��%��Ȉr��J���
ݒ�А҅�������=��!�fSa�y]1=h44��k5������f�[X�yL���^�_�)l6��8&h6�����x�������葎���\pg�;�o��u    `w   ��/I�AI)� @R��u�f���J��Ζ���{�v��$�|>o�\fxX�_�ZM?��u 1��:��=��%32�-��ʎ�t�����+��w�
J=�~>��ؘ$]�X��������J�rR:���H��+�e��&a(�V����������n����z����uEA����NSo6v:
[-����^�ZV�)�+�,�� n������ߨ-Na@�^p�;<�	���|Uҧ�C    ;X�  @�|I�Ò��:�NO�J����Rki�:�	&��M������Ξ=�"��u�~H����J�:
�����t��2e�-�g2Je��KR��N_}|�PP�6=��������rJ��=�)�� �)�_�qp��W�;v:
�)�G���R�	%]���u���Ջ��^�~͜���+	��Z��f    �w   �ѯ��;�k�O�ʹ\p�ذ��8AhvvV�O����4`We��u�u��3o�u �(�W��t� o��5I^h�_����n�H .Op�NMYG0��i��>�$��u   �Z�?   軏Jz�:���>r�+��(���8aj~~^����Q̝�������1   ࠎ�I��Ǜ���a���;��5y��Lp���%��!   �kQp  @\�� @R��i�?|�:��(ԩT�c$REZ\\��ʊuS�|^�~�ǭc   �1mI���IW{�)y��F�0h<���Kn��H� ���n�   �
�   ��ߖ4kH׏]�9>����n!���׵�����I�ǿ��5|�u   8�)iMRp�Q����G<�_+g>�N����oJ�Z�    nD�   q�Kz�u 	\���z���M�^�T*���S��QL�2]x��c   �5u���͛�;z����C���Ppv�.�-�!   �[��  �8{P�}O w���]��M[o�o��P��533#�����8��k�[��:   XE��]Ӝ�U�T�G8��Lpw{�؃��=   �w   �YK��1��/�;�i�K�VK333�<�:���~�g��f�c   `�D��%Uw���/~� ���/�>l���ke�.y�~�:   p;�  w�&i�:g�z�:�������u3�o����y���vr3|��%�����  �JZ���YʕG=�4p����>���2`�>$i�:   p;�  w��k��f��(��c�I��w���6���@333�Vw;crp����P��Q�    ��I�=���ܜZ���.�8\p�
���1L�x�:�G���  ����  �$�e�}?pF��<�:���Ó�\޴?HQ�T*iuu�:J_e��u����   H������>�<S�qO�H^�l����%���˹��>.�k�!   �;��  �$X���u �\߸�;�y���
[-�kmmM�RIaZG�c�x�&�雬c    ���$���_�b���E�֖B��>�n���d�.0�   �G�   I�K���Q`���q�?|�:�)�)��Z�jvvVA�ȏ�TJ����)��Z'  @�T$�K���C33j//� \䭭YG0�?r�:�)��������	.�s�!   ����  ���;Il�+��o޺�y��fS�����8|�N��Y�   @BD�۫=|�ʣ������/�9>��52`~�:    ��  �$?�{�f�i���޼���4==�Z�f�/ο�*�=k   1HZ���J�&w�����FB���/J��   �nPp  @�|E�'�C q������:�o��S���W�\��r�2Ţ�ޛޤT��#   �ZGҊ��<w��y����t�/w��;ׇ@ w�    ��%   ����=��5\߼s}:��+�"-//kqqQQ4�?��_�"�����  �j�[n��k0���w��H\���>f   �-
�   H�/J��u n\߼K
ʎ�X�0��潕��M���+C�(��ߨ�s�1   #[��$�o�
���/O�����Na��52���  �D��  �$��b�;p6卵������j5=��3j���QL�P��{ӛ�4�H   ��$�%m�?3���V��2����s��J�r�1L�~�!p+��C    {��$   ��Ie�6嵐�G�#��ln*
���<O333��ڲ�r`�_�B�}��c   �P iUR��_4����c���H�����j�1����G����R@R��  ����  ��z�u  Nؼs{���P�r�:�ӂ ����VVV����ox��x�:   �%-o��[��;����rG�XG0��&�%=d   �+
�   H��H��u .ؼ��o�z��� i}}]sss
��:Jϥ2=��~I��I�(   裺��ۭΌ�=�^�b�:��6r|mD���u n�,i��   0�(�   �~�: l�Qp�8>�.Nj������y�u���;����Je2�Q   p�"I�����m���&@�x��6�:d�C ��\��>�   �~Pp  @�}L�Tb�N��[G0��xi�ۚ��V�^���s���mzο���1   p�u��׬�l�<��v����9�/��4��Á{�1�   	E�   I��� q���]�RGAhnnN�r�:J��+u��~�:   @[���m\T\�,��#)\/�9~���Ӓ�e   �/
�   H��H��u��wRvlL�|�:��7��*�"-//kaaAa8X�.���s��_Z�   @�՝�X������׿n	����Lp���u .��$�:   �_�  0���Z-E�O�K�����Na��M���T*���V��9�����_�ox��JYG  �=�$mH*o�G�����p���t>���us�IҌ�w[�    �w   �?���u�R�j�Z�1��>��[_�\��!���fffT�V������/��_���(   �_Ҳ��u���|���wQ�N�l��L��.>w`ۛ%u�C    ���;   �/X �����������ڲ����@�RI���u���.=�ۿ���﷎  �=h�[nOB������u�XgsSQX�0�s�T�k�>芘�  �@�   ��c��h����wx��$uVW�#`�6775==�N'	U��y�s���ާ3���Ki��   �,�T��&)4βU���<�_9|���v��0L�w5�@�Y���   ���   $Lq�Ӛͦus.Op�����I�j���3Ϩ^�[G�t>��?�S��~P�^�2�8   ��@Ҫ��u�}�Pp��^pg�;� I�%��:   ��  0H>.���a�T�ݯ��w�7�(���jee�:JO_��ox�[�>��o��8   �֖��}�D�'�T�k_�F{�^W���K�I�(��  `@Pp  �������<H������O����s�G�"=<Z���UQ�.�D(R'T�
��ǔd���� q�;��f3�8)(pT�NcS(R�yĳ���Ν����}��>�䏞陹w�ޙ{g���������<��w���s�?�&��7��upp�����}�Q���>������}���Z��oQ�T2	   �ZLn�My
a���˦c`Dy���F%ggMG0��;"�MI�b:   pU(�  `����ϛ��"����V̊�[ݨO�w�mkmmm"OV)��z�����������~�r�=g:  @$�*��B�Y�B�K_2#ʉ�I�)
��~����  0A�    ��G%}�t঱�'�	%�e�ժ�(F0�}�y����u���kv�	V*��~P���$�=8P��W�~�55_yE�k�E��/  �u�I�J��}�Z/�,�������E�=q̲���1�8�? �^��  0a(�  `���?��u�� 7�E����ld���E�	�����d۶n߾�Dbrߤfg5�u_���;�����Q��W�~�U�^}U�oȫ��  ?�����&cj�I}ۖ��ʿ���(!���c��(�K&M�0���������  ����R   D�'4(���DdPpH��J_���F��/�Z�7�سm[+++�}��
���87&����Ғ���_��o6�YYQ���~�5uVW�Y^V��  �&_ҁ��'U�O���;N�� 0Ø�$�G�eI�e:   p�(�  `R�{I�����
�Q_����Sp� ��kssS333ZXXP,�����J�{�J�{���WwcC��^�����ʊگ��   $�+��A�}����e雿�t������F���LG	LpGD}RLo  ���  �I�II�d��
�Q/w������n:�X�ZU��ѝ;w�J�L�	�DB�^P�N���﫳�*{yY��^S����Y[��4G  0�BI�4�H    IDATI-�AnH{yY�m+�ϛ����홎`T�O�?±1D�$���   �u��  �I�ǒ~G�_6�	L�HG|jY/����q���iiiI�R�t�����Wj~^���x����,�+_�����ʊ:��r&  x�X"��[�28�������j�w~��s��$�Fj��ʩ�|�6�R1�������;"�M    �w   L��􍒒�� ׍E��d��nķe�t��kkkK�v[KKK�,6)��x6��߭��}��~�%��=uVVd����++r��%  Qu�Ȟ�sG�Ýjro}��;�8��*�ے꒢�WM��_����������qLG n��ux   &w   L��H���K�A��F�} E��t܀F�!�qt��me2�q�V�XT��P��8u�W�����Y]UguU^�f()  ��\N��S���%��W��畽sG��ɋ��w�}�Y���I�����/����E|�;��v�m:pSBI�4   �N�  ���W$�M��mۦ#��x6�D.�~D�=
����������Y���)���41���*�ר�5_s��~�9,�w��e���������� �sS �y�ҰȞ{���4��S��-�)_��>�����EYǕ[�ʹ_�۷MG�p�>�}~�t����1D��J���   �u��  �(ؐ�����t�:��+��L&MG1.97��Ɔ�Fx��B�S��"!CU*ٶ�۷o+�J��4���J�}�J�}��ϓ��'{yY�������Uu���w��� ��K$�^\T�ΝA�����{W�;w��s�ʿ_�T*j��B���GZ��B�
z=�[-�1��g2���c�
@ҏ�   \7
�   ��OI����� �u�v��%�ԍh�]a�^�2����v�Z[[�����8�c%��E�~px�mo���������KowW
C�� �E�,K�%e�yF�g�U��g�}�[�{�Y�������8��߿�^���K/Ezת�گ���}�t�V*�~m�ZX0adt�w��I��!   ��F�   Qq_�/H��� �ɶm�J%�1�K�͙�`���O�=�|�������nݺ�x<n:R��,����_{���;[[�޻'gkK�֖��  DW�T���Nc�ܹ��s�)������ժ���xc��y�j����\����k
�P�X�t��홎`T:��@�x�'�uM� ��+�GL�    nw   D�ߖ�m�fM�[1D}zY/��Q�j���tt��-�E�qp��KR��TwsS��uu���ln'��L$ ��ųYe��N`ϼ�-�>��r�>���(�y��߿�D��������m�Y_W���LG�A�J�t���%1���K��4   �	�  %MI�Pҏ�\��>����7����{��ijjJKKK�,�t$\B�TR�]�R�]�z�1�Z�s��`���k��=�ժ��  ��XL��ye���Hvt�޽��̌��h4���+���|����*fY
������֫�Rp�87�����#��> ��   "��;   ��'%}����� ׁż�T�w{_�ǱF��N��۷o+�˙��+���QrfFů��\W������A�}kK��uVV���QxNA �qb�RJ��K�J��=�x6k:�S�}_���j�Z�|^�XT����YY��d����+Z��o0���,��@�pL�ӒvM�    n
w   DMO�/�gM��yQ_܍��:��y�666433���9��O0+��������~_���CSߝ���ܿ/�� �Q1AS�/��ji{{�ܩ�*��=�%�o������MG�!Q?�;��@���!&ܾ�   @dPp  @}Z�Hz�� �Uc1o�J��,��5���A�
�Pj�Z�u���#(�H(��3�>��x��l���Vo{[���������Y  .#��>T\O}|���T�t����vww�h4.�y���j���o_S���;�:++ʿ���(0īTLG0*57g:�H`�&�ߓ�6   �I�  E���-�L��y�Rss�-��m[~��8%f<�u]����\.kqq�i�J�J*�J*��ҙ����JE���`�������ˍx� pZ�TRjnN���S��SssJ��+s�����9�ͦvvv.<�����ަD.�>':�����#ʷ�H�H���?�11L�5I?c:   p�(�   ����?���A���bޱ���1�q���}�Y�10����:���qaV:=,'������m[����)��﫷���ޞz�����ȭT>Aq 0�,K��y�o�R��me���^ZRjiI�����L�tʑ��������S��,��.տ��+L6�گ���o�&�1`���g:�Q��Y�F�b���$�t   �Qp  @�����[c�01X�;�-�{{{��HLs�U���ʿ����S�@�����m�������}9��rwvԫT� ��� ��,K��Ye�����WfqqP^��W���ܜb��c�i��?����Pp��y�M�a�;DN/�;	���MG}��zYү�   �@�   Q��H�}I_o:pUX�;���"��E~\\�^�mۺu�����8�T�����c�m�7�r����ߗ[���ڒ{�vog�I� ���2w�(57�����v��vzqQ�KG��*��?����\��g�NG�榲oy��(�aQ���c'qLꓒB�!    8J	  ���!IQ��0X�;�)f����#��icc�i�0.Q*�P*���w��x��r+�vw��j��jU��=y��p �ZU�4x �,%�����UzaaXX?*���攜�Sjv����j5���_����Rss�ܾ-���+������?��AQ?����1v5�����3   0��;   ��O4���#�� W�żcQ_��E|����4���%
�q����q��^\|��@����rXzw��O���]�k5�w3���,��'>N��S\q��jgg�ZOF.����%��xCs����aQ����Ob�&L 飦C    &Qp   ���W$�M��y�R���YVd'�2�O��<mnn�P(hiiI�d�t$��,kP�������G>իՆ�w��@n�"�RL�?8�W��S�K������Ai}zz0Y}zZ�����rY��Y%gg�ω����
�p8�=����w�S����~�q`���0 �ܓss�#���a����?6   0��;    mK�I7xZ��(C�b1�Q��%�J��r�U�Q�p+)%�_�j��Z]]��ܜ����w�D�{�[�ܣ��W��_��wp�~�.��c
�@4%����%�SSJ����J����GL�N�����z��~���]�����q�U������+R�0�'w�)�Qp��H���   �i�  ����I�L�F�v���r������\d���k4�,�MG��}_���j4�u�2���H�Q�r���?��a8(�?�_���j��l*��"$���s9%���8,�/SSJ���"�Q�=Y.+��������U��� �|^�瞓��r��w�o�A�=B�z]�癎aL"���͚�12:����U�I��C    �Qp   lI?���c`�ٶM��Pj~^��6���>w\	�q������i���˲,ӑ���]����I�fspi��5�[-y������u��~���u���G̲/�,��׉b����ǉbQ���aQ=Y.�J�L�ǘj����ّg�l[x�;(�K���5��_k:n�[���`'s�P�㘎\�=I?n:   0
(�   �~N�#�]�� Oömͳ�)������r/�h:&D��V�j��Z\\T�P0	�8V*��ܜRss����qN�O���}�VK~�#���]�ݮ|&^b�X�⹜⹜���٬���`��ai=Q*)yXZO�J����|��q]W;;;�m�h��;ߩ���=�FAgy�t� wo�t��~��$۶����U�1I-�!   �Q@�   8H����5xl�|,��^w�tL �u����B����%%�Iӑ H�2�3iaቿƃ��~�5�}���q�s\��v���o6�?�۽�.��)�H(Q,�J&ee�ǥ�lV�BA�BaXZ��r���y%�yY٬���9��b��	x�0U�մ��� L�Qᥗd%
�}�Q��nn*�<�x�	�����1��L�d\�?����C    ���;   p��I���?o6��X�;���bo/���p���VWW5??���i�q \�D�(�W�������W�ݖ�`�q�8
\W���w����}_�mKa(��|�VKaʷm��?�\�S��)��z�|�Q��Gz��J��d�3Y���D� Y��nK�%��g���s9�D9=~XN?�/�HJ�鴬TjP@O$�(N}O J:��vvv���LG��i�^xA�7�0Ũ�����T�LG���I�O��Ϥb�&��5�   @�  �����/Jbl ��z�2_�u+�0�|���Ύ������LG0B���ҍ�0��xI�������Q�~xG8(�? �<��D�=���g��R�?��dΝ:|4%]:<AR,W<��pF O��}U*U�U�Q�Tx�;#_p�${y��{DD�=/�c{�����6   %�  ���I�%�æ� O�E�c��Y�,Ka��GQ�f���8����555���%r`N̲*֟]��	�P�ZM�JE�s��K/��0:++�#���ߵ,��`:���X�\ �c�C    ��2    Q���G`��w,fYJ�Κ�a�{p�p�8�<�FC������W���   <�N����U���t�]��o{�bKܣ!�#���M�����!�ܯI��L�    FG�   ��ݗ���<	�NKFx��0ԏ��?n^�T*Z]]�  0�����߿���u�z=�q.��d�}�Y�1�s����x�y�ݭM����L�t���n3�c˖�I�!   �QD�   8ߏKZ7�,
�����MG0ʉ���0���iccC����<�t  �	�P�jU���j4��\ZᥗLG0/���0�׬�������=`��O��   �"
�   ��z�~�t�(���^\4�(w�tD\����ʊ���Dx�"  }G�[vww��uK᫾�t�����4�,��u��#�
�S�����   ����   <گH�C�!��`Q�T�'�G}��!U*����u<  9��w�q]�t���g��$ɡ�>�܈Op��~�31�~H�c:   0�(�   �����st"���iQ����옎 �����Mmll�qX�  f�����=���L�NX�RI��%�1��nl���k��`��8�1�G�~�t   `�Qp   ����[�C �ԪӢ��ۣ��d۶VWW���%��L�  ���ժ���upp�0MG�R���*��s��&���E��n2��=��;�L �L�    Fw   �b>*��0��z��%r9�1�q��$�Q�fS+++���S�Y
  �~�v[+++��ݕ����\����f:�q���abE��7�'�?�a3�*鋦C    ���;   p1�%����E��}��k:�HIEx���8�M�1�sA���-//�^�3i  \�n����umnnN����[�j:�H�nn���k�5��tcb�R���c�۶MG .�%��C    。;   pq?.���E��wZjq�t���]������������;Q  �+�y����"�#s���T�t�(�O����M��K���##Cu�]�1����%�   �
�   ��9�~�t�"�Rܸ��o�݋��?Ƌ�8Z__��Ɔz���8  `LA���}������b��ܳϚ�a�s��*��q��K�Y�Q�c �.��   �
�   �����k:�8�OKQp7�4۶��������}�q  ���P�jUo���*�JdK���7�8w�����?ۨ�x�b�|T�!:    . a:    0��O�Kb�o��v�m:�Ha�;w��0U���h4T.�577�x<n:  Q�fS���r]�t��/��}�!���Ja(�b�������LG0*��8Đ��ߗ�/M�    �	�  ��{E�?5x�N�D|�;�]�I�{{{���
  �f۶VVV���E��P�LG0����5�c�D�=nj~�t���w�W��   �
�   �����aha�OK��*��n��19� �����|�MPt  �l����666���L�)��%ųY�1���옎�k���Lp?�c`?���    �@�   x2uI�t�<�v�t���,�fgM�0����j��\����������u�ah:  �A�nW��ؐ�8�㌤X,��3Ϙ�a\oo�t\1��T?�f
8ށѶ#�S�C    ㈂;   ��~V�M� �B��a��E��br!&��y�����ꪚͦ�8  �������-���ɶm�qF^��]������I�E��4Q,�bw�S�}��	I��   <
�   ��%����A�����T�'��L.���z��  �`������Z^^椶K��.�"^��DQ�3M�ϛ�0rx��EI��t   `\%L    ��J�MI68�Ž�E}���wD@����Ɔ�٬���T(LG  O�u]��h(C�q�N��{��Гȉ���Q?y�,È�%}�Cr    <
�   �����o�T28����R�r�wDI����榲٬�����MG  �ຮ*����&����wɭVMG��E���4����m������/�   �3�t    `lK�	�!��X�{X���^@4Mt_[[��E  ƀ뺺��VVV��~Ţ�h����
��t\��O������^#�@��4   w�  ���^68���E}8�% D��D���5�M�q  �(�_��3Ϙ�`T���o��o������Pp��[��   <
�   ��$}��5`\�ݦ� +����¾m�g�������E� �A���en�2��~�a:���n������#��<`�|QҧM�    &w   ���;I�a: IA�q�1FNfq�t��������j�L�  r�~///Sl�f��Y����u�pE���6��w��1B|I�'�6   ���   \��T3�آ�,��o��2 �n��{��iyyY�jUA�F,  \�N����MvS�Aɹ9��c����{�������1R|�W��38�iI_0   ��  ���'��H�ϒ��w'�e �<��jwwW�����ߧ� �k��Z[[���:�SnX���\&�O��ܣ~��Yl�f��I�0   �$	�   �	��J�vI�3����,-��`��2 �8�~_�JE�ZMSSS���U"��3  �D�j6�:88`��A�%��&F����8'Ma���$~�    W�:   �ꅒ�[�I�΂c��aܣ] .��}U�U�j5�J%���)�J�� �X�@�z]�jU�癎yɩ)Yɤ��Y�k:�H���F���Y���$���   ����   \�/J�eI�a:��E���MG0ʉx ��0�h4�h4T(4??�L&c:  #��	b��#��R33�~/@�}rD��c�cga�F�+��L�    &w   ��|L�7Ib?pA��a�\N�bQ�V�t#���|�V<�7;�v[�v[�BA333���  I�뺪V�j4
��t�����
���t"�^��F�#�%}�t   `Qp   �OU�'$�c�AM�ϖ^Z���xooO��7[GE�t:����J%Y�e:  7ζmU�Uʅc �h�^�t\7���c�s��xǾ`غ�O�   L*V�   ���O$}�tDE��E}�Y/� ��z=moo��7����<�3	 �k����VVV����{�1��;��&���c:�Q��y�8��!�a�_��1   �TLp   ��wKzYR�tD�|gKG����w�U�}_�jU�ZM�bQ333�f�� �-�    IDAT�,�~_�ZM�ZM��K�"��$t]�p�~�vԏe��c_0���;�C    ���;   p�ޔ�S�~�tD�|gK-.��`Tԧ��%C5�M5�Me2��̨T*)��� �sG�jU�fSa���'�x��	����3��tďe���D`HC��   L:
�   �����o���� ��Ζ��Գ����T*J/..KK��Y���x�DpG�������fff455�x<n:  ��Z��j��:���8��d�t�b�e:.!�<9;;������UowW�Ύ����������p�)I�M�    &w   �fx��Wҿ���*n�|gK/.J���	�~���믫���=�,�.�^(���y�vww����b��r��|>o:  g���j4��j�x=Q�5�(+�6=O��=�vv�;,���J�Zd߯?J�O�?�`�%���   @Pp   n��$���΁�`��lV&��Ԕ�z�t�������u����z,��+�������J-,({�2�<�x6k -0>�0T��T��T:�V�\V�\��4Q ��m[�z]�VK!�҉8��F%J%�")�}y��Ⱦ�'woO�֖��-�*)LG+��Ʊ/�0O��H�   p(�   7�I���9�A0�<ϓ�J�R�������K�۶���ꜱ-|�T:������2��J--Q~�������J��b������*
 �aG�����܈O����OpONO��0��nW��}����"{��{p@���X���sJ<�����/�   Dw   �fU%�-I?o:���m
�g�,-����cL�ٔ�l���=�(�e���A�}~~8	>Y.K���Āy��^��^�+��hzzZ�R��� �k�8�j���ͦ����o4LG0*}��cͫՆ؏�ݽ=9{{�7���EBja���g�P�n�tDǺ�5   �
�   �����o�����`��mM3��!��E�"��l��lJ_��C�Y���33J���������J��LZDd8����m���\.�\.sr ����?�����Lǁ��=���=���#-�}y��p��Ⱦ�����|�11�2KK�#�$۶9Y7%�`g֎�    @�Pp   ��.�3͘���n�MGI)�GB��K�W^y��D.�ԉ�{rnN��E%�畞�S,�4��>�����@��r*��*�Lu \Z��t:���j�Z
��t$���(Op�,e�y�t
�����JePZ��=���S�Z�(	����#�c^�A�R��   Dw   ���%���>e:&�}gc��x�w:꯯�����������`���|j~~0~fF1�p��t:�t:�,K�BA�rY�|�t, ���<O�fS�ZM�癎����H>�!��$+�6�������^�ȫT�;*���˫T��>�R�Bw&۶MG@4�%���   @Qp   ��1I�"�ݦ�`ru:�{���b���)u�+��j�j5�7z8�+5;;(�/.*Y.+Q.+����Rssx�� �l6�l6�N�U,U.��d �� �n�U��)��!�3^+GI��MG���ɫׇ;`�G���rww���D�ܺe:�H�wn�J�1   �"
�   �9}IU����&Lp?[,�TrzZ����(�&����W^y��x&sj�{jaA�9�������H<Z��S��S�RQ>���Ԕ�Ţ,�2 `��8��jj�Z�}�t���W�b:�Q��^2�B|ۖ{p0(�N^w+��e_~�k:"J/,��0�8��9I��p    �(�    f}Aҧ%}�� �LLp?_zi��{�����Ɔ�g>��畜�Ujn��r�qrvVɩ�N�f۶l�V<��ԔJ���٬�X �k�y�����\�5�.�~�u�)���{�ՒW��*��'J�L`�y�dr��w\3[�w�   Dw   ���I�O$�`:&ӬΗ^\<s�7 I}�V߶�-�[ɤR���%��Y���'��Kp����}U�UU�U%�I�J%��e�R)��  W��}��m5�|���ښ�j�tc��R70�:�v�V���ZM^�2���pB
�Pj~^��L�I��5���5�!   �(c�   0ϑ��$��$V�p�X�;_fi�t����������9��e)Y.'���ӳ�J��)53�x>é1�<������N�U,U.��L&MG \R�J�a���1T���MG0*��sO�5B��֫U��U�*y���JE�Z���Vi�]����p�� ��   Dw   `4���~C҇M�da��|)�q�� �[�>rbf<�VrvVə�gf�����%5;++���Ԙ$�^O�^O�JE�\N�bQSSS��㦣 ���:����Z��� 0	�,)�?�����Zm8e�;|��V*���f�f��H/.��0��k�J�I�]   F�   �/�/J����,���)h0����߿/��}��yN"�S�잚�Urzz8>ux���x�N��N����=��y�J%�EY�e: @��[����|�7���/�W���aTrvV���a���$�����H�Ǳ��1���'%��!    Pp   FIM�G%��� �,��/=?/Y�D�#�����ȹw���$�E%�����L���L���U�\���0�n��n���U(T,���)��
�P�nW�VK�fS�~�t$L���|�t�6�LG ����1/\��%��!    Pp   F˯J�/$}�� �Lp?_,�PjvV����(�S�Z�Z�nl��+�TrzZ�rY�rY�%���}��i���X���$���h4�h4dY�r����Qj�Mj����o�a:�+�a���8�+�K�.I��     (�   ��$���Y�A0�Ǒ�yJ2��L��%
�����Soo�������4��������̌�l���&A0��~Tv/�*�������
�P�NG�v[�FC��(Cm��n:�+`%�J�̘�1�Z����,?-�ߛ   �w   `��H���~�tL�v����i�1FRjiI��M� FB����uy��#���畘�VzffP����ߧ��(��MM)��t�쾳��l6�b��R��D�C� �8A����l��nSjǍ;��?Pgu�t W ����l���$2���H��!    �ƪ   0�~IҷJ�K��`�Qp?[}�׷m�m[ν{�|^"�ޓ����RGS���?ڎJ#�NG{{{��r*
*
J�R�����}xrP��V�#!��z]���M� pE8fq>~��
���]gL    #��;   0����W$�L�Sa���X\�a~k��᧦���^'J%%gf���R�\�oX��m[�mkwwW�TjXv��rL�9�^O�v[�m���(Cӑua��_�E�m�t W$��h:��j�ۦ#`r���?0   ��(�   �k[�'$��� o,��/�b1`�E��V*����SS�&�'��rY�bQ�RI�x���G�뺪V��V��,K�\N�bQ�BA��L� ��v�n��j��y��H�){��_��/���
�8)�\��Y��q�!    ���&   `�}ZҷH�z�A0���~�����DBA�o:
��\W�����&
�A�XT�\L�/����RrjJ�bq0)~jJ�T��O� �n��n��ŔN�U(T,��dL��'�����7۶����H��0�Z�7��M����jU{����x �X����8օ+H�I�A    ���;   0��[�˒�L�xb��|1�Rjq񱓣��~���'�Yɤ������J�ˊ�r�ۉ|^��'�e�b�kN?��0��8rG�JE�TJ�|~x�,�tD 8�єv۶e۶�1	z����NG^��~���m˫���j���ZM�fSa����dn�6adq�W�$�k�!    ���;   0�6$����1�m�-s�6w ��SP�˫��\+�<5�=Q*��OM)Q((^,*q�b1�\���u]�j��t���{.�� ƹ��N�3,�3�O-�Z�[����z]���뇷�VKn�.�ٔ��N`%r9%��uq�u�)�I���    ��;   0����Lҟ7�c�E�G�ܺe:�1x��jU^�z���� _,*^(���;yl�'����~pp�x<�\.7,��R)�D@����m�V��7	#�h��QI��j&��w��fS^�%1e�SJs�⑘���h�c�m:   �G��   ���Z�˒߄Ka������u9Y��^�s�dR�|^��i%�e�s9������\���|^�\N�ryl�����V�5�=�L&�e�|>�x<n8!�I��	�=�eG�o���u����m+8���uy���Ng���s�q���8օ������    ��;   0>6$}\�ϛ����Gc��(	<OA�~�2��L��'
���BA�|~X������'���t��T��U?��S�����p�{2�4��8�@�nW�m�����*Cӱp�~PBo����v[^�9��~j�z�%�{�S� �,&�?Ǻ��V$}�t    C�   /����J��A0>�j�h�[��XL��`���V�W�]�s�������D>\�?|<Y.�ͼ���u]5�A�DbXv�f�J��7��h�}_�nw8��qӑpI���n���~4U��t��>5Y���5<��E���(��	���C�m:   ����   ������fM�x���hV&�����j�t �Q�Ò�X�p
�� _(
�'�]��Aq>����>]�~_�fS�fS�q��h�{&�y��`<��}u:�a��B�hgX>?����O�ԏ������N�tt I�6�h���)I��t    G�   ?;����_3��qy��d2i:���ܹC� ."�o6�?,�_J,�D.'�����﹜'�;�(��\N����*�g���%��Ȳ�������Q�ە�8�t:�<�t��z��ݮ�nWA��~�#����;������`�z�;��h�z��0L� 01b����#�	�$}�t    �C�   O�.�?���M�xh�ۚ��6cd�oݒ��e�1 `���`b�e�Ɵ`%�2�uT�?Q�?*�ݟ)�T��V~vV��i��eşr�<������E��R{@q��ǑT8?����*���Π�~Tj� )��,�'C�O���J���5   �1�;c   `|}��HZ2�������7 ����W��%Y���r��r��ޓ�����lV�lV�Bax;��*^,*����f�����YY�����$�	A �q��;������X�+�r�U��
轞Bו�8��]Wa�7(��z���=x��s�'&�+M�T �+���#ٶ�	p���A�M�    py��    �*�{%��b��`ıu�x �H�I�۪�n�KJiP|?y�+���EY��p�|�PP���BA�\N�a9>Y*�J���dK&���Ǖ(������9Yf?����p��ف��ͻ������t�z
<O�m�.�;��^�tY�u�����Τt �dn�2a��Z-�0>�$��L�    �d(�   ��%��������ߣe��5 `�/�{x9r4�=���y�S�yO<Y�q���V*%+�>��RJ�J���LF�����K�e����s���N+Q*]K~DK��New]W�^O�^奔n�y����*����=oP&?��^����bzx�sN~�ѵ��*d2, ��̝;�#�4�8��I�&i·   &w   `�}����DC�b���Ţ����k*& ��p����,�'58�j�D�ÂŔ(%I�BA��N�����$��%)���JN���5���<*�[�p��L*��n�%&�'������.�;�~o\��u8��v���;8�#�}��=|^��ɒ~��0��:ͦz��^�/Ƕ�t:
�pX|�@���P����NG
�S���W�8�� �f��#q��)I��   ��Qp   �_]ҷK��n�c�1����ܽ+��WM�  ���J��q��d�=�1}Q��)��5��*���aq�AGS���fK�=�X����ʑ8�#p��B�9N������G?�p��e�N�8�:a"�`�wx韸/�U  �E1���8ƅ�I?i:   ��C�   ��F�?����`41���2w�E� pI������cY|Q��E\:]^?Yh  7#9==��g���ǨK��Ĺ�   �أ�   L��J�s���t��/{��� �	�?�<8���q���?q�NG%��$���  0+s���#�!x��!i�t    O�5   `rx�>"��҆�`�Pp�w �$����U~?�X�b7��+������\4  pi
��1.<�oJ�g�C    ��  ���'��;I?a:Fӭ/s���I!; �xT�]:.��u<�=��ǘl��׏.G���S�y% ��b���q��ؒ���C    �:�y    ���I�zI�t��/��*5=-�Z5 �3�����w�k���_�?���m��� �l�;wLGyLp�I�)�n:   ��C�   �<���HzYҔ�,,�]L��]
� ���x���U~?Y���ٻ���������Ԫ�[j��v����$�sI�s2	K��b���f��X*�!Da�:��0a��@0vLX0v �f�m����j9���T�%��ڪ�[���zի��VOKXu���ƛ[��ք��o�sk,�7�ڙ�  $&�oC��wH��u    �E�   �M�K�F�_ZAgXZZR�\V4ʟ��2p��Z���  �\�h]��>�)��W��=�M�o|4,k���:�^gJ�jx�U��^�݋�:  ع��b{�U�
�X�{�n�   ��h6    ����.��t� ��lV����1:� `c�&ϭ���^	�\��p����  @'�3��y�)��QA�s$-[   �|�  ��v��GJ�Y�� �L���&�]d ��A�  ��ąZG�x�|^a��Wѧ�X�w�C    h�N�,   ��[��<I%� �Ǆ��\t��2     h/&�o.��XG@����Y�    Z���   @�����X��=
�s������1     @�I<h��QpǊ㒞-.   �4
�   @x��Sm��8	�5ɋ.��      ��7��H
%�T�Q�     Z��;   ����J:iv8	�5�    @;�����[��xo��[%}�:   �֣�   �%�\\��oqpk(�    �vJ\x��u�������]I��!    �w   ���.�6��A�}k(�    �6J:d�+Pp�kK��-i�:   ����   ��k$�c��I��I\x��h�:     �Ƀ�#t�7��)I�Z�    �>�  ��S��,I9� h/Nn��D?�|�     �O0�}k�з>%��    ڋ�;   П�Yթ7�#�ܺ��/��      �ܷ��}鈤�Y�    �~�  ��u���Y�@�Pp�:&�    �vpA�ā�1���S��I���    h��u     �^(�;�~�8� �ϫ\.+�O�͜�ԧj�c�#Zz��Q��U8rDa�h     t�H2����8tHɃ5p�%r��u�������FIwZ�    `�V   ��U����I�LZ��rڻw�u���S���ОG<bպ��\���������W�P0J     :MtpP��ϯ��/�H�C�4p�E���/�u��㽧��_�4m   �
�    �"�M�^k���d(��RllL��1�<�a��S|    ��D��?p�"{|�~�"{���y�ah�qJա,�:    ;�   H�i8�%�q�1�jL�j����œ'����Zz�������C*�rFI    �v���S��A:�ġC�B��C�[G��L�:�#�t���Z   `��;    �:繒�#i�q�'�/�����k��_���˩x��
G�h��-�<.<���D2     ڮ6�=>>���.R����m    IDAT!%�Ǖ��Bɤu���І���>a   �=
�    j��rI�gA�p2�sD��4p���R�5,�岖��Nz?zTţGU8vL�G����`�    �n�@��1%�?�~�8��(y�r��uDl��}��n�   �3Pp   ��vI�I��:Z�����E�J:��Cڻf�/�T���N{�|P�ǎ�xℊ'O�3�    ��\$��y�)>>^-���WK���J<� ����`hC�[��lIe�     :w    k]'�1�~�:�������b���+>>���=lպ��{� ��w    @�	�Q���;�Ğ<tH�/��8a��3���%�L���    ��   ��,�i��� �.���u��{����ܺ���'%��    ��bgJ�T����b���9gmD����*���!    t
�    ��CI/��!I���!����F�9�}��	���ѣ*;��[��)��    ����٣���W���_��Ptd�::�i���%�z�    :w    ������k���y�v��\,����J<x�:_��t�t}�{y~^���j���	-?n�    �-�XL��1��ǫ����j�}|\�.P00`]�ϴz�iI�K*Z   �y(�   8�WIz��߰��`���E"N~����K���|�v№|P��e��    �v�)~�@��~�@���r���/9g=�ϴzN(�Œ~b   @g��   �\BIWJ����Y�L�B3�Xl�����{��qO�<3���	���%�m�    �,�w��㊍�W'��LaO��+z�yrA`}��{ϙ��q�    :w    �yPҳ%}ZR�8viiiI�JE�H�:
z�s���)66&��/��ڗ�*��Uo�����'N�)��<)��Ap    �/k'��FGSb|\�/T�LZG(����Iz�u    ���;   ���Sқ$��:v�{�\.�={�XGA�s�h}��z|�������Z>q�|��Iy
�    �����J�=>:����
	��9�>�BO8&����A    t��$/�Y`�9�3  ��0-��I�]�إL&C��E"�	��^z�z
�    P�^��6�=1>.�[Gv�vEBt����Kz�:  �l�9�=u6�����D�I ����y  �^ҳ%}K��mSt.�^�i>U��S��)O�T��)�N��>?uJ�S�Tf�   �V|�>���W���طO���S���߿_��1�1���ϲz��%}�:  �|�{���uΕ��1�$ L��  ��1/�Y������'�\(v�y��w��~���ƗJ*��k��q��檏W�����U:uJ�B���   � �~qwtT��������⣣�_p�"�1s9���>#�u�!  @נ������  �  �v����$��:v&��ZG :���W|||�m*���Ǐ�8?�����Ǐ��R�/�8��'�0lcj    �":4T/���Ɣ_�<���ׁM-,,XG������z�P  ������ �{   l߻$=Aҕ�A�}��.24��K/�F3}���ܜ��N�tꔊ�N�x��J�OW��̗ͩJ   ��ۻW��1���Sl�߷O�����\$b�	\���-Iz����A  @W���9�})*i�: sE�   �+]%�%���A�=����b�8���n�K%��Y���|�D}|�$��ɓ�L�   ̹HDё�������QEW����W�HXG���ڤ�oY�   ]�N+��sŨ$ƈ��  v"/�
I_�4b�۰��h�+.��c��4p�nW��T<~\��y���U^�_>v�Z�?uJ�B���  �����|tT���jY}lL��e�����s�Q4`XC�z��[�C  ��D�@&*��;}�{��  �Sߓ�2I����.A��L��!\z�α�/������U^� �T������   :A��_��k(��
�ׁ��gY]�I��  �k�e�@���s�   ��W�/�j� �N
���b���+>>��6�X��S�)�O�������*/.��r_:}�i�   �
��aE��O^��<n\߷O.��
�E���uNI�\Ҳu  е�}�9G��$~  �ݻF�#%=�:6G��m.W������sn�K%��Y���U����W�'�ðM�  �/�CC����QE��_)�Gk����S�LZG`la�S�]�"���~b  t/�����[@_��/D%�[`�	�  �	J��.�ے�g�&�٬���!���X�:�rlL��Η�*g2�"|�˩4?��J	�V�/�<I   g�����퓋D���Lp�*���)�  ��A0ｷ���B�{�R���Z   =�I/��7���Ypa*��jdd�:
�.�ѭ��P充3S�W
��充�D�LFa�Զ�   ؽH"Q���g�b{�*:6��޽��ۧ�=g���8���(�w�;$��:  �~��c� �;��!������  ���)I��������)�h*[*�K�/�T�fם
_Yy\���>^X���
  ���}FG:�xp���A� ���ҒJ|I��'�ْ�  ���!�6}�h��� �oι�3  ���&I���	t���E:t�:�>�je�m��+�|u�ܜʵ��\}yinN��E�0l�{   �Dѡ!EGG����QE���<�����\|@�[XX����-J�\�� @S�e �A&����	�  ��^$�$=�86���t��2|r_̩M���r�"|y~^�l���\N�S�T)��   v.���NR_)�G��_��)>:Z/���V z�au�P�K$��u  �;�0|(� y��Rl�D�Zg   =�(�钾!�|�,Xӯ ��Zl+*��J*/.��ɨ�ɨ�r_�d�������E
�  `עCC����o������E��>_YU�LZG S����pno���  �������u ��sG��\r���QR�:��s�寻��zի��  ���SUK�wJJg��l�: ��*28(]x��Y;!>l�_��S%�����r*-,H\= ���8]=:4T��VdpPѡ�U֣{��E"ֱ��Pp�h��4m  ��뮻����lN�֦� �5�l6{$z�WV�������u" ����s�3�  �U�*�zIa�1� vf;�%ɗJ�I���p�_��S%�[��<7�r>��w   ֳ��RllL���Ue�h�r�Y�����d�#`}�I�B� @�9�|:����_���ĿNOO������s��;Ї�s?��   zޭ�-�*� 8��� �.����ƶ�O���J6����٬ʙ̙����a>_-�g�
�y�\� �u�������aE������ޏ�PV����� �rI|�  Z�����HRT��s?���J��� �v�Zҿ��k�AP��A �\A"� �P���F���+S����Y�++��Tjѻ `g6-����^[��/� :�au�Pҋ%��u  ���}��io��n��	��  ڤ$�i��t�8��A �E;�_C9 �
�� ��gX���>j  �X `�6��Vp�w�?�a�]�  �oU�ҵ_�4`���qr Ш���|�z_(����J>��PPX(���T]�˩R((\Z�$ (:8�``@���"��)20�������Y���\,f�  = ��XG��K��  ���� �����Rp�t�a v|,��:  �+ߐt���I�[��r��*��"��u @��M9��W*��{>_-��J����*���2|��r>��Ғ�ʶ�|^�� ���j�|`@.�P$����P�L�.���Ճd��6+� �	�#�껒�o  �H$rO�R��2�w���=R�:�>&�Y" m眻rr�g�s  ���vI�X��w7�|����k ��
��d�����Ҽ_^�����׶����+����"ey ������x�\$�
�zY=H&I$��j)=����I&:�>�~G  4��^/zы��u�~wRң$��:  �/�t�~I[� �>��SSS�3�%�^I�m	��=Wo   V^%�%=�:H?[\\�� �9A2� �lʱ|���X�����j9�P�J�z��R,V'�
���R��_�X]���P��T��@�H�^(b�j�<���bՂy2)�U�I+� ���W{��W9�� ��r��v{EI��v  `�Qp��s�;�Ǎ�{D��+ι{�3  ��Jz��oJ�y�,}kqq�:  ��b��b������%)U�����j1�\VX,*\^�.[ZR�
W�=��Ru��6a�$_((�T��?�o�,��,I*�r-y����䜂DB.��F$�s��E"�y4Z/��h��.��}�x����F��@��� @��+s^իp~�:  �Oι{���Y� �V�Nk�����s�& a~�:  �k�&�+�F���%N `�V�mU�~=�����\�/��Pa>/I���aX�4�+U
��~��佼���l/��~e�f�0�>,���3�K%I���W
�>���b1�$�)�K�Ҹ�j9���ʿ�ιU�>G�����A��A+�DV&���\<.9��ʱ�����Ū�^  �>�2w���b  �/��7�3 h�z��^p�F�_�pY\���a��  @߻W�%}DR`���p� ��S+G�sl��T�����p�eE���:ˤ�R����S*�R,n{�F.Qd�%�`�~��DB���.�P��^�֋��}k�r  ���d�#���$]o  ��H$�5:�@����x���t:���ڞ����R���  ��M�n��o���+���      ���������Y��G?��(I���   �����{�u mq<�J�_{�jB�s�i�@���u   ���t�u�~�,      t*>�21/�2Qn  �{O��_m|����8�@o���  �I��+%}�:H?Y\\��       ���{ە$=O�?[  ���
��U�ֵ�/�7 +��/Zg   X#/�ɒ��/(�     �S-,,XG�'^�u�*�  ��A@��ι/6>_Up��rߐD��}����=�!   ��SIOW����     �N�gWmuXҭ�!   ��d2ߑt�:����ݸ`U�}zz�,鮶F`������:  ��.�E����2�      �T|v�6wH��  ������s h�/^}�ե���-��_h_ �s�� �N�aIo������J���      m����[�3%y�    �@��}g���Up�D"�2 z\�R��:  ����X��u�l�:      ���^�\�:F�{@ғ%��   �K�tZ��Y�ֳ
��J��v`�7�p���C   lы%}�:D/[XX��       ���d��u�^� �2IY  ��J��>� Z�9w���_�Ok��Up_qG�� 0���u  �m(Jz���X�U�L�:      ����u�^V��<I�X  ؆OX �2��knTp�У�s�| �ns\�S$qV�8Y     �N�gV-�%�J�'��   lGtހU�T���^����f�N�G�^t:��~�:  ��#�
U'���8Y     �N�gV-�vI�X�   خ�.���%������d�K�X��>==]����F`����u  ����?Pu��daa�:      �
���[I�[�   ؉+���"�S�9 4ݧ������V�[p�$��_�. ι�a�  `��-�u�^B�      ��Ϭ��^I�I  ]�{O��=vZ7,�g2�;$�W#�;Ng2��[�   h�)Im�W0      ���{S������A   vcϞ=��t�:��Y�`�+3lXp���.x�?ޚL ��{�����u  �&�#�k�Az����u      `
�M���TIZ  ح����$���������VnXp��H$���`��g  �c��.�t�u�n��B      t�:�eU��m  �Y��t���qΟ�s�?/�XS� ������/[�   h�9IO��ەL&#�u      ���6�J��   ͔����S� v�X6��¹68g�}zz�,�}M�����uzz:��  �ߗt��/[�s�P�L�:      P��U�v���u  �f[����:��q��������Yp_9�{$1��^�s��S  ���%�L_�ۡ���      �$)�˩T*Y��fwH��:  @�8��-�b���y���f�lZp����Oҗ���ϥR��X�   h�H��ѭ(�     �S,..ZG�f�(�b  �a���?u�}�:����)�J��f�mZp��S�t!~~ @9,�ϬCt#
�      �|V�c�I�}I�    ��!�8�Km�ӺՂ��%��U" �d2�  �F���:D��!      :�U��IO�t�:  @;�r��Iz�:�m;�G���
�K�޹�H ��9w���t�:  @��D�g�CtN     �S,..ZG�6�Nn��u  �vY����u �㽿u����-�%)���$��@�X��6�   ʒ�!�[�A��ѣG577�r�l      }*C�������M
�~z�u   ��,��P�D"����n;G���y�s�y���ݜs�MNN��:  ���%}U��Y�&�x\������p���e���S$��     �W*�4??���y���i~~^�\�e
��:n7)Kz���X  ��N�o��R� ����T�[�8��#G"���aH��|�9��   ƎIz��%���t�b���Ǐ����n�Q~hhHCCC���ݻW�m�;�      �@�RI�\nUI=��Ջ��|^�lV���:u�*��u�^�%M�r;  �sA�=×h�Þ�_o������N�ӟS�$�s}"�J=�:  @��UIwJ�c���b1kppP���;�_+ɏ��)����     ���zc9}mq=��)��knn�:.�7H�c�   � �NBғ�s 8�ϥR��������aRp:�s���   :�ݒ�%�c���Y�V�T��ܜ���t�ȑM�_;~m1���      �MYo����y����0�����KQn  ����aRp:���Î ���wy�s'�h-��g'''�:  @z���K
����b��FFF422��{�jxxX������p}Y���Ȉ"��ul     �-	�P�lV�L�~[���l~~^�LF�R�:6Z�IO��7   ����J��9 �뫩T�7��ӎ�����O�d_ ����	  ��}P�!Io���*�J:}��N�>��}�񸆆�488X�_�_�5N�߳g����F     ���h�z�V[����癰����LQn  8KoÐ�;Ё�0�ӝ��k����J�����%�.�J=�:  @��Y�X�@����ke�Z9��߸|�޽rn�v    �.P+��������/..�R�X�F��O�c$��  Щ�����o��*_K�R��Ɏ;��.Ia��];�@�y���:  @�F�IWXAw)�*����ӏ��-�S+�ixx���񃃃��S�    ��ڲz6�������z��9�J%���}G$=Q��  6s��W��d�!�s;���9�N������1 4�GS��3�C   t����Jz�u�Q<��𰆇��g����hdd����|dd�>9>�LZ�    ��,//+��)��*��iqqQ�LF�LF�l�~[XX�/+�ֱ���U���    �`vv�����Y�  y��vjj겝��	���a���`7��kIl  ��%=Iҗ%���Y��b��ӧO������/�kttT����&�7ޘ    �F�MU����eLVG+Hz�(�  lY�\��H$�d�`�� ^����L������s���q �s�=���/��  Ѕ.��}G�1  �IDAT5I?k�0A1    �.Ձm)Kz���X  �6�����޿�:�ϼ��}jj���9Ʈ����F"��I�� �H&��  ��QI���$���Y��+�:~���?��}�Ѩ���544�꾱�QQ>����     Z�\.�K�k��ճ�l���:�e^�u��  �#�H����3%����%�ܮ��KM��.I�t�5�^ߌcضT*���  ��%���C�������V��Q�   �&��4�����yy����O%M[�   �f���)���u�9�^399���g��%)����H��f��}?��l  �|S���4h��Y�bQ�bQsss��w+��������    ��YA�\e�b�h���$��   �6<<��L&�I��u���(��4e`sS&�KR:��\���:�-��T*�)�   =�ɪ^��6,�c6+��b�U�4�Q$�~    z�z�R��j�FS�k��9�Iz�u  �^133�D���s ��{����Ǜq���%)�NR�e�<&��y��zjj��9   z�s%�OmV uk�XL�D⬩���c���\S?�   `h�	�[�XT�\^UP_XXP��o@g�KI/�  �kfff>�{�u�OܑJ��Ԭ�E�u I*�˯�F��$i���p��H$r�u  ��I{%ݬ&)@�*�*��������hT�������@��xK&�J&�g=P2�l�   �O�P�ߖ���������jϗ���%��햖�����n�t�u  �^��s�	�Ƭ� =.罿��lzYcff�Z��ۚ}\ gx�_>55u�u  ��jIo� �'���q�b����׶i�&�F��GFF�p�
   t����R��b�x���b�x�T������|>�L&�r�l�V ��g%=Iߜ  h�t:�rI����kS��;�y��ܧ������������c���_J�R�w�y�,   }�m��� �V+����z9�V����������
�   ��4�΋Ţ���b��rz���Xd_XXP��o ��+��(�`  ��y������$��u�G��%�\�W^ye��mz�]�>��0h��~��Kz����}�Y   �Ȼ%��: t�x<�d2�d2���!%���Z)>�Lj``@�dR�DB�DBCCC���J$�u�d��<  ��R����e---iiiI���*���rZ^^���
�B}������
���Ţ�����.--�X,Z�% �Tߖ�XI�    �`vv�%}�{?h��1�A�����w�}���%ivvv�{?۪���9�����[�s   ��@�G$=�: �x<^�_�$�ŔH$���k��'��b1+���  �Wզ�7N;/���k�����޸_�9 ���Q��>o  �����WH��:�c&R�ԟ���-+�OOO��ß��V��O�s�����]眷�  Ї��>&�2�  ��i,��&ȯ7E~``@�H�>y>�ippP�hT�DB�dR�ht�z  ��h,���e
-//�\.+����/--�\.o8=�X,�P(�*� ��}�~K�1�    ��{�fgg?!��M��r&�y���tؒ��5�>��=����u�>p2�<����:  @�K����[ t�Zѽv�v�|�4�Ƣ��}�N���bP�o ��q�I�R�����q*�z�k�d2��e� ��K�͕{   ���9���W��,@�[(���馛Z��MK�433���Z�:@�{F*���u   (!鳪NY ���ɤ"�ȪR�����Ѩ��䪩���d�^�w�ippPAԏU+�מ'�I�	 ��
��*��
���0���Ҫ��|^�{---�T*�P(������B}2zc1�v,  �ਪ�)~�:  @�K��O����9�n�����[�-/�KR:��M�K��Z@zG*���:   �%�)���A  h����7>n�H��6����ݯV� t����k�����Y���N9�h������=^ZZR����  ��iIO���    ����}�����9�n䜻mrr��~�h�_@����5��ÿ*��x=��|#�OY�   �*YI�#�K�~�8  MQ+�r����f��J��488(�ܪ)���%ihhH��D�H$$�>�c �D�·$��yI�O$����eU*I�����ƥ3�Ͻ����Z2_{  v,#�2Qn  �(����L�W%��u��ܛ�d^Վj�wI:|��	��nI{���@����?rjj���A   ���$}Yҿ�  v�6U�9�n~``�R}�|߸>HZ]�_��_�p/UK�ιUy� �?����N��]S�T�pI�ޯ*�׶]�,�X&�M��kiiIҙ/�ݿq}c��{�J�R/� ��������  �����o�$�~K�� 6����T*�/�x���%iff�J���h��]�{�655�q�    8������:  �/�E���������U%�D"�H$R�v�}$���kje�����x�F�S�%����Z����&�o$�������^�X�>�B��0Ϲ�\.o����V��]�����Xk��a֋ݍ�X��1����k���s�(j�r  �6[��4I��  �����<�9w������gMMM��v�`�(����$������snzrr�O�s   `K~N�)L���   �}�2Um�   }�(�Y�n�  �����L;���:�ɜso���|u;_3�|���f�$��~]�[8�n���x�u   lُ$�����   �}�Ţr��9o��  �NI�D�  �k�R�?��W�9�N����_���~ݶܧ���J��\I������w�0|�s�o�)   :ȏ$=N��     �~U��BQ�  �*�9�U��oZg:пT*�g]y啕v��k�ּ��o�� �.i�U������R��X  �����/I:d      @�����  ��I��?#�$�o��'�0��n��/��	�5+o��%�2 ��9�w�]N�  ���P�c%�      �-(�  ���e���Y���{�U�]2,�KR*���s�Y�ʖ9 c%��3&''�n   M�CI�%w      ��Qn  �!�T�n��S%�� �*��799�U��wI��������9 #�{���ħ��   ��~�j��A�       Z�$�E��  �S�����bI�:`�{��T*�Q��wI�����{�z����LMM��:   Z��+J�      @����?h�   -�J�> �5�9�v�޿~jj�f���4J��o�t�u�������&�s   ��~A�%4�      `�(�  �t:�FI������R�ԫ�C�tT��{�fggo��
�,@+9��>99y�u   ���$�)�u       ;V�t��X  @{0���9������9�u���:@#真��|�s�6�,@�׉�����   �⻒� �u       ;R�v  ��399y���V�@�/�ɼ����R�ܥj���/��$��:���f��-   �M��~�:      �m)Kz�(�  ����r���N�,@���K.y���thd-g`#�{7;;�g����4�-����Pn  �{�"��ƭ�       ��v   �{���t�97a�h���r��+:��.up�]���g$MZgv�9����ɛ�s   �cPr      :�v   �233s�s���9�]���́u�sq��T*���:�,�y���)�  `�{%=Q�	�        �U�t�(�  �����[����Ա�``�K�R���r������ξ�{�.IQ�,�U$�"�J��    �XWu��~�        �j���n   �ivv���wK�Yg��✻frr�V� [�5wI���}��y��� ��y�������A   ��(�      �#�t��w[  @g���y�s�%��l� ���T�#�A���
�t���W�T>���l�����SSS_�  ���I�%w      �RIҋ��v   l��Ç��'%�o���iIOM�Rod;� �511���_��]�,�:���?�r;   ��ے#��       @�*Jz�(�  `&&&�Y�T%�n�,�:�T*��r�ԅ�kn��ᥥ��K��:���x���^{�u   t����I?c      �#Iϒ�q�    �N333C���{�u`ŧ���o��� ;ѵwI�޻t:�'ιת����wν5�ɼzzz:�  ��w��%�_�      􁼤+%�a   �m��z�s�?K
��9�ޞ�d���NkO��ggg��޿[��,�;�J�R�  ���_Ւ�í�       =,#驒��:   zG:��\�{%�ZgA�Ytνtrr���Av�'
��ַ��� �����:��s�[�J��n���Y   Г�I���GZ      zТ�'K��:   zϛ���K���_I�5�,�ߓtE*���u�f�K �p���f���{�u��;��=�v   ��iI����       @�9%�E�   -r�M7���G�m��l6��^)�K=4������s�s���;��N;���^�|   �FR��H��A      �pR���m�    ����Wx�ߩ�U��f����������4[O�%ivv�b���$=�:z��+��U7�x��A   �w�n��{�A      �.���'J����   ���������r�=�.�΂���H$��믿�G�AZ�g��w���/s����~�:�V�{?���f���C�0   �[QI�t�u      ��H�$��:   �S��*鰤!�<�Z���?��NkO�k>��0o����Y�]�s_.��/����?   :���IWY      ��wU��~�:   𖷼嗢��m��ߴ΂�� ^611�]� ��wi�7_ҒF�w{�#WY�a�y�lw4ݖh��J
H �!�"	�E�`P	��L��"d0 m�j�����e�ƽHJA�!����B�@����s^?̖�B-��3;�/��O�yv3�d��yO�ս7��v�����I�$5� �\�:D�$I�$Ij k�3�7R�H�$I��Coo��1�>��{T�Bo�y��3ft���WS������t���
��OC_Mݢ�B�]�R��9u�$I��7 פ��$I�$I���j�`g�I�$�}���N�1�c�z�է���j��ŋoJ�2��n�[WW��B����-�υ���啩C$I���t=p-M��N�$I�$I� ����C$I��������cS��n�B�~�\�e�
�RY�j�?�̙sKkk����@1u���c��X,����X�:F�$I�VS;}��K�$I�$I��� J"I�$�U�Vm8���>88�:07�M+��V��;w�hɒ%Oݓ�������M�7�,u��M��Z�^�hѢ�S�H�$I�ap3M�%fI�$I�$i�/�� 1q�$I��O�-[��B�p#p1������BW���SǤ���]����*���S4�	!,,��Ϥ�$I�F�%�π���$I�$IR
X,N"I�$�����c������N��wb{$�pU�\~:uH���>z{{O��|)0+u�Fݟ�<_|�UW=�:D�$Igw�S�H�$I�$I�(ݩC$I��Ѷ|��,[
���E���,��J��R���{���}
��OO���Bx<��e���H�"I�$�����O��$I�$I��� ppG�I�$i,�lZ�n��ٽi]�p�!����9p��)4��7��:;;M�"I�$�������C$I�$I��1�� x8u�$I�4^zzz����v�ow��Ú��/������<� ��{�v��ʲ��\.?�:F�$IJ�j��;&u�$I�$I�4^�6��[�I�$)������y� �pPLݣ4�̲��T*=�:�Q8p����ӆ��.!\��G��B�}xx�'�-z)u�$I�T�����$I�$I�F�������C$I��Ժ���B����G��B��.��/��i4��Coo�G�<� ��"�=S�����b�����J$I�$ՙ"p�Ӭ$I�$I��F�8x%u�$I�TOV�XQܵk��!�K��pӚB�ܚe�ݥR���A���(Y�|�Q�B�1�K�i�{���!�;B��J��R�H�$Iu���8u�$I�$I���B� ���$I��YOOϡy��Ͳ�{1��R�4�7��Y���T*�K38pe�M�6ͦ6�05q�D��}�q�ԩS�7o�P� I�$��� \�:B�$I�$I��.S�H�$I��R�dmmmsB���n�(Bo��1��u�9pC�J�#S�L9;�x�`J��&� ������ϟ�+u�$I�����B�I�$I�$i/�\
�C$I��F�bŊ����Y�o>p�ہCwm߾��J����A��qR�TZ���f�.���{�x(�xo�X|�Q�$I�4�����!�$I�$I�D�F���!�$I�D200Pشi���91�s��S7ձ��6�+ݴ��tuu�B8�p*�}��6�1���;;;��:H�$Ijg@[�I�$I�$�}T��"u�$I�4�uuu}�6�$NJi;�ݴ�MԌ�ׁJ��2y�䓀�B��Y�A���ҫ!���y��zƌO���WSGI�$IM����L���$I�$Ij<o��N"I�$5�����ƍON˲lv���'Sw�����1�'��;w�\S�T�SG5;�u���o����,�N�1|80u�>�
��1�!<U(����x!u�$I��w<��C�$I�$I����M"I�$������j�:;�xb��� �׀gB��<_����dGGǆ�Q�_�H__��CCC�gYvpp��u0)a��B�q}�e��y�>��lKK��lI�%I�$i�<�:D�$I�$IM�e�,`m�I�$I{���?mxx���qY�����!�#���zӺX<�����I�&����x%a�>�@�Riikk�B����4`za�[B |l���:��`ʻ~�v`�mvQ�f��#�7�m1�W��!��b�[����3gnnoo���)I�$ilM� �N"I�$I�����<�:D�$IҾ(lذaz�P�B�c<8(�p0�ݴN�G���M� �-���#�Wc�[��Y�m�1nޱc��J�2�� uG��\�    IEND�B`�PK
     !M[���  �  /   images/a5640015-ff5c-4848-bb8b-6d4b42e5489b.png�PNG

   IHDR   d   ,   ��U   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  eIDATx�՜{��U�����nw�����n[����Db(����!J�Mj�$`$��	j�/�HH��"�JA+[JHw�ew�m�5�;3~?w~w��tvf��-z���������y�o��з�?��m���G�� 7Z0���,�HX2�������0s�k`�����gL��b1�f����㑑����6444�f�qM&��cL�7��Dr��vy�ZKK����Y}}��������'��sm����� �(q�	�@�N�b��z q>PH#�T�����q__������?�u��	��O��&��-�¿袋�q�TKK�1	fX�Rz`�Fzz,%��RB\+�Vs���ga�#i�C�ʈ��}P�C7�ߊ��=��`	>œ&M�z�~��u��z��s�9b�<�=z���L������Dr�x��R+M@ )	s������^�A����n#���֪�I�R}0�c�l�P��r��S����J�0�N��@��9Ӫg̰�E��a�76� b���p�4���O���������_�y�B\'��MҤ��->y�%Ĭ�Vw�V?�;&��9��2��i� �H��wX�=">t��4�'-Huu9�<�S�[�}�;���c�ſ�'�ZXQ�7�+�0��!i���n3W����N���&����jC�����[l�YgYV��0+��  �=�����G�3�/�o}b����s�lD L�D�|�����\&4�<@��Y.:��EHQ�P|S�A�8ٙ�c���o��2��>�Z���A��Д)6 �����>���H��ng�`K�);?"��-h>��
��O}�x���$-h��얦�459-�;�d�|�IϮ��a����Q�+*�E�-���Y}8rV$&#!�'$��r�PeK�Xϛoھ��[--�K��Z�T�='�O��0m���6�	�n�<;�3�i�
�1]2Yh^\��u�0@�͞]HC P�U�E����C�+
��dav�@���6[~�A����6._n��l�SW�����Fנ
 v�{�HpI	�J�̀��(�i��i�P��ò�������NZ��� Ǥ��ɣ� "�el� ].���e������4��T���g͝kS��q�B�u��G��S�G�Q�'?i�n�����oC��oq>C+��3���f������a]��u<��(-҄�{�؈�cQ0"=�Ƣ�Ծ"��"�� i_:�I7Y	���Y2U���r���@�*;팸V�k8o) � 14�A�(��ߨ�5��A��t qy ��,]Ӧ��BCF�8>���9>`�� �����|"�G �`B�	>DH|c��Z���1��@V�X�����6,�&���p�*g�d֪,L���߽��B�O=ՙ(2����Y�;DB��X�@�"�� �;Iya�e�D�:=Q�V��p�d��ciiW����O?�&�U��d�;}_���f�\�L >�4M�%= �)h(c,Ah�� '����Z�ż�je�Ah��� �B
�Ci�7�~��,sW�� ��*�Qڂ��g�~����8�|�����SOS���.���[�mVA��3����Ѐu)EM�.��������޴�!�iO�򓆏ܚ���<�'���=0�Lr+��g���6N=�D�7��_Jj}�U�*W]~�'l���g��Qѝ�h�RI%:r�t���$p�������euO���]�I��Y�0xH�*����KQji�����x�&]3Yf�Gt 5�i�\E�J�mmc��ʕ+[�j�U���$>W��1����K/ھ}��:�O�3=_��de����R7�U*�]I����-3C����P~��m�Bט�V|���u�F��b�sk)6R-�)��B����1Ν��޽{��r�9s�g/�䒃ZhI{o�:�ϋ�9�%u����t{�0LҚ5k�D��/��PEݣ�QNw!i���  ��LBP��@RҞ��Id�Z�Iq"(s�DP�|�r��瞳9k׎�'�@l�Q��o�V4֯�1��ء����~��2�oY���������2���+1(6|�+����}�'�
�g�����Kve<�Ջ��w�H���,%���.S��1�FM���_�+�H;b�2/cb<z~��EΌƂ�� 1��˗��/���XF P�P08�$�k �yk��U42R�J��g�e�m[N�EV�c����D��G>��d_.g��-�K/v�Tň�1��^{�R0�xo�] Yl" �bb
�Q�!�wA����Bo�A�s�Ǜ��@l89ߔgr�#��^V�/sc�̵��{����TN ��wK����S%4�
6�<az��\�U_�u	$f�>P�U4��b�	Y=Ŵd�sD3ʸ�V�@�ԡ7�d�?��")@I46�ayb�i���DdUDK�[�'�HT6����|��n׮]�lٲ�N��e��%i��֦o����U��͒3��o�!q9�r�(��b;vX���j
 0G�Z������R�(*1W=�����7���q*���EN�LJhU��e�y�66��{�Զ?��+� ({ �I��ͽ�Z��<"SdQ���/�}()A'�*�2ǃ��H� ���M�M��%�r yD|��h��I�s�9�7�|�o�k6m�d\pA��p�:_�c�z��R�B�4]�S�|�8܅�ҹe��\~yY������h��ڂl��~��kL-B3H�������>�쫷n�ZN��fϯ-�f�K� �
�*u+��+�D����k��?�p��ɵ�]g�Ѵk���e01��2x�%�F�DZ�(���=�i���g�7n̕��!%Bj�sؕ�b��������y���u_:��Γ@yiݺu��\s��I%��@F��o�����B�'���l/�7EV�|rɞO����$h��K����Ü�~�V����My8t˅����wu]��v��YR.�za��(�j�?,�Q�a��ʝ�ehE�D6Y�A/����-�A��4r6���ݮ۵t9�U+���c����z�Jd龺�-@��B�\�@J�5�_�
S�t��*��x VnB��z%�&�0�����&sqP~ �nݚ;nc��;gv\7#�p����T���Bh�pM�g�� �*2+D�l��j�p����a�#��+��;��i�v>��l���4c��EPhBF;�ۦ�D^5���ٮ�|��E#,r�-��r����m��	M�d�E@Q򨘢R��*"-V2N��cr�����ޯ�P�7s�jg��?|���`r�#�	�K,`�*��lL�������=�a����i0�����������$b�|>1�l��7bss�[��Z���7��d�Ιc�
�iX`˷���`��Q {-��^�����BX��}o�aIi���뭍����(�8�'�����/���g9γ2�l��Y"D�S��̟o�
����5b{�g��Wd���C_sN^��5��hM����|W!�n	SV����:��6�����G��H��l�+^��ɲ*!ПECB�݌!%_-�ۙ��cG^y����uM�԰X�'�\��#��a�V|�|KMk��+D}g�v�l�fS����~�1p�؊h�,��E(����Y�%hL/��#�z��L{٘���e�}J��D5�]k�2M��6[����C���fk^��E:߭듛7k�l����9GF!3c`,ɠ_��@n$��mQ
,j@v[�}�;��zI �n���Ӝ�p@��A	�[��0�ޜ�f�r�k���HؽA���@ �o�n2>�W��xj��/ �d�@��"��x?�4���s�&K]�� h��x�YǾI�s���3v�h��ӵt�Pv���]f)�c'I�\I�p�_槏r(��O�$�ڰKI�7y��aB�]�?, ��[�T �w�{�%�M�e�L�daR��"�=$a�g�#�� �3�\c�@��X!�ہ�Ycc@�+m�sh�hX��<ely>�l�ާ,J�@���E�)YX,�x��������l^����%ָt�h�@�:׃(	A��nE��������$AnłHilp�����'De����x�>c��O���q�z^^��+�~a)Y�I��\�g���ſDCz�!׽A%տME�W��;��"$ڄX�$w���R՚��1���;��(<�G#�9���1�Կj�{�/r�Q ��x�xi�~*�b�#���klx��Ɯ@�������?����z���|9�8����0ή�R��9��V��� d��-�h�'D��x�����{9t��r�1���x�Ȓ'����Ev���,'_@�g���1�����b>8 ��D    IEND�B`�PK
     !M[�wp�&
  &
  /   images/1cdb40d8-22d5-4761-8204-85ee5f97d036.png�PNG

   IHDR  �      ��֗   gAMA  ���a   	pHYs  �  ��+   %tEXtdate:create 2023-04-18T17:15:54+00:00SMK�   %tEXtdate:modify 2023-04-18T17:15:54+00:00"�=  	fIDATx���!�Va���1�l�tW�&l&�f�=�Y��`uF NW܁#8�~��2s��<�N}�KߝB$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)�/8�{����a�$_�~^t�a^;'yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yHYN����qr�݋y>���y��r9�WC�ݫa?+����C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C�r���-��.����`�<�!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)�L��<�i���l�6�8�n������f��5IR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR����? bw.g�����9���<pM���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�H~���p���u��$���y:���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E��8�w�q·H~����-$yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)�#=Ng    IEND�B`�PK
     !M[!��Ů  �  /   images/9ee875d8-7c7b-435c-a3d9-92ac29f03ab9.png�PNG

   IHDR   d   �   ����   gAMA  ���a   	pHYs  �  ��+   %tEXtdate:create 2023-04-18T17:15:54+00:00SMK�   %tEXtdate:modify 2023-04-18T17:15:54+00:00"�=  �IDATx���]N�@@�� !Q���5.ـTg,<;��r��%��z�N:6��0��Ch�1��Ch���ǲ<"�ؕG��U�Ǻ<o�&�3�?"eL��s�?G�G?9�i�1��Ch�1��Ch�1��Ch�1��Ch�1��Ch�1��Ch�1��Ch�1��Ch�1��C�?�-E�w8�%��>.{t��.	ǘ�;�k�2�2������#g�"�*����;�3�KJ��:����o���א.6�*}�v�zju}�.n�&�O�'�aDR���gxA�1��_�ԫr�|�����MK�2���b���:�C/k�u�Z�+���m�����t���.�ʧ��qV�޵�lخ��O;�w�/j�m����ȯ`�!GƮŚ�RC�Y�]Y�|w-��M܎�g{�Y��k5���9rd�}��}���y)����>�4#�/��1��Ch�1��Ch�1��Ch�yQ�K���Oz    IEND�B`�PK
     !M[����� �� /   images/99708c53-ae63-4787-a3c4-6dca09af2b7b.png�PNG

   IHDR     �   �U=�   	pHYs  �  ��+  ��IDATx����s�W���7�|/"0G�I1��Ė�
-�f�gzg읲wm�z���*�]�����\5Uޝ��O蠞n�L1gI�D"@9ދ��}�K�)0h��{�|T(�Ó�s���$           ��            X�            �2�            �.            �p           �e�            ,\            `�            �             X�            �2�            �.            �p           �e�            ,\            `�            �             X�            �2�            �.            �p           �e�            ,\            `�            �             X�            �2�            �.            �p           �e�            ,\            `�            �             X�            �2�            �.            �p           �e�            ,\            `�            �             X�            �2�            �.            �p           �e�            ,\            `�            �             X�            �2�            �.            �p           �e�            ,\            `�            �             X�            �2�            �.            �p           �e�            ,\            `�            �             X�            �2�            �.            �p           �e�            ,\            `�            �             X�            �2�            �.            �p           �e�            ,\            `�            �             X�            �2�            �.            �p           �e�            ,\            `�            �             X�            �2�            �.            �p           �e�            ,\            `�            �             X�            �2�;� �y�,�)�K^�c��+Y��%�J��>������Y���-N�-J�T����U��6=&���H=�V}�H�d}�5�%��Ѽ�֯K����)i�a��k�o��:�����/��B��f����t�a��wH������Ϛ�S���:<k�gH�ĺ�����4�?U_�#��{I����w_=�������{�ǥ�|y�&�?.�?U_����]��S��������Z����6������hm�������>�z?�c�߰���OJ�T��e�=��'�b������^������S��S,�`^/���־zJ]��?���{��������Yϣ�I�d����?��S��%�.<[�jۓ��.��B��y��8ݓ��h_=H��t��1�?)��i�����?ԯ�Z��-�'�}��ǥ}���i���>!ݣy>k<���|{\��_j�>m,�[�}q��ߟ����7���-���}B��K�ԼZ���V��h�b��~�~���������	���������1u}�>�D�g��~}�w ��]� ��������Jv�mjj2��me��Y�Em�������O�P:u||\QUU��U���zg!�#��"�i�ҵ�t���%��y*�Ұ"K����H�yq��������TY���|?O��]�n���B]�6�[-�~P��_Ҋt���|��]��[��u��5ٶmo����k�<]��D�{�W���A�r�G��T����k?��p_=��*��������~i��eK����C�ԣ�!o�W�����+ڰV����%���~��n!�ln6�v�ݻ��ѹzl{�׻�A_=���������}��\�a������E�K���|x��s�|iגu�:�POȯ�R��zj} r�f�����C�􄾪�kO�����+�?��v�,�n�R��hދ��I���I�5���~�� =���/�_�߫�R�_H���B���m����GY�W����z�b�{���?v�����Pދ��`�	������?ݿ��R���u?O�1mz��K����K[�Ã�>��:ż���.=�y}��ګ�8�,jW��ǔ�POe��o��1�z�1�/Iߞ[��c�K���W��O�W���=�����۵T�G��P�)����(���I�������x�bO{��S�Y��b=��<a�<��<����/��3b�2��aOzr�Jҳ��]ۿ�����Kο%�]����_\�ǵ��\��W��������ϒ���G,<���H��z-����.�������Yd����}�A]�������:<:^��賺x�X�]�4"Q�8���f�;ŸOZ/�ٳ�ه�%��{kh��o���lҢr�e��&�o��qqH�L�1j}��vzЯ��ݏ�����D��~Zj\��˗�_=&�� ���}�ĸݟ��o�Ï������ER�?<��=c���ǍO��Emzڸ>v^=�V�_=<�{�&����[c�h}�����(�:c��x�q�7�bΔ����ǟ���V_}�y%�ֵ�ΫG�צ�|��y��z�P���Ճ���_<����~Zx��H�,����������W��m�I}�K&�`K���h�oΣR�ܴ��O|#���Z�gL�.���5h�{���.�ڙeP2�J�h��9����~Reu�}���{�lC��A��#}��&uxx��{�ն��	�0�E�����9K���E��w~mmm�} �T�ǃ�»�6���(����y�B!��S�E��ӹ���w���~���^��]"�B�Z��|��s�·˗D�3!�|U���\iWۋ�>�'��N�~5+�&�mnn��(m��.��k�1#vKK��Ζ�y����?��q�iffF��yU�9�������SSSZNωZ�r�[�U�*��<��w�W����u���WEў��ֵ6��:��e����C�����~����:��im�1s@z�|]�Wy�?�?�܅��+z�}�>�y�׊���K��C}�������O��``��s�"�Jm��V�~��\D����"�����|�[}��S�_��r�Z�x^9�����s�����A�E��=�)ϫ��,�9�B���?��ޯ��K��aٟۏ���%�����>�=~-���Tm�Z�9ʒcu����~a�H��|eM|��&�R��A���߬%Kŭ�������6��ߧ�  <������2����w�}�R�ܐ5vl���¡|S�� 6��eY�1��W�ѡ����@��%���_zy�A�`�AS��:A�va@����W��O_:hn[����'����"��$6'Sl�������i'��̑p�,��ڜr�l���p�������A�,��j��J2|��1#�����nt[WLVw��bj�Vy!��*����?����׆����}��u�Y�����$�����jn`pb4���/��P^8�ۍh����;�-b�AQW��Z���R.x�n��X�>1>!����ʾCf�.^u�7{I���� chnȘ���'�s�۷���w~p�%3[�g���dʦV�K��g��̲�/[ɹ��f[S�%Қ"m�]U��8V�8v�^�l5�ɓS�/?w�ڶq�i���\G*KrA-��R�x��_�tFY�q��n�_����m�܀��}`Vն
�dr2�O~�WGޱu��}Ր�g�6SӢ��y�5U%iYZ������̧������\g�n�\5\�}U�hE�jE���*����'�����]������l4G��?R�*Uut~���K�H���y��^���k��U�5j�3�N�,G��	}^��S�)���r��[�s��W�z��Ǫ֯S-��GG?
(���B�+��{�kwXvL��hW�޸����ޗ��v@�d��|����G[�z1�����Z���g����H�6�k�ۜ�w��7l5c�&�o�u-W�4Ռ]���{�����x[V��66�Y�-�Z�^�*��:.��t������1'�k߶��춬��yC�I��B SK�O飹����|V�4���;����zK�U���*'�?}��Qu<�w�҂ޏ�noZ�����k���*��tV��6�D�j͖�}�v:�k�MqPv�_��6�K�M_�ڐ����<�}�5�M�K�~����+��뽳w��_k�6lR�4�����k7Y��W�����5�d������'�k+[W*��;ϵ�:�7�c*�m*��j��k�RV�����BjH�>��]��\ո�r��0V�������?c��Ҡ��~�޲~�U�3��D]��$�̜vs�������+�{�������e���1Q���k���s��~��U]n�3�3��j���/�+Vڢ��9��fuU���5>����5m:��7w69?|��V���9�߶�̋���1~��G��5+�ш;������܃y}�]�Xڍ����_�+׮S6�X�no�h���8�¼i����i�#�PX���{p�n����t�:8S(�q-J�Ը6&�uk�f���_k[�?'��7�lX�Ռ����?~_�VF?q�R����?�ֵ���}���pQR�U5YH�����h=�{�#�I�_���R���+{�8���?9?����G'/�&'&�+}Wܷ�����3m��f\�^6���3��H�i�s5S��]ͽ��{��H}Ú{/Je9�����׿�pL_/�jM,���|P��)������drL�[���C�_�Hk[Ѫ�5�s_|.d~�W����@�0o|v�~�Z���g�����퍛6ZZC����tm�E�΍������꺆6�ï�[�m�j�f���6�sssZ.7�ߞ3���f�eu������n��t�^��κ�dRKOM��t�9��z��}��?y�-��>Q��*��Z�Ԋ�u��1N^:jX٢��9o�Ȁ���}U;����V)���bkW�n}�]�͛�&��{���Ě�yb���V���ZV���A�w�W?�uA_�n��lݽ[��k�h�B�D�US5�w��Nն�ڭl��z;��b�}j���;[�UĚ���%����ȕ�֦�қ�Vn3�m�C�]�
�"+ʍ��x�E<��._����o��z�-{Ut��?~�"���u*;���}c*W�nt�P�7o��8���*� ����pm*��ZgOg�z�u#����!yw�f��^�@CU,���S�K�W��hӑ3���V�'���~�n��Zk�5%�;�$�U�?�u\�\迥5niSԬ�Ŷ����_�߈g���51?����+��Yc���,�`�s;����֮�x�F�#j^<��Ã��_U�m�(�Ҿ�޾ak5�3��l��KJI5�3z�P��9<�_�tFݶj���C?���W[b�����c�����	��Ѐq��E�Ц�ޛ/�"ֶ��a$�|k���̌�;�ktܺ*�>28"��s^y�@U�F�y]۳�<��������;���&Es4��X��V��jq�_~�TRǒ���+�+c��Ub^E�絝/ګ�6�s�Z(_��������'�'���[�+�|}c�~+������c�~�b�_^=���u]߽q���/X;7o�D�Յ����&G�R.�}���{玲go���֗���+����y�[����Mg����˝�t?���/x��8d6ǚ�����{�J-kn_�O'��Դ���-ܾ�}煗�HscUķb\��RIQ�L�1�\<�OfRz,UIw~���Z�ہ:˟~��Q3���ɉ���I"�4_p�~]��W�~QW���v�~5>>}T���6V�۠���}p�󶘟f0�������a?5~��g��Qu��v�����M�N�g0*�V��l5����~���,��Wv��vo�f��4�k���_���'��v��i}rnByq�>�}�&[�Bb\����A1���|&p��O���������m/�Q?n�׫�������?:��Qk�mZjX����Ko�+E��bn;���5p\�C?��=]IF<�;�N��C/��|�y������ǃ��i�H+;��ζ�Vcc�������2�Q��J���ӕ��i�&inŜ�O������AQ�����vZ��x/`y�rcG��o�N{]��tt��f��yb}�紌S1>��#m.=��~�w蹽f[��+�6�9b�RG�sF�ˊ9s�H�L+��?�.��P8T5��-���S������)�hrJ9?$���߷kqP���A�b~�~�����G��Wh�[�u+�������߳\w!RԱ������F�M�y�h ��޼�n�W����\�e���S�)�g�*h������M�&��wU������ռ�7������cc�V���Cކ��mݟ��,����1}���{ntk��W˻6>g�6��139�]~���OLLhw����m|��gb`U���a���=U�����Z���U��4>�<���7ث��#�#�^m��q�.�1�����P�g��*�v�Z5[,Jm�͖'U�<(Ƶ�M��1<`��z.�n�f5=;+]5�:/�}٬o���>����3�6<?e��c8Z@kTB���]�K/����m�����1˹�[�WG�46m;���[��mkEܺYĭ~�ۓ��y�ρ�̬��W�k����u�Fo���ʕm����#��Z����d�`�ï�՛C	���=��];����ߜ{�t����]w�1��]7���V��C�Z�XQ����?����'RS��ǿJM���Lʛ/�t����f]�ׅ3�h��������-�i�J5�Lz�j�}y���>lޏ�݅j��w'?j��j��$��yi�KfD�7���g�D׹��K��C;�h0 �沵y탾r��ϫ*�K�15`|p�kc��f��q���}�]n��k����?n�g�����'gN��DH/���7��7�b����Z���\�M�k�}��-��y��5������N�*�����'�|�a�ܚ���(od���]�L9\_1ĺ����U�P�q��u#�������ou��cE��X/k϶뿿��f�<��G�����뢯ޙ=h�i�Tc�|Q�B-���FGo�~�ZG`��%��;Vn�׶���W��g@�AjA�]O\>�辮n}n���q�sp�����J{�<&Ύڼ3o�ｩ�p�غj��rj�޵a����Rۇ�����Ym|v���;�+{o_���ЛV�x��\�.�1uH�ՙ��B�f�ʮ���O^r�P}�c�u����8��疾�!ݮ�ɩI����y}�aK��M�������~���K'Tg����N�{��>����٢]��v��;�!�k7mV*�ko\k�ܲ����{�8����N�8�}I�{�Oۺs���9�W����x^�O�%ѯ7�u��.j���7�Z������+�<6��\�j��k��H��ysU󪪈��C��zr�n�s�1������FѦ-{���W�1���U�@�1SI��6���_�jw�m�Yg,Ksl�\\�	�,K�6�k���c�V��J��n_�n�ZMݸ�^T���D,�a�M���������g�g��ݢ_���R�R���3̤g�#�N3���m�F�[�v�m�f�+_��A��+�����H��ޝ;��X#W�V��Z��hWE��v���:Y��G#�Y�_�2�{]S�X���=�+��ꛚ2�KS���C��Ĥ��}��Җ�ٜh����9_Q��s�1S.C3�z*5-����/��`�_�����%b ���?7L��m&5��������L�M���{cP���W:�c"f4F�ɩ9��]��v�����g8�JE**E-U�_���rF�ƍ�
=��0b-W�߭} Uki������r^���>�-�fok�T;a�3��p�l�󅂖�ҁ���6�'����z��[̍k�P(T-<'X������1c��]�gf����q^yn�Y_�*;�S{�V�đҲ���A#cov�BV}u�A{����ggM��w��|�������	��E�IŹ�U�y{{%���B�J^U�*�]ҏ�篬ZF�XV�ǧ�6>缺�Ū��,��(�VQ�T��/>}/t7=��nY-oo[o�������U5W����T�v�ˎ�~���F Uwn��on1����3X����9Xπص����G>E����m�[mm[����gS�L1c�R�Ï���������K��T��R����q]��Ѿ`��x���#�]�o�S�+�B����?����v����(hj��`�V-�7��j0��b^Uż�=/~Z�,j����Bz��]��+K����6������o���5%��/>�u@��rK��~s�VK}�W1_�Jmo��̍���`[k��n�zo}z���% �T,������畂6_�7��9���vx�c溶u�R}�q�O���p(�������4c�?ϒ��r�"+b���3����OO}��i	��x˖WZe���U-�������i�j�:��k���7�N����<O����jJ���nCl����4-gI��{���ݪq��Z�"�b^ϕS����ݰ���'���M�ۯ�]���U��	����Z�������1�}�v5�D���Uֶm�L?nw�������Nf\��_�2������Z�mc���"n���_[˒�n\-��Pz<����L�E�}�w�/V_4�W4�b�4�![JAĭƩ������6{��[֚�5Ր����{Q����w30R�\뽥F݀�g��؏�*Z̏Y�qFl�jU��9}`h �,f�+�z���z����nkkD���!���ﭙ�L�ק?	���@����g����\�C��~/fs�����"�n\�v�ز}�"�Y�*��^����ߋ.�õ���b\C'/�ӶloW��:g�ѧ᪪[�����P�I;zn�:��ϵm�w�����̐*��Oe2�ڻq~��f���Ͽ�Zˎ��C?�7��X��Z5�j��g|G��3�!1n�SgNU�з_y;�u��\,��SZ���]� �aiXOY��]�Jw����c'����������iB�wC�jϻNU�������i$;�ꄴ�[0�+W/����?f�n�:�����Yvճ�G�~����O��r%!�t목�'F&�����&CR(%)RYz�ɷ��������ۭ͌�}A�p��Վ����_��tSk[�V�eZ�������j�-�י��]�e5E���G�.��u�|E˗j������������sCV�Ī"8�8�]������;�p8QpuŒ]Y��ź�ׯ�����И�䢺�)]s�Ί@C�z��;�����eWu�Y}t��.���NQ,䕑ёR�.�{�}i;(�7E�ڶc�Ci�G?Iܜ���l�����64Gr�W�,Z�^2%SD:v����O}�XT��P%W�퉑����'���ez��_d+9%���&�v���U'hD#�'2IN%����!Q��I5_R����?>�y���h��,#��V�V�F${`۞��K������c���~,5QB�:����Ƈ򥲕߷�='FU�xJ��1>�x2~u�?zwr,깮:]�����C9����E������R:��ٯc��w�nOߍ�̊:�9ok���e����+�U۬�c��g��wߎ��ِ.
����H4T�$Vg�bM%O��,�W�t��=�~,����e=$,��]����YFI(9�Rˎczs��ȇ'>�]����bR\Z��l��'���"W�]3�Kk������s�K}�"�,�5�B�JX1
��{)��"(��j��ݞ��鱏����h�h��׭*�=+�g��BX���L����pw�LOg|`x �I�:���_n?��|1_mι%�t�ܜNM?�u.127��+[=UM��e�_��bJ"+&EU�K�*LG��r&~��z}*���͢�C���n}._��TP<�*����k��}��T���Դ��]��؏�m�miq�-���:|�v�X�ٺ������!Mѕ����t�)ޔk�k(��U(����\�l������������C����7_x%E�^ƶʕ�!�`��~�8��Lw�j�f���D1_1�{�>��Fœo&;�vܽ>�{)28v7�ն���N�l-����5%�D�h[�SV����g�;c�g����ª���b�2\-R�l(ωya٥�>���|x������D�R����*���k�2�=�wf"E�*[y��v�tD~q��h�pf�lԹ;Ћ��ޙo��91NeSD��y���y.v�έ���<[V꽠����ۇ�(&"b�(,�\ЦJs�s�;�Nܼ+�"��$e6�Z������8_뫼�Պz�΍�ߝ��nzn�a�4�F�D*]~�q3[�l��b�NՙNO��
����gok[Z6��5���w������-��SR�����Ѯ�؝����U�dr��_�ڣ�Ȅ�т���#�����&�tw4fJ�����4W�5���ݾjK.
�o��h������W������1'��������%�r�*�Ͳ2:z'|��Jå;7�
�qmG���V\3Jo~3�b����iI��𑫧cz�חJX�Ue62j��܋��φ����/׮�������W�̍�_+���ND	��b�P�}K{Ұ�.;�9��ݮ��[�3�S���m}csE,��^y+��qة��yd~*20{'v��b�ݩ����;�|Ӥ�V����rbmˉ%Xl%e:?z���g{�"A,y���&����\v��]��p(�,V�j����O���Kuy���O�AO-5Ś��D�*UN��ݺ��}���xC�-�스�ut'����F.�e�J�V���h�؍�u�#}q�F%���I�-�X8���9Ìd%I���9x�7���4t��Y�D$9��OΗW��d���$�sV�hNg��3=�#��;&R���d���� 3���襷sa3��ʎY1���Xp 5�����l2�����V���b��C�L"�ȉm�l�H _�����~u��Ʃ�d�vvBݺz�]Ι���v�;�1�)�0��no���?�����T)����z!��D�uɂ\(�5X
]�j���H[����Z��I$�o�z5�y1�U�q���d���s��7�z��Q�q����� ։��/��n,)����8��씿g�8;x�A
k1��������ܶ-;�L)�s��jV<�Wow�}t������Ʈ��`"�0G-�0�fJvs�l�J���_X��}|����b*��D��f�.V?��5z+ҪX��<p����y�z���&��+�;FK��LM͖����P8�P���������+�޻����d�nz�3T���q���bo�@ś���ܼ���w�a(53M+4:3��5��+F&�W�R��liz>8s�R���+us�L}ѭ�KN,ȿ���l4!ϻ��cm[��L�?9�uc�@�J+��%q\v�ٕ�U+�k���m˞7��2o�����'�>]1:7ק"z\���)�~|H�v,%���8�{i;�6���i���S�d}d���?��r����|}�)c{v^�RN����u9q�������w�iu��U�+���ޫ���/�re��So��/�u�ZW]���Nf�%WlgM���D���HѮV���\�C�����uw�F�˖e����br������D(��z^I�l�L!:�q:�9��8�OFm�2r��vL72���OD뒞��s��ȧG�h�0t���z	�8���խ+�r�଩��b����g{�4��:WW��x0�"�hUw���/��j�z���+^�K���3��'�w�n*xvL��YS�so�f�ֻ�9��X^�����Ş��O/�������m�1\W)��������Jv^�v>�V�M�%:�o�wu_o����Xi�M��^��էZ��W���v�I���|���������"��ln��y���U{��y��j��T���\������񑙱���z���r�LQ�z �Դ"�HNіly*7���=w��N%�=yf�\Ӳ&�^3����ռ=��	\�;�q���YQ5�c�����ᷲ	=��TG<-%i�8~��G�7�ܨs5E��HC��8��wL5ƛs����%m���D,�ť�+J�F�J<��%;��/����1?nqcJ�5==�s���fW"���7۴���X�mm^�RKjɫ���B����8z�|b$9^�x�1+b�dn����C��9�"�����S�/n\�N֋X#j��1mf-G��/o=0�4$�z�,�A9�MF>8�I�������|����|.Yݽ��\��")��Bծ��r����L����	+ 'D������S�ڛ]QהW��ު�ǣ??�Q]��@��2�!%�E�D󋹗vN���%����293����̍�	wP�ԠҠEͲ�﾿��|�
��_�[څ��/����5��$irh`�ɞȥ��}c�\k�5]U�9��dĺ:�}��g�?X�1����1U��vNoͽ��{���D���Υ����;5ϔrQ�V��w��텃�{ӉX��=�R���{��?�:]�7���\>�zJ5�����热R��ԬX[��dJ�N%�w^X�Sݸ�ƴ�뺚
p8����snQ.���341}��Z;'��:w�) �4�b�܋�΅�[���JI�����Ѻ��T�:�2�kҚ+��e���ٰθ�ee�i} 9���L��������PLJf3妦�억[��R4Ͳ[��7;_��b&���͏��V�}�ŷ�����7�qh�w|f<xv�z��nOÝ�ވ��#ɤ5��Ͽc� #��y6WDZE�?�/i�MM$�f�ca[Q��y���!��IE׊��9S����Ku_]>U�W�x�u����U�����ג1%���fI����X��3_��}y��#���3�l�yEK���}�p):oU��Z.�g�EOu����ۯ�'�h�I5
�wJ��X��V���S&���/.��x�Z�
��jЛ�OV�2�֬�hN(g۶S,�ǯ��~���B2r�Jj�Ѹu��X�'�I�U�kӪU)�@�KND�?�w)197Qwk.�&[��|1�q���Q+Z��XeRsڭ��������H���C�8|��jTf64�ɉ����:)ր3]��_]��8�b�Y���v�)��ޗ��hcRRM?���d䗧?Yqj�Z�2'��*gfS��H8�}�Y��6U�\%�_�K�q�n09Q�kA��n��Jm����;�'��*�Y�K�Lv6��/��_K�#lh!��Y�U-�3	GI��Y�óT�.�L�w���\��;;����������?ʴ4�ȋ�hI����݁���'�޽�P2��¤|�i}��-d�=�34#�L3���5x+zy�f}��p<��E�2�b�ʖCN"�nݚ�.�Uu�d6i�8���}-�r��cj�b�n��/�HEbuYE2��&�3��ȗb��u�Ŏ)"��T�W�������{2�Px^���|��_�=}��q,=�eCv\�1TD����τ*1��V�*i�"n:r�x]�h_C5(�tO�s�喺�x���e�Z����po�ï?nIOD��C�u�Nd]�>ε����BF���jr(����#=q�R_�����,�o�^|��L�(�,�T%���sp������u�j)؟�Tv��Ru�^�-{�&��^s2��q�������d̒�P�̊#e�p��`z劕IEҋ��L%/�Xg���v������C�3��:-�o�v��A���|��w��O^�X7����T+�ؖ425V��V�ͻsa#����m�emd�n�s_�ߘ�u�&����M�%]�1]K;z��9Pt����7_]<+��E��k��M�̖�Dn��5y��E�z�'�C��2�7u�����3���Ds�pZ�W��WPC�8s;�rF����r���ݾ��ؑۙ1ye}C%Ә-���W2!#TrĞ��"Υ�kю��ѡّD٭�);�l�Vz��@f���9M�U����\�襯�o�jJ���h�:�����a��ӣ����bɪׇnFO\;�0���f]qzU)�a�nv�T�F9X�4Ϯ�Eu,5�����[3�u�!+ו*ي�r;��yC�qv�Řk�=W�����!Y�F�PP7%ٝ����i\QXٺ2#�F��e����Б�S�;C�QǱ�z���7s�P���ײQ-\r]�L�ehj,t��L��ୄ'��@f�ٱvK�n�����b+%K�!����'�}c�uC3c˭�S3�����\kӪ�j�Ղk�������u�&b��tĳuzvڪ��/�5�iMSKUǲ�fA�519�u)64;�W�S<e2=mF=�5I�`0�ϔ�x�n8����`:�J `�^�t��%���iE�J"�s�ޯ_������hΏuI���4=3^i]і߰bmQ2�J1���*���7/EO���/Jv�vvT��LU�s[�-K��r�bm�퍾w⓺��dX�e�Nv�Yۼ�<�6]8�sV�m"����vq�z��Pw�w�/�H�6Q�w��l,�`3�Xג��$I�����g���N�ߝ��8�Hr���ض@���B���e+w3#�����'r���V�AI�>>w���Д]-�)���X�^�R0�ވ����倔�l���heqmjJd6)��x���8�J�8�������gE�_:2\�+dS����BK�����(Θ������u���D�19�kA�)X'��J�Ǉ������~|��M�}����H�H��ۦ��ה�;�vo����8�Z�Y�슈����)���&��+6�9�7�7gUY���-��O?�<��1}'6:=7O��ϘUqz>�i&��ܢX�\S�N�~������X/��aG���J9�z8�"��L%P�QY��_���?h(ʑJ��*�����1P�9I��o
����Ӊ/:N��r1�خ�W�a�R��g�O-T�(���\~.�Ź#�3��E�
�ae&��7���vge#���%Ή�������O�ӑ���!��H��ŉ����C�]��;�O�'��E.�uƆ��R2�������wJ����ʖ�9�T
�8dN�L�����w��3sՓ��\ʪ����^�EB��X>��h��3�����R?[��Dd��=�͗ӥ��m�oN*�^�J�c�s��??�ai�b�b��+b�����K2�FҞT�?��Ʀ�#�.�;y�|��{QqH����+���_��/�̉csQ����D��_��x����Gc��*�w��[�VgZZWM{�^p=�rl'x���_�e]��T�e#!E�:;X�w�?䶬ߔ�l��� ����|�����6�r��D��B_Q����B�1S��87y���������[�^�/\)�w����=;�N�]+��s�X_��Y���?�K�����-�"�m�3ө���?��	5���vR�$q�s��.�\��3�ke���DcR8�u�������>��?�� ����. (�t"�_j�3�w��Kf�\!�D����g����G���s�o&�����9i���j�E<ŕ+A-����|��/�1��М��a�Ե���/]ifKٳ��)N�z��t���>}��s��������OV_�Z醤U�۹�K�8�U2�� �/�g3�PJ2�_|��%z�GW+Q��q�T���\�o?�i�O��ù5ͫ��R^��z���	3�dNܕ=M���W��fә\r���|Sc���洎���՘�rM���TORʅ���
��8������US��}6���#�Y�X/����y���J��,[-R�o�U�uɽ���������b��^}-����p���h�P>���Mu���h��_�sJ��T\���,[�;3T�� ����^�v\Y���鎿���E�awuUWwtO�BR�F
=*B?KzV�DLLO���,Z� pa���қ����
=H�y�A� x�d�����2��q�B���ټ۸���hȞ��E��i��d�"�����/��d�n�t۽�qo~R���5�C�Ot���"��/�\�'�z��չu�t��}�u��\�b(��Z�N����bux��<?�n���\�©�u���b�<+C1�ћo����:�qn���ݏ��%aK�&@V�=-G��c ��_������z��0�z�fgJ��R��
��q�&^��k���:{u��<�����m�����yAh��W�!��������g/�(@P a3k�k���γ�^V
�&�Ie��E�ك����0�{p7<nmOL@�ĥ-t]�����Ք�r����<�#1����G�۳�E��%bdS���,�Q|4�'K���hp����A�oGe�J��5;챌�4�߹�f`�m�m{�7d�X�P�|N{$8���Ʒ)��я_{'"�S�m>���͍x�Ph�T�������������sq��/67��vC�/��� �����i�a;��+�Ne�˓t�~y���~t���Μ��w���'d����o�-;�=�|�l�����\�(�n� )������	 ��b�\�LC>L����'݃���� xV *s��$�&�o�$������{�ig&�nEY�d�'F�Ei��y����Y������ݝ�ޘ$s�,+Rv��ft�ɣ��0�E��.D��t�i��x�{ZL�G ��p��l�[d�����(<���5[�h����~/5|�;����jq{�qtۓ����ᶊ�|h>��y� >�gM�Ĵ��L���������K�K��ֺHT���:�i	0��ζ��AqZ}��z��b|��;��a4t/?��p��#V<eZE�y ��N9���O�^����H>;�n<��tr�/
#;����$M��ɻ����������s!��*��Q�x[�a����t0�V�%\i6����`�󴿷���*�
�������hu~)�<Oyo��{�K��jNj�sO�[���|g���o)��q8s���;��p�uԢ�N��g�Ͽ޼�y��t����n�T"������Q~:��̥�xeU�O|e��w�OJ�1��O��<wR.�~�Lo��jS��i<�&�n�I��r�d�{2ޙ�غ |9���qY�2U>���� ��=^_� ��!���=���||��$&���"����r6���d�\�j��l�k��F�Qt:�.,_����Σo�g�O
G.��Z.ނ��<ʻw�����4�xgx`~����c�X�|~�S���ў��ŵD:N�ԛG�IUj��X�Վ�|9s�p��K�� ���$��ן��_�)��\V���c�z���H��������Y��4��;/Y��&_�>������E����Ko�eU������n�8�.�T�E-�%��Tp���������c�$��i{����Tg�ܓse%@VZ�q��I���0���`����h�;�JE��&�=��\}q7n�콷�
 e[����|܉iq.����AFs���3��q��Da�VOɷ�;�j6_zf�_�P⛒�/|eE1y��C�o>�'Χ�?��N�/f�8�9��������ϢJ�A�jD�<���oz7�����U���ZE^�+�R��޻�F�"|�n��A{}����|�@Е�+�W�yY�o^xm*��fU���'���O!VUK�[��B GQ�i���&���hFų��dk���3��Zf�f@���x�5���{o�7���['���+=H���S�T��7T����G���f�dii�N����ms8�r�2āe�Ц�S��	��7^����iE�44~��������ӯP�Rg+�+>����_���M��'�;/�ϧ2�(���

����oG�!�^|c��Q�392'٨��hs0݊
�JQ�H�L���J�o��`��KX�n�}o�[����B�s��eģҩ�?z���h:-׎7���nwZƫ�*��=W�	���Mӟ��� bp�d����v+���L!�,K�M\1�񣯳�~��]��F�EIDn��ێD��<y.Q%��Ǖ�<�:����\}c8�<�%eb>��Eo}��r��UI��CH0��������*~�I��h[����p�s�2��论�q;V�����l:��G��%:�n?\��_ �3Gs�/%���mT�,|{ᕉK�,�:����<����tE��V,�UY~��z\�j���k�t0-<�6���+%����#r����H5��;L���v�w����v�/e�_�I5��!3!�t���d���-Κ~P��>}p��e� �rp�`�`k���S�fq6|��w���|v0>�ݹ<���Hm.��1�!c�w>�����
O|��hno,������T���R\Y9>�������8)'t�x��p��*��%�s�}�SU��e�f����7#BI���l�;7��[�|yQxz�)l���F�$���7fǃ!�8��Lv��hU�jA��}����DʿT�߾��q�oe/�����}-�I�T*�L]?�MOE�����`�ޥĝ^/���4���t�<��[)L٣�����M���'o�?��z����sm�F�����J��F����~��[�F��_3V%�<��n=j<?\_��
0�� %H�矿���d���.�#�O�\�[;z�T�|�
�_2y\U��*�&��Ǘ~8Z�_(�����\��f�$j�p����f$�>��yb\5~}����"v��އk�,�l��|�*��G�c�6��x�?���O~#�;�W[���7��.�Et1�l�4�j�+&�,���ӟ�����ҹb�d�>9Y���}��:l�K9�@�{�0e?�$���7�IH�W�^�=~�rɧ�J���8t=�/����?��Y�o��*��o}�:(+�\���'��p嵍;)	��+��^>V���Wϭ�.Z2R�|]%��珮E��Ë�s1�,�?=�n�x�8�ђp����6�U.��x|-��^�??����{�� �|wP�V���d�n+���֧�?���6����x��l���dr�"�@L$�Fa��|���h�9�=}�L?<md���p����>��i'�1��z��cP_y{�sw�Qg(g�B��l^����o_��ꏆ`��,�Օ�_7��p��"3x&@3�<��8���x)l4ZYX$�O7>���TM}���k\�Cl�l�jT8lvq~ertr�����;���+��|�4S�WV_�]OrQM�si�����q��;ɇ����S%ڥ��D�O�>��+��aൢ�]�?<j��{���|���^�SQ�<�7u��w:i:�����l��<�G������Z���a��_��R:�f��o��C��M��9[Nk��K�N�J���/�--,DQ�˫n6y�(?_���!��R|��M��r���;�v>e	���ǽ��͋�Ǘ�"�y�w���í�C�y~~):����[��'w�
�?F!g��8��9
u_AV���|8��8�om�Io?�/�X0������E��������b�|4�ä߼���RA����Z� 8O�(�W��/��YL%�w��������t�P�jU�a���F�ʒ8Y�^�&#v��q/�0����Z�ȣ�����g�N�����ƃ[�a1Y��2��|^�Ǐ���i8��?��&`��~~������J֐��$s ͡`WWB���V��OfE�l?m\���\�s�5s���K�+>����x:�t�A8����Gwz��d)w��� ����������3��f	/8�)���s1��s�-��ZZ���D��_����r��]�X[+��<-�*��WE1K�$�����/fGG���s�8�f"��x�,�nBҧ�-VA���xiy%9���g����\A�JB+�Ͳ���X��N�h�w?��aoq.��T}�Z�����[,U����~��?>�2����q���apm��BF�"��K.[��c8I��ڕxN���R���LE��yv�{��.W��#�k������$��i��� _���Q���oB�,p�,��	��rR�.ǿz�/bϸ���`Cu�tkp�2!�Ue��"��4�U�'+�/���}y0:���~�$-�>��E�i�3VNX�f�ƅW������w����s���P�!���Y����W�/������|��Z�����m�̨� �+9�u%-�,��t!��Ll�_?��b�~��jRm��
��ϲ���yo>/}.�*�n���'��.Y\�\�#{�>��/���,�--�@���ɖ��/{�a�]�3���mW��$��w漪��lӻGOZ��`���AVmS(
��O�eEYD�̝ˏ�|+9t�Ŭ��s� d�̄��E�������t~a1���3w�ŬW�X�c��B�(P%E�7?�e�8�X���W�Gf�\!Yǥ�s̸��ϲd΂v3� =9��l?��� gs�����ɓ���֧���~��y�I���t�]��Ugȧ�ң]�H���M)g��Q���>��`C������ړ�=噞rHOC���kDʪ�}�q�W��98�A�K��Ak{�ߓ�� �5*.ȋ�>��kH���C�mΧ;�[jgt�vz��d�$���/�2^T��0=Gѥ������|:��O�q'�yOj6�=��	!�b���~������:���~g'��s��.��|���|�"�yy�RTi�7�6ݻ��;�"\b�W���y�^n��*��?��iQ��_�o4�lܟG�7ҝ�R4\횭����O�����xna.���/�W�nα�\��c؛y>���Y����D�IT�1Ym�vf{�`�=PS�j�0����sIDx����Q�e�<�|��
��]%|I��i���q�k/�[����!�8a-*osv(#�����_��p��P=�{w�ak7�/�.�/t�>�nE\��t4���V��.���3�I�=��0b��|�~{����k��\|+v�����^�~�x~{n���q��{�^�����k���ݿ-�-�)����|ռw��j���Us W���`/����`��D�2�8	p����`����ZQ�Ѐ�?K��D�_�v����$��~{.�9�W����t�
ZV�����t��T�����O�S6��&���Z�&��+�r�e�������?D���|v�3�v��3�z���2�u<�u�������t��koΔ1���;��h�{R�ː{�ǖ�J?l����>��O~1��z1s-?��Y����R�E!֚�����z���?���_��4h�������o���I9\�8�*�I5 n�����?�/����/s݅|�D�?��{��j�E�t�u}z�D��۟L����N��$M#q0;m��?�����.A^_Te�&ձ�_����_��pyny�'��v�Z�ӵ����Qt%b���q�������ԣ4�&��|��܍�/�9w�4��N!6����LrS���N���\��l?Zܞ�#rQR����J�?\���_�����!a�\����?]�ϗB'zÑd5�[ݶn�Q�w���#�,�������|�������o5 ��#���Ǣ�P:�%HD��@r��͍�.�&�w~����?�����bڒ�Ȉ�8��9KRzD<�xy��Gow�.�53�*riǴ��-����J/ĥ�͟^���\�,�{�݃h�u�.`�6��@���_��O�~]�&Y��ۯ��n���7��u�P�Ce�50�;����7�%$z1	'��p��<�*]ل��PH��8*��g՝��byyIO�G'M��tuK*�;�����1QL2�O�{?�iYҫϮ{-��>�@1p$_6x�Ŵ���[�<s}���P��Z�R	�5�a�Qkp��ѩ�����g"���)| CM��O �xӌ���ю�G��5V����+���$\������O/=��EQ�g�]*�@���CwM!����(�'WF���9�F�T�hҠ $��<LO�鲔�I���1o�{*.c���@LU��
�@�a
����bv�����mu<;�c�" �.�&km(��9�?>H���-�ȿ��m7qr8V6�J%����hG��Y{뱐�Y�N�\)����)q�ǵ������KO668ؠ�MNp�ѯ|H-F��a��K@l������ {u���a^N��(�I�}_л��nM��&p`.��;1M���wT@��8W��Ԭ����T�s"+S����g`��Ç
�u9;��d�ϭ��V��N�#gj&��H#�E�	�,c�-�>y�D�����f�:�g�\4Q>v��Ӑ��h��{m�8TEE�fN�3H7�k�#�g�������O��+"��ɘ�X��?�,���ut�s�ᷗ�jkE�3��O�ʗ�ۡ@��4SyT��C~��x��A����
���Ђ1��JDy*�䳶��;CH��*=��>�;�*�^���?x*�A[��@���R�C>�
-U1/EC6ߜ��pr�T.G4�d��H�(��r��i4bM'��s�$��e> \�� /�T��\~��W�v7��\���ɤ�������I�{�#�f�fbp;�Z��4��DNFK�"UC*�kE<|��Ha)Nn_Z��O5��4�I��
�	rQS��et�^X��漜�c��)�G�2�A�r��:+s>Ig���#A��vO�i��<�|?cy��Yr�V��7���_u�cԨ�t@*��%�`��Ǌ����;��d�j|�'^iS	��qJ��A�Vw�3����R#��e}ߴd��AA����zy�L����䕕���JIFB��\3���4`��X9��*:�p�̈́]�[���ň���>o�fN=�q�2���;�N_Y�,�q<ѩ��A%� bEPJ�^��n�����2'��~8$�����.�,ӗ��>��b�_;;-N]GM�>�ͫ(k2��9AɁ��R$�����:-LgR����t*�r�ˍCT���~����~�+���}2�@Bd�4dHX�3y���֧|aa��E�Q�\垠UC(�mRA	k}6���G�\\~�A��tB f�McX�@֡�2�a����O�l�7�G ��l
z�|�Y��7�bKZi�'lv;��tN4:r2���zA"��P���������o-0Ȣr�M!��2�u�¸�I�:�t�v���b��+������«\�+��{pZ�E�_��=>�)!ȝ���ȗ�j*���H���P�>����\�-�$�ʜ�o0Q������섈a�����tP���J	ꐃxD�����1C�� \��?��Go-^X�W�
���I\�E�q�[� ��������3M�<��1/Q`WF��$�7�Sia ���V��֘�y�i��%�� �ҠP ���\~Q]�z���[Cb��c��}Qy�3[ё���o��{Z��?3cQ�8D4+^ba����>#��ҭd���E��u�� ���.w+�d����~a�y����9��틖2�ՠ���ʫ[w.m�U�V�:L�z��Te��h��0.�!k翿�y�Ԝ/[������2U4�O|r��S���2>z>���:�M���'^E�ȵ�\�u�<��o^<�
��	�9��~��&׼A9F���/���Ճ��Ҙ8��"�'�QV%�6�F��xz}v ��I��1��?�\�4*V5�	K�^
��x��vG�j����t�x�&9��̓aTS���/Ŭue�[�{4x�A<:��F���d�X��q*�a)�G���N0��b"�@nIeܐD� B|shX0A�l&l�Y�^[�TlB��̚l�8�	�" SI��S���H�:�
���18Ϋؕ��)���o<?�e�V���\%�����mPQ�C��E�E8�Y��O=	
_G���R5 ��Z]'��_Cq:~���&��� ��|� ��g�9�#���o޻�sx� (�~6҉SzI�KDClǧ@B��,+���~��5�����n�'�*}� �A% P����<��g�j�n ܤ"d����d��^��퓋�hT��t�c���KU�j� ^<(Dޤ�Rj�0$��lw�o��VO����DT�yC�CʾJ�]���蕇��y�ђ �7R�6 +�C��	$�@�����tR=�_/�z=���N�U胖Z%�� �ц#ag�?�q����k�T|Z$&5��h��c4� +��U"Sy��ϖ���;*�99I�>w�WX��W:.����<7Yٳ��j�;/�ُN���!@�Q�w�C���(�+���k˯�**�n�O#S�MG��� 6�����7.n��T!f>�_7S�c|��ڰN��Yh��4bO��KK������L�W����� �+(�����&`l���(<���$����/�&���<\=��!E>*C==��lq��d�4�K�[�^8�9�f�v�aqJ��4 ��fW `@���Y�r�����{�Ŭ��i:r2]��_K݄k�ǆ
�����Z�W;+,��ThR��K�7 �@�� c���<xtast��B���Ф�n2�f(8��8dL8'�@99��p�u�]1LH�>♠�y��w�F�*x���'�Ϫf���� hPK3�y�821W_o������%EnB��x7J�
H��������7�tq�s!���cr���@^Ѽ�r����eP�|�y��ꐝ�i�O@V9�`Pf�p !Z84��r~8T+�%Q������r&��$���w���^ؙ�Rk��O͸
�ҭ��-M�ϘCѮ��l'�O�;U;h�Q8%))�«�p��0�#�PIU����kCfp���Ư$oh! �C�3 ] ���_���#_y&J=�f. [�-@
�+�QT���xup7��<�.3��19����ڒ ��0�+p�{�O>���҅����Hs�A.ص��q� h.Rz��QŏƧ|���*^舧���)o�-A�Q�����o�'ǻE�k�q2�<�B&���w��5�E��c�d���^K�'�$��9� ����*������Ƀ���X�g��$>�f	�k\\�p,S2z¶��`�b��tXF���� 7A
0���t�~�ʋ�'�+�`W��C`��� �
p�Kh1�����������V[��t�-��� �)�[%����1;?wA չ*i�2?7�t�j
�o{�x\��t��p��W��$���-Ae*�+�ׂ���LiJqe�>�U�vG�	�B��%ప�H�� 
^��%|t/d���D,�8&�&�L��� Q��2v�y�݆c33+f�Y��� �}��lܔ�Z	���(��ٜ�x���.��_i���.�[�l���9��'�/_� �Ñg'SpF� ��T6^�`]��7W��{�<.]���pb���B�.S��ÓW.���W�����s�^��!^Cn���S_m�=��x���^혈^F� R$�+�7�� w.���S1ט�SY8��!�W.��� �f��D)�w��ω�t�C"��X7�aX���I��Na_K+�`vB6;��AȰX8�4���ח��K��I26�G!?�ȯ�_*ee�������������(�KY9�l�*|���	=|;��{�6?:�_8��O��|��:�cy�֥ ߺvE2��������^����c�Cd+�;�?�`O3FJ�4ĝ����W朮�S�v�2�$�_��;�?��f>����h�:r4�̌\�8b��4�Q^A�s�v��?9��jtH��S�40��y����R!?<~�O��~��*3�2��_BlǺ��u.��<W{���}t��u{db"��"ƃ�I�~vE������������R:-lMRi�k��.��iBκ���`[8�Qc5!E�݂��1<��)��S��A17�<<��Z'���e�V�����9�� ��H�b���x��	k"���A�X>0(I�& +r6?�Õ��]>���=��r�6�&q�׈[)�O�;���xe�=�3	�-)�[��5�`x�ǵ���~����ӭ� �d8jV�na�< b��������݅���7{]���C7�r�%�[=�A�KA��P�<���ps��RD����>�D��m!�A|,��{_,.�]�m�26(���Da�+�B�N���٩�6{b4←��_��w����AV�(�d=/7�rgE���8�h� 0J v�sC�RW㝅���|+ Ho��cZ��=�����LBC�����׋�_�@����(9q��y.w|���*\<���������K�%9.C�?=vY��ܮ�*�MB��	|G}����� ��+�7��c����|Ou�I5wp�����k0�e�B����/`�� ���O�_��=9�Mk,V���XЀClw�B�q����]�ܚ�v^��~� >�eSP���Z'��4|0����D��	��W7@?�+.ط��`r���b��R���R}��5s�-R@��x�� �_���OW��nV�N�o�F���&�����0mmBU�Ӈ_�{�����i�i�Ij�-������o��_|����{�奋|kwmНЬ	���C`ti���>�/!��?aO?6��-7i�ć8��"��T����_^Y?���[/�!.����'A����M��s@W���fu�����?��γ�X�����S�i�l����J�@���P�����d�*������1�w����rQtJ]��m����%��2/Im�7(m��#D��?���|���|� �ח�u ����. Z�F-�� �Q����+[���[Fbi�M(#�� b� �g �g�%Bs2��ѐ%D���	�_Jc�8��M$�v|��)�Z`��j)��&|� ��7�OE
 {�����c}g������Q����MXD(��G��p���j��R(
8�Hv�Q �IhARX�i<#��:�  [�c�-w��,��
��$�|l�]!�D!�u(�x,���j��h=$!99�CHۮϩa;I 'M5��3���7���H(D<���Ua��+���H͈�M0�tp�%�@IyD9��I&�vmz�#��)]�I��4,���jϘt3�b{�#H0 5]��q�q�]>n���k�@� '	��s�('��KG��I�W�L�W>�]q�7U��Xϵ{�\a$"�QL�D��a<�V��x�� $#\�ra��3�2l�SS)a_8�{i�
�%Ln�� ��7}��ڋ�Z�aje��p� \��,ڴv���
ؿ�c�M�7�[pn,�f�xWj������H��
~3��TI2�~ �~���������%ȩ kg��I������ �h6(|u7�� &Ni&�1��V��>Ų��j|+���� �X���*����
�n����
21��v��\k��g "O`]H�^�	�r��/��{�x*�k�xm�%�B�,A����k5������c[pq���2��(��	 �Q{>ܻՕR��23�)�\�((z��eX}�S)9�"�+�D��u��P����̀	�}KKc7Pb�ɠ���� �
�!��� H��U�4F�+\+�oIP2�x���L�b \�k|�/�����@��F;ɫ�. �B��u�����j+Wm"��I�P/`W�hW��4�r��R�q��i�+-�T?��<�6�־t����/h++�1���m��Inv�ko˧����g�:Ю���h��8��Tm�~l�Je@�X�I'zfN�l��ڠ<u�xE�cXR#�d�f�[�����^�h��_�]��ñ�9�Cb�?\���l�2(�/�B����Y��l=��I�2���A[�L���9�@AhL�������:�p}q(�JU6�vL:p�))��86x�W��gֆAr�� �}P��K����2!�yfp�&�s
��G�r0&�?���l
`j�WsC�+��X@| �Jꥉ��ˁ���	�x�R�X,��^�sJ_�c1#��7A4�J	���Im<詘7I���K�(�z�z���¼C4���f2=MCk?�JW<V����ǝ� \�P�H����5�*�c�2�c��!b��t�q�S3(Sbe��֫������Ò$>��?�Av6نH����SH۰?|��eR�Q�����`���ZZ��+��%!�F��u��R�*�s��8��pj���m
~��:���
�G`�k�r��_,�0����{x�kў��[�_9� �L�W�F!�R��(S�C0b,���B��!��M��	:��u惘�ȃ�
�(����T�Km�����}\c�g�W�V}�c��V�O_�6�������1l׭c&H c��*X�?b�e����p�k$���bF{JZ���e����J���%�E�; �Zׄ�eFNq���0��
>�}��$$��c����=�?e�.�/�n�:g�m�3,h���5Ѓib��W�� 3�� � �QT��ͭ�H 7|U#b&�����hR3.3kg�f4��.V�@e��Rr�+�C�s�� k*lr`��L�8��
����"��e%ȅ���%fq�u�yr �wF!T%��xC"n�����X��� ��:u46D�͹��mp�!v����@�fy�Kq�㄰�Uc��1�R�kq
�����b��F�vj��v�We2.
�S�U��!Na~��9�%%8L�� ���o�K�z+��qS�kq��"�a��L�^��/%��-q90n> (w�8l	�AA[��
y����`�R�7T�R�!�{�A\�}7S�C��yqy#}�ף%ɪS�=���9���ub�@�
0\7���!"��@[��zu�W`�#XW��I s�]Tm����m$�u���Šz��R6�(e�"���~�@�!)L4�%OF�6/�Wnc0��#nN���9d�9���W���0��C��m��3s�"��з���]Qk#�T�?$x� �4ȱ �S���ޭC�=��n��iZ$ ��,D��3
01�@a��g���x��������M7�-'d��q�v �BdT�5%�*�%�Wc���@�`|E��Xd�!�$�+�q��_�Đ�ce�!^|j�!6�K��1���:��7�B\
�W��	}f��#��);���!��rA��C0�@Ĳ�������A�@��i3,�_��-�F{〡r5#�Qll��a�Z@���F-η�)q���E��܋xvC�G[|��K�N���kL��7�s� |����3�ǌ�^)�%��;������*��Z.b�7�A��$�Ga!�4�ǀO[C=`���\#�#1;�1e";0^��b�~��z�����p��ì�W�"�s��E@�L������*ns���.hR�kK���3� e��c0�gis��\�d�fQpv�7`,��$bo���k��w�� �!��#�I}��bH�v����*������1���#꾮�k+�a#%�<7|�)?��T�~��7�/Dl��&�des#G��MQ�w���<�B��c��Y&�5ϳ8�,�-���%U33 |c���>��%7`��j���9��N	�kD��+8X�B'дFc#S��(��Ŀ`CXρ��D�M
6����CId�
1�0�Ե�#u� �
ߏAD�%��$8m�@%� ���9;v���pӨ	�e�}-��"�l�$ք0�lʁ1'c��B�U>[,H��Z�;�)��ī� �U��m\G9a�m>�cS94;������X����qE!NF�M
�)G�j����x}����Ԟ#w�ݡq��bv|5'f ���8�xm2�+nN�����,�/�m;�7�/J��#���p��ɾ�+���^��pm��לB����eX���a�M�|-�[<y�~TňO�z<���i����C6�����Q�9Xϳ q�*�I�`�Qy܍�l1�7������q(�U����r�7 Ntj.䀭�Xi�E��v��_��*n�9�S�9��q�K����o��I^�L<��[��`�;�OTL-��x�v���@�����J�C�#	�ɩk�~������W�����of�)/��4�E�
���0�`]H�Zy t\Ol]O �5�Zb�`0�i�6&���Us!���{���
4
�~��&p��mm�,��֦,f���;�J�E���x��v���:�Xk$9�c�� ��!w6��/��r�[r�����K�M`\����-�ֳ�@B�~^�%gkz��Z��u�d�kF�Af#w��f��Y}��I[�$�_1oW`��6�!����Z'�ޱC.FpX:�@����m�/HS��l��5ɳZ��I���lX�c�3>l�q����d�W�Dh`Xk4Mm�4���ژ����$�@78��3Q#6�Ե+;�Z��u|�Ԩ��X�hs��6�X$���2��C5���%�4�_!׀�L� 0h�~
��^�ɪ�#W�<��9����X�Ǌ�LTATO�<	6�m�΁4S�h�(m|��fB�)�l�vl��ce��9 ֐� B�=e��jkd��Aº��n_�m��m\�a����=׭�jp��[��M���X ,������bj�
�W,n�d�4Xշ8�7��_��"����>y<�78%���W��_�W��ao�4O ��}��ϰE�?H�zV�9�u�����/w����ڼTu��6�Y�f�1�\O����X�\��
�Ra�W��+���nQ̭�?�?�
���)�21* c�N������"�@t4�;K�Ծ����?��??�-� @�0��q8� �r0��x�:�� b���� 'H40!"r��7�B�&�'1���10bb;�Hr�zf��X�ξ��u����\d�96��gx�4��%�%�����, 0D�9�w�*
���Jk�9�.���%�<X���bAA��d#��Od�+Bf,�]C+����n��B[v�u([6��h	*�Á+��%��hcs���z��
���q����zl?'yد�;@�2||�Y��H��S���JcQܣ�M���bc,q�J�	S d���
ǵ��3us΃�!�4Ʊ� <I�9��,��&BDl$aM�^������+,`���&X5 hZ a\c�)�B���+j���~϶�\���w�fY7��|
���}H+��;�	�m뎛����x	,Ѥ�U�}i�B-����" D����G�9�6�`���!��@���0pq�=�_��L+!aA6^�0���:.������zג%��v Ă���Xy���: ډ�>���"��IWl��j��[��į��3l*z��g�*�p���l��.v�p�۞��4`G�*B@h�����-3$#�αE�*���VGXH5u� ��U]�����C��l��'���kQ]��;����`��E����B���\
ۤp��3"mV�6�,b��Ҍc׆v�E$%X$%>> ��*4����Ae*�.\[4`#Hv`�v���ʟ��5oT��c*�W]7�������i��i����{�J6�`��E?C�
�6Ȭ_��KI��!�m绂��$�hkT�X��Z��;l�XrE����=[ܲ
�V('��� �+Z����~,�ca6nA�'�p<�U~��ԅ5�<m��긌�½�f,6�]Z�#1���O`	�؟;��ȳBBE������a���..q�r��A�-ܠ��p�oԗ�M�#�Ɂ[��u<�cG���wu0�J۬����"?�dl@������8�� ��q�2ua��$�ne� �8���ب5u�
���uq��+��RlHQ��#c�({�5W�cs8��=��q����1�ɶIb�k���XP����D���~��Z��z�{�{������d���
UR���Vl�r�l�(jmm@��T d��3��Z$�զ�qr���3���dM�}�tla�.ح;�*Q �j<��5X#�p��z�YQ�i�W�4��uR�c��HזamN��-:�\�q��ΣHeP�t��ym�lٽ�j*��4��M=�Rg�������G�3�.�A_���u,Ï�)���c	��)�&��<k����\�賵aC1!DTO'�z`�ځMb%0B� ���K,�,l!�2�W�sV�	as��P�(��l��;�P'lZl@5 ���b5�j�9��f��L�d �)b �Scm�����]Yp���N!pp�
ؗ�wka%�����{r-ީ�a�,N��
'^ѯ����8mK鎱E���V;�鴍�g�YS�i�!h�%��`P�օٺ���H���W\n�)�X?��@appѵ�������{���
"��*[^đ@�\�2��c�_a�Y��Rڢ6��z�����5��g�`c�X����[�Kj��8]���xG����b��k����_���zh=o��4���t��-|֣,6^�F��A�nv��e�%D`��"�-�����<
�v�0=k�#ni�:�r���X�x��A��"�Qv6�l��yj��ڵ��:�Fby|�:��ě��ک-[���P��z����k��x�,��1�a��^c��ܜz�������}��\^'|���*\�G�]�☟�Ќ8���U�ިm�"_ж&���lg�-o�����}�y�#��4�c��$����b+�����8x,l��f��,�0v�mE��ʎ�hhc�k��6�"��[�g��nq��K�K�x���� �n���zH�.����6m�k��R���YxJ5�~iY�������kc�.����q�-��pk�S{g=�Zs��E߶�C�e8�Zs](��r��%�!,�,=k��+�gX����kb����ü��9k�;`�Y�^���cv�
�j�Nߩ�g�g��"l�ú����yg��w��)`G�
��ŷϒ��zt�:��b�
���)^6rZ����7kg<�%�U4ۨ��!5OA[E�k�Cc�g�^�u��7R[ [si�W�i q�Y k���Nmӱ*�C�g�
<o���3�#vpl=� �����(iPS�[����ݱ�X��r�8�M
����3��k�������h�J�,*G��}��5v� �쮕�m��a;+7��G����mR|��{�5�%uCc��u�õ�@�����
��y^��g���@m�":�r9��C���ͼ:��zh}�6�-H�-�m�"��[�+;4�lrkP�M��@46�T��l���[�i�k��8� ���&u��)��n�'��h��]�:��ځ��������kL[g>�ɊZN�mc3w�y�����aL�:	���P�S߄�i2vp�6��Y�ڦ��8�����cuDkW��� �x@��Xa#�Š�TD'���ؑ!����m��;�P�w!,N������c��x�n���7�Y=��r��x^#�� ��2�g�}
�W"�O��AHe�.�È���x�>8�p8đ;��▸E��D� �9d;W��j���7XԸ�^3bA伸7{#�/j;@�g����F�S�F��d��mF�3��������W��#9㮶�tVנg�ݎo;���`\v�1��\���]ͺ�!�_�?�y��9˯�mk���7[Tv��ZB��<����A>ȉ�)�vh�;��yP���^Z7`��:8��zQO���-q��]���3�>�;�C�j<k�ֵeac�t�4�n�Y��Z������÷��j���c��(b.���FT6�R�5����l�j��vn�/0�"��<em�ZlaoȰ��z ���[��Wv s���k��ȿ��Ņ�Z����N]r�2�g�h�0���c'qo�9T�SS�������g�S��� �foC�$�����M�uIv�2�9���Vuu����۶�9�0q 0`�G`;  ��� �8��lal0[�d��jI�U��~ܳ39���Yk�}o	1h��{��g�̕+�ǳ>�n�.<|�뙾���wOnm��������VRU���v�K]R8�/�����Cx�߀�^�Z����ז�?M�k�W���X��m���n|�x����ђ��d��~_�E��(�iOd�y�v���>8��<s�[�>^��w~%(:��_{[���~Zc���@[��j9���l(lّ���t�s,^YE_�	z��`w��e���7�݋n߭}�cj��
[�1�������}层��Z~���CM������6���T��c��G�R.��ݖ����}�V��ûcPb���=��Ê8E<|��Akw��l��>fw}���|�?�u�ʲU|�0�����w��@���6�|���.#�6��^�m%�\?��W��2��y�����}\O�u~X������?�� ��f����y�^�������� ���v�^������w�ί|�O�=�����6>�j�rw���0^ �땋+�\��r�p�?�� ��,�/`x5X!��OK��xXF�!{})��!v�Þ�1_>�]/����A��]�ޅ.WK�U8���ݼ@�%� D�b�L�u��8̄�{p�e��g u�=Ǭ)��p�
-{��,�+, `/E�y���Se�y�I7B@��0��+/z���L\&�rDW�W�B���>����_�]Z��|��CB�c��L�����h5�I�DϬ\>r{z���ָ���AY .7/��q:\��{��Ď�/*-<����������Vf�1��HF�6� ��XO~��pN�5}��.��"д�1O�����NA�I�ټ:���Z�Q��'�-˲�p��eL���c�\���nwCǍ���ޯ�]0]]2:��P����L-����lj[�s9!^tC ����Z��=&�h�r^��1����޿��pf�x0���'���SuG�a2ǗQ�x��@�m�5���+��t@m1�W�l�o4�=�Lgg��2$j��lt'��~!º\X�/hw����op��X��_��w����.��.���5v�������!���^���N��:��ƀ��z¢����|�m����-Z^�u��{0��x-м\<��X���������$�$q>���>����J�A�ߠ�����=�"z`�J�x���|�l�r��p]����_+�Y����u�F��uar����q�����w�X`��c�Qg���iy�^Yt�|�	� ���+'o�}5���>�	��3��̿8`=�:�}�5� ��ksFI�J��U�|�� # �9����f�|�X����u �k�2V�T��1�c	9�J7���!�4��Q_�E�InȖ��}̫�M�E��%�>�H��*���I��7#��I/LPZ�T�9�=��H�^`��-Q��6�/����|�B�>8�7�)����0ȃ(^�
\����L\��r	{K���6�iG���X<����:1/���
βWV��6.,�x��|Mg�>����Q�0��ؽ��
`-&RH�ks�|r ���@B��z���0w28�`�'�ޫ��u��Z���n����,�<<�:#9Ń2m��u���Z��EN����0nc��`�7� M;�'��.4@��sW2�y���G��k��`<�k�������������� �t�F�b����z��
��;d�=��o��y@�ұ&��޸��겱*���v�q{`~U4y�=����ECCm�L&W�ಽ�d ���%�)�����u:@[�0a �N ƫB��>>�%&�*a{�����-`z��Q�:}�/����a/���$�"ظ�����>.�� �� -�T�~h��a��,M�#��P��{����"��z�������W����<��?���Ɖ '��m���10�׹�u���O|t}=XIk.�=����{' ��V�`�w�Xɮ�TxM&����'h�l��t��R�m��rF ���D�mhӵ��?��}�$�~��m.Z�V��s�O�'��{y���cn�X��} A��ھ�t�v�� ���t�����P���=�vxք����^>��K��bJ$?"xJo��? �k0ɋ�SYz����_+	iɆ������x �F���}���
�׫y��s����0�:w�D�� Ǔ۴�_6� �$�y�]��[c2�-�!�Ġ/���=���c���'�[�����!��]μ{�!p�$���=���[>�t�V��Xqm��9�����r�z�ɴ���kR�z�ۄ,V9��>-��w�����3:��$s-~B�lv��E�֘���K���rj�EO�4&"z ���>ٸ}\}e��:�Iy�l�U����k��|/���&��X��|���.�1k\���@?"Ø,������`�/.�ah�>A�,lؤ7�������Y���eҍ�@�����z�5���F�[Cu0�\n6�V���`���A�^��7���s�r'����5���4�0��5W��J"Z����X ��?K_��95G7���m���.��� ��Q���u���^�$!��	�F�)�v��pPz��NS$��=!f6Op�HBr_�����<A�7&�@v,ُ ��+t���J�����F��^�'+u=��!P:h�78~��jwo��W�ф��l�U0�/ٙ�1:�ZMO�_g��Eϧ�^We��q�Y>؅͖�&����%�/.�s��q��sjL�6���1J��&l7&���-v݈�y����Y����9.J§u�n����ֲҜ<I�E���[z���ū-�I��)���C��o��|`����K����Ɉ7{{� ~����KϚԵ�-�v�o�.q�=$���`�vw�SN�`% Y�L�fH��=ic�˥)������	�p�!�#�C:���3����S�3ݐ�rx0IH>�ĵ�KP	d�߸�w�������°`����@A_x�j�'��@&�B����������x���t�S��\��e�x�|MC��z���&>
}<����-*y�����i��u٤@��iu$h����Y��'�a�xW�;�lQ��F��9��߼��WI��\�5�9i���No
��A`����'>e"����av������M���'��_��p���l��@�}e��jH������;��:_@,�����^#�ea��	��S��v���t�h�q����YgcRϓ�s����\ǅ�Q7�4�e./���tuC��`[��'_�)��ES��d��
��
$`G�`qu��}bTn5�����N�x���G�E�����xų`�ΝC)��� �ǻ,�f_��9�[N����	[���a�ZG�}^ ����;t���S?��z}|����ݽ�^�x����z�^�?���� �o����������7��~�?_MȽto�ӡx���T�.��*a�^�!�x@�vԝ��z,�B��_��.�7\��5�Uj0��4d^�Ax�DF3o��qe�M�M=�M���r���=�_F���x��r<��p&���W�򕗢�ܘrE.Ђs"��e3�X�՘>�D�Υ1�g�yV%4�+T�#w��Pm0��������pa;��*�ƀ�;��"����p`��2���羐�4�;��nQ�F���Y؝Fܸ �D�څ���) �Ƶ2�I!��s��"e�*T]�M_u��-�;�57:B��,�t
o�xl�;x��+W����'xp�y���Ҁ�-��z��X-����󯠲� ���J~�+��,�2��9`O�w{4���P h�� 4��r*V����>�;7�Q�@�`�-x�Yk���@� �р����[����=��d��|�zآ,�sP|Y^ ���aG��a@s�k@ @�B�����r�hh��C��7�*M��˰�C����h੬>� �wLfM3��].��6�X��������=c����8ݷ�\�0�=�س�/ �V2�!��C����1�E����ASw���h��?�BN��� j�A�AمJ I>�������1�d�A�[�mz<L�#�D$:����e��Yֆʆ�%��c��?8ۋHf��8`�d���r�}B�tʟ�3��K�~���M� ��z�L.�ޜ����;ӫt��b+���"��I"�r| ��{B�� &+LY�=�&w���}~XĶ��}��ګ�<X���g��0��v�b���$��T���+4�!���S�B�����}�`�Y�v7_I8�^-�gnNb"�^ڠ���4�Y4X9G H{�ȿ���COz�{=d0�ӑT4����J����#�	�P��73-b��ٗM�Q�M��+4QX@�F0�_DCґ�.X�^����޾l��/�ս4@S�Xʭ����".n'�IaHYxN�'_H�#@=�����ń���uʆ�g@�;�x�����s�A�3Ό��S���e79�=>2y�mo �`����``�Y�m����0N�hW{��ƿ-Bnau��d%�ԛ8{i,7$�y[��䔢�v�vt��d?ڽ�c޽j&m}%D&�c�ڠ�&�Ǻ�J[��a��D�~U�Mw�rJ��L�	:8m[����q�(�{}��jƽ� �A�A�P>{�v|3$�q� /����b�m&�䗃��[�v��_$������e/u�����aݥӔ$8(7�t���2 *��؁6� ԝyૐv꾍{ş� 3R���������
�R���֠�c�X�R/-���>��7��E�f��Ǩd�#���*�ǆ�i��� Vk��v8gtp,��l�t��7�~B`:ǻ ���M�n�'n�3� �������� b�Gg�������5����]�NBMb
~{�@�\Ѝ�B��c���J[X���Ķ������ �HpRR��l�7�`�]0j�ú�&�}ӃȾs'�QC��.�B+3���H6%�� w�א/���A(I@��� 7��������:����t���<8|�6>���@Aln�����T ��#C��d0�<�t"�yҏD�@����-��C^�O��R�#H�q���7Opԁ[�X7�\_�6��Fb�5Oh��7O��nH�ž���qR�ҁ��f��2��<#�r�:!W<�8�ʃ�i
$5tzX�wRᾎ|!c'E����0`��=���;��l�C;���Pb���9�d�yB9�,H���7��c�_��g��]vTU�ӿs�q��t�V`}N����	��s�7���#�w(86�;��6JC�AY4ǌ���J{b�xE��Q>7������g����>���;���5�G�v,��DՉq_'�]��װF���8$���tA�\3&��<�����1q��;77�t�Œo��c�nn��ֽ����ox�(�Ad9i뚔�=m(�-�9^��u �
r4�G�x {ɩ+ʕ���a[�&[xY�;�V��܆�L&���y�d`�OCÿ��¬f�dQ_��5^zą�x�z���Թ�SW�C�F��<�)�9�Έ�wŚ��&,M�l�6C�:_�VY��Z���B�:���\zfx���2��فh�K&f{z�4�;�u׵�H�*�;����z�H�1ڔ.�Wr堌r̔��&�� 3/�#�`5pc2P���>�Y��W�!��c݌���8�o����֡_���˼��C��hS�[4��
m����g���&#��~)�Ɣx?��5�
׎����-��n�q����7)6��`f�xc��&D2��ZSG�l��L6!�e0��F��r��$=W��&F��JWr{n��b3�}�'�{Cq�d�+:K�VF�	�)��s'��|�I;� ��&<Ø�p��M�L���h�	Lr�|�m��Z6\�D�F�|�r:�9q���i[^�h:���!�6�q�����,�a��G�h���֠�шc�]�k_�/�����|�?�w��/}���Ͼ��ˇo}�[��z�^��돸~�	 �����'����|e�~xk�O==���*W7��*�A���Q�� w�\���;z�T��ǋ�F8��3���" �B����f4 �� �-�*x@FJ�@�R|�	��^BMr��W�(@���jCc��P|��Z�]�ۍ�(d&Fa9f��oi@6�?zf�`
>tV߸�¿�T\���<PmaC��q�w�6Pd��Z��,�V@f?� V퍊�<�#�;�֧:��N��
F���T@�&���ϲ��\j�@.�2�*�D6�F�A�)f�z�0�1O_cC�T�����e�-�q�	=�x���ss#a`ok�Q�!�N:iO��?�tT���ZUGh��H�w��L���+�� �XpqG�٪���{�Dot�A `n2=�j����:׳M��
pt%��⦝�A5$7�8�2�����#w=gRސ?lk�O�[L0�˫[�hw�t��������Yk2����	%#4Vp��j̰��\��V`-�	�;k�A���G�8��E��C٨!��/����t9HG�.���tb�G0�d�˩-��:�:��-�n��Q��厎!�0���p.�󰷃g��s���R�W@+�?? ����5%'�z�R����f0I�)�@��(��kL�#xK2��#j;�I+�����b����74	d<���~��7�Q���W�k(�).�,�	�Y<a�ZӸ�ܳ]��Ƥ�%3�����m$�����)C�4�`�Bl��vJ���K�oL�` '�2Zt2�@c���zf��f-6�N�aF=i��3by���3y�b�]	ЏU�c<�d�c��C��m�F GU�3X� 8u� �%����U�.:���m\ȍ6�`5�0�Ⱦ���I7o�?Օ��oG��A��;9���FS��_�wPO'���L���'
@�
�s�
�#�7Yt���\��}H$���3�#~G�ٴ�l��i@ `�L�]���=d3��7%"�����	�[�;u\��a�{Cv��� &m�<��I�S�������)��Z���ڢ�|a���d��ʦ��M�f#ǡ�v�����!�c�oC−���=A�2׌-(Q�)��`c�f0��}��0Ӡ���ϰ�ݾ�%��̔p&^�~aP��}W]/m2�c0ik�;���Zz ��-LF��NZ� S��n!�ե	��Sm1(({����X�c������~FR���L$D+T1�'�z�]�����SH�e>cXc�Iv�������N�t�;�N���p"�a�8m�UR̓��C�-�x.^���u��H�:�ߠ���΍>-�G#P:�w��\g� �U�;�����:���Z�o����O%�YTą1��^[����Ic��;7pQ$r��U֭jE�ɠvg���]�4���%kUjM��d2^ʾn
�����Z$��~��%���ڰ���c d���R�]�w�=�b,H�Ď�z�����n��1w���Lf�'��?�!V��Z���Q׭�v��e�:�h��o5�Ma!K��&�u���4��~�ґT��;���|(|G�JT��P����g�e�T��O���b�G,��Gs��ؚLr�t��/���H���(�6�i���2�}&O�������/��W��������e��qm���0��F̄8����k��³"Y��q��i�1����(~@�ЉB�v(l����>z�̎-��[�{%��!;_r�bJ$Ҟ��~1���Zj{&X�n������=���]��E@�#^�s�ش�����i_Hփ\��*�����F�}�|]�x>'a{��%?4_����]d5��H�j~��9U{�Lc�'}���@�M�I=$���7P��=g��$��\�)��]j*y�vC/���&�A,d�������E��V���Ð���D�����AX�e2�L�>�q�1�g����ڸU���Ph!"��[T�'����t���[ѣ��b!5���8a۫8�Bo&���|%�NҎ��Vr�z��ɓ�L���VGǷ�#���x[|_���f%�p$L�&���߹i�0׮"hF_�~��j�B�"�C�!�]������N��:�S��G��᧎Yw�B����כlB~0$�K�*��w�dh��Pd �� ��7ni;�S��ą��{Ha#���çM�����á^$����'8v�-�,:;�M�l��E�-�e��(	3�^��-��	�S��|c�7�y�<�N6�����>�ˎuV�&T�4��s�h�mҎ�CJX��e��96�_T̉-?+pW&�5�������ݥA���{������������W���}�;���~���k����z�^�p�� ~l?����'���_��/��1�*6p<qk����Q�O��P�@��<.���9Q�Ȱ�Q� �t�r)J�G�q�e?+�	����I�>!W���3C?�r�`���Ɓ �6�9��*yf��k0�e5��+�����QY7�Lt*{$�J4:`w���D�,gL�+�C�o"��aPp�QIBx�����2��2��15V���4v������nju���P���2�e���o���هp�Gj0:�LLV�t���+��\o��*JQ��Z�	!=^�R9���ƖGr��'��J'@=Kt��� ����e�l��8U=
����śj�����<�ѣ�˔�D#i�;3���n~���q�H�g8֨�]F�F @�rR0����
<M��G��!c��kz���'b| "b��|16{5�9�v+ T�"�9��.7<����j�x&��ؿq������k�� ��rM������D�1�Ads`F)�瑩lߦN^ '֐��h�{�-�H삅d �Ko i����������7w `��#G_y�&#���v�k^Wkl���4dЀD�;�t�}�l�mS�.":*���D���� mW����Wv��(�L�A�t�S9lCs��M�?��+	��#]�H��
H��Q5q,}]쌶5ŏNOu؀\cB���O����3����8Ȭt:����R8y��V]�g��5����K�h�tޠE�o!C@[k<-4�愛2�� �g�/}5+l^4:c��Bh�]l�i1UF3`��+� �P35u�\<��2�� �Ց`��v���ȃ�r;� ���3�v��;��7��y5�����aAȨ�j*\���r�6���J)�1�[:�V�C�tj\�8� �rg�Կp!h�SB>�J��t�i�49po�{͵�������$}G3��ƅI:3溺�H' 1F c I��J�td������h�#Ē��E��RYc�f� �ў���ߙ�JE��n�!���� +s�(Q,�y��p6����
��|�aWt�W���]Gu �ܯ&MC8*c!2�<�M �Q)%��4�L���ZE:����Pni�(A[�L�kF�D6��G<u��"�6Bgпu٬���]ŵ��t.D��溮7Q����	� �?���wvj�6���&�Dۙ�N�N�H�Ȥ����
Q�u���=��3��?Ϩ�˫	�qvی6|��*�#��<i�<�����H�8���W%�Iԧ�?.w�_8�r�����0��W'ZJ�
t1T��k2��y �u2P�Z��;� �D�iѡkQ����L/[�%�(���hH��s�r�e�<��(�AX5�-s��`3Е�}�؂K2�� l1Nt
��9%ٸ��dQ�\��BI��hHp��D�v�-�G�KF���n��b$�M(��@��d���D��UYH�A��?u/x�5�z�� ���R�<8L��ڶH��	J��$���1�l����J�W&�3J[$Tҡ�Ib���l��#;y��$t�Q`��d'!���ԗ��^ESZ!���x��M��a`���;=n@������>uK"_�k|��};��@������cڧ���X���h2a'��v'ܐ����~����
�ʷ���,��Br�D��f�PGM~yLbZ=�~�WdWwx\���|���m>�&L�1tEnM��O]��WӪɂ�����fQΩ�e���[�W��O0����I!��,G��7�C��|�Vޘ|4ul��m6r��9�jjW8��؏S�4d��?�\bcl#j'��${�x�y��6%1��F%�\'Au&�������l�X��9�:Dɓ;4� vp�����I�8�:�ڻ$�]�7b�t矸Hy��|�H�n��c{R�m��\(�p��!��rrV�{�H���ƅl�&Q���b�dז�=?䋴����Oy�}5tĆ	�Y��y͝I�+�
E�����#����2G`��h��m�#b��>#?-��n����,(���D�N�S;}߂�'��.���h�21wj���!~<���l�-`د��@J��.;��ܻ�XbEi@���Z<<�_�m�v�<��/�Z����ۦ�y�pb������F���9��]�6������c%6t�'��%�#��J"+�;p3��6j�	ldS2�J�Z�u[Gi>�����^Gܶ����\���$j���M� Ǡ*u�IZ1��:�����6�� �N6�\�ζ�C	�aՊ���w�d?~���h���1q�r�����<j�k�)��sk3{����:������?�x�'�vx26�7���&:"�g�ј��k�!��~'�+�v�6��ƣ�L�e�<�c�#y�L�
穉c�&uR������.�oY���'�����G���������/�ۿmo�g�����z�^�������' l?����?�~�ٻw�ܝ��c��U◻�b�`S�^gU����w��x�2����Y$x��+\���Ʃ��]�Ш^�_��*׹���M���Ymr���g����?�aX���6�� ���Exi��m͖�Q牺�!�p�1����o=�9'�~��m�� �#�Mp|����e���a|��b0lQ�3��f);���ñ\I� �I�"�F����Bs��[��6��uh�@�\[�ަ���5�;-ދ� ? ���-΃j����)��yM���� ^��Ā�R�9V*�h���u���eno0|u~&`r����]T�l��<+ΝF�d,�X���U�$醙��p�f��V0r2��Ǵ��"`=���1c�mWoˈ}��}6x>�J��U{��dtsj�l1U�|$��h�b�E;3L!�t֪��'1����T��!�����;-�9��r>�D�y
���4	�3�H��+���V��`p#�b�c�d$�A�C<K�&�H��k�[p��Zޤ�)k�*KҔ�¾	�@���Wxļ��h!�+A��^�
�M&�tz23�9�oH��؟��li�č�%�ژ�0)6ʪ�G���qy��ؙ���8�I 1���;Hk? ���A��d��b��I'~oF��bm�U�P�~hy6-��/��L�(m�=d��8 /b{M��aL�N�	RJ3R0�q�2�ʔ�n~N���S����"�c���؋ Id|@�) <�/�\�fr�f�\�~��@e4C�f]�M�baCռB����3Z�G��Ev[�g�y�#A)�T�m��5�՝��
^��L�䓐q����}B����6U��*�F�rs������[Ns�NE_,��(h�v���n���f�Q�@��~�`���0��p&3��A(Ƀ�[?��(���Y�}2 �cp'R/V��P` �FOJ`7�ܧA�b4�1���  �D�G'���6�س�WC�A�����)n�4���4�߽���~�i����d��fg`�+��َnS11��>j��(�8������
��<��O�'� \��u�e���G�Lk����P�������Oje���\z�f������$����t�����t�V�:ٌ`��W2s%�4����O���A�l���1&hm��.0���ѣ���`�z�07����S���' 5}gr�SCv�j�8A}[���Wҹ��K���L�4�:" �Lbj���O�T)����7���]
��cN�
��(t�Ԍ�
Y{n@�E%>a8p���m0<H5��^k�$C������ּ��'�,��D�e����ν-��GIV��2ڼ����	䁅Ѷx�`o(i3_ˆ���|��EK���@�`�8lh�=��oWKq&�C��˝Uɴ�eW��M@�?r��G��n��[�a��L�~�����c?�.��QԺ�/4�!N�k4[Ӣ|=B�>���;� �E����&�1�����J���R%�t�[6���ڛC3�Ni�.�쩍|�q� �3���UФ��eGw���B�Wf��p�J���6�Zӵg�]>�d8L�&��ͺnz�5A����հ���uZ��	������߶��0&`2P����{���WO|b���};�P�v�1gT®�_p���&b5�(L ��]�]���}�3y�Jw�䷝���G���v��Vٙأ~��Ԛ8� #��� h�6��!�)� -�}�
�ֺKF�-�jL,�0ʿN����+a�10�KN�o�m�u��G�����K�o���Yڵ�dp�O�~���|�ke�0�"{�Aav�˫lX�M�/A����c5��Uh嶃h���6x��L=��p�O�]�C;�����Й�a����?$+�V�����D��ɕ�)Ֆ�� o-��2Ig��6�y�L�xsJ�t�=l욧�[�w�
��^=�v�.?�f*����L�&;M,}��S~4&O�����]�3�Y�U�Y: �Uxx�LA��`�lK�����f��o�t>]v�����O?�97���&m�>��D�x�9��v�l���>1�LO�u���"��C��"~�D����A�M�S��?3���nt�A-E�:�ev!���{e'����*����!
�c�!Hn�K��7١�#X�U.<r�#:7�x�����:b#~9Gڷ�b.����}����Ԝ��8��$�5���n~��3��쀎����\bV�4��؃���r��Ĝ��Օ��А�*��}��B�FZ����>��.�um����7$��L�ݍ��Χףų�'uJb#�ec�m���a��p��곝��8��� 3�>yLA�k�ؕ:lums��Lx� �����a:�t�C'���&���g\�A[����8��D��ꡣWY�h�5a�:n���d�l��St��]��5�����	xG{�ޛ��_�v��÷��?�⋟����>ٿڷ�>��^����z����E' ������a|�O��|��w;��� ՞���@�H�1� ����|/���Ӊ\��@��a�y�*X�/ ��Z���J{C*9?ώ �
�_:��4�g�N`��i�	�\�d?�>��z d�����nQ�cWE���l1����bx���d ��8M�9�"3C�5=���P���#��}�p�2<�F��"��D��<@%
�x�hcm�֖[k�fMȔ��9<�Ũ�\}J
��;�K�����J�`���� L 
� �����3<{1� ��1��#�=5���BC���M��]Q��/�I��ZM	lh�B_f����6�j2��[�3+�aDX}G-n�����2cծ<�q*J���d0� �n�<��Ɲ��r����D���S�F`��8��_�n��Cъ{8>׺�-�|��1�Dq�n��ӳ�Q�-��q��9��H8
>�&�<B�X2C�e�`hS�4�?�ѸW�S�������l��C�&�p�
��=OrݎC��`� p�'���|�^N�7�v��F0�(�B*)��a����Ǟ;c-����B�B��*��b�m>>SNz?�q�<�,�;	�e �dpA�g�#:��]�D��������R#.��p	Y�=��d6���@� �;���챶ZԹ����\/⼙	Ma��)ᘮ�g;�& gcH^�<��cu�/@f�����1�dŞ �xd�!/��^���;AB����`=��:,��fU���5��ü2{���*�� ��F�Ƨ�q�c��L��^T�ʔ�ON2�����ȟ�l1y6��)�����g0��͐�i�.��j�/Z�	�����SJ�4�V꣐��Ȑq?���:+��L=�Ąⳅ4�)#�&�w6�Ă�.�)a�d `}��~�m����|kfH�蜷���'y��-@e�&Q��o� pF> �6�7��_~��~:a�ւ�)e+`#{��6��IR! �il�ҢM���ln付}Ш&ЋA9o5N���uә���;�ؓ��7zS�*��(褟uO��E��8�v��A�і�J�0G�K�߯��^AR����'b)7�<Zl��1C@�4����, ��Z�BciL��|�ɝ-Ѹ�hhI�(H�8Z�A0=g����d,�o�����?��t�����*V�,�o&��]�l�*�oH���q6���]r��"�kGpHv��i���,{�e�ϩ��!w?�WIE:JM��M��Oy(����,�r�;��m�3Mm�U���V���6�e;�����Y��*�:YO-Y�!`X���UWa��5�b׫���e��g���x�N�ȗ��>g����<��h=!��b<�+R�4�uu߹w�.���.�	�sUu���l�^xI��6]�{��u�%�#�O6��dї]��G��2I:�v׺��w��� 8L�,�zrGX��v-�g�S�j�k�=�ָ��G'�2x�^�"��m��X��) �l�t�d�?kg���J�&o1[E�'Ҷ��SG�dV 0v��U����oB��ݐ���$]}M�}[�n��į�vix���#�/<���.�:��kbL��O�	��ǻ��䲃�E"�;g��U��P��s���0٣��ɝ��~N�0�l.��>H�Va��/�cB7��M��O��mg-�ۋ+�0W7�YG�Ӑ69�QH^< l���|�@#_A�A`�7�z�6��JO�&�3�?� �`�ӟ�B�h�Z<���(��`꜡o�g�<;dF��,ɖ��#����)��UGB쮙�!�vJB%�)��;��)�8�I����!Mh�rMy-�E7P�M[���ҿ�	2�6�����w�~!�'��iƿ�M��%F&��$�&퉍�����1G��|Lc�_�~�j�ւς������s_x�@�!�T�&����/��tQ�崰�Ù��[ƦcM�)qƠ�A�m�n,�]-��iO�[�)�[�tJl�t��䏵�!��[3|_�T@�η�K�\��:���5��<����Y�(DLvp
�rgs;K6���S�ɼ.[w��nsli�ӿX��N��<��={��񊱥/��ҕ�oj���PG2�z�J�w?�6�?�1#/�`��6
�����ltn�G���x��kk����/��������'7v?\�8�`���?mߙ�����՟=���˷o�¬{�^����z��E' �k��������'�~�w��?ܮ��u���gҡ@�.�˳Gb�H�?��M�~�o5�vc"���&�5h�֎&Z�� &�C6�	
���������C����Go�r& �d�Ռ �׏�k�=���U<�=4�g��U�@a3�������*�����µ�  �l��FZ:�m�1
�G�ă�_�s�����Y���La���*�:�;�~��'�8D`�4H#0��l�/L��� M�oP��>I�-\��41�O^�ܮ�!���r���x���Xjե�Sh��30�yX�S����
rg`2i�k�[X+��`�>/ʡ�z
x���s⋲|��ҰZfyȓ��W�x�jtȊc�� l5w�J��#��A���g�	P*�lƃґ�t��G����i�I�b�7V!�`Ab����K��9
<o
J�O�:7�s�5g1�d�(q���ȍ��E ώ��od�a�Z�1%��_�0�����,��~͵���5�*g�
��؎�r\�+�j;�Ŕj�g�W��3i0s��)�-�F �o�HPy��ov�x�n��*Z�;Cs<�L�/�,Y��X��>ֽe ��~R�d�^1Ui����>t7�B�D␤:ArƦ��W�N���Vch#�!�
Y��)c�|��/����{]��&XAV��q�k%>9&�b��]t6�+2g�o pX W��$�%st��&���^�Nk��Z�Ӥ4��'9�)֫��[�|ѿI����Noͥ�+�´ń�a�U6e�C2z�a��m��H����Q��p�?Ư]9���)ZA#s��U�:��ZG/A(�j�X�<8Q�7���ĹΡO�����L�j3m2�]J�8���U�E0�G�k�R	`�x_+p)�� mk'�V|�?�������tt싘f7�{5�C�	@*�쑙É�i\�%Wz�u���_Ak̺,K�����l�De~�#z�a�f��+i(V�*{n��oR�e�"�J�
��XC�p���T���Ex�Q&ii>�9�"�v�ݲ��߃����t�V;;M&7���#�noI� O�_�>�h��k�)��j	H���z��&*�� �9�q�	����S��}.C�����e��>��Ya�ⱅ\;�\j�z�q��Fy�7c�u�p�>d�F:�5�?#���2FI�Ӹ[�uUujz~��*A���2I?
���X�3�@����������*'6SG��DɄ�W�E�O��j���JoH�գf����Ԛ��r�m�c#$��oX䀋�� �r+���Zt�����A��A�'s��C2;uf����q6��=\�J�kt�>�7˞����|̱'�c�c]��5g��8�R�U�֔]��n�$���4�l��{��4�ʅ��4�A�-����'6�s?�m��F�Fyh���CvP�d�d�T���M�����[�+�?{�kڳ��ȱ�x�S�P.*yZ#��:T�Z����G� ���-����x6�ں�-?�B��3���?��fP����Y
n,���X�.`��.���&V�6ޑ_Ҿ2����ܣզ��Y��'���y���m�[򠒵�@�Sש�k��N��'H��(-+��i�F��#1��e��ևE�ʝ�[z�;m=ҏ��'9�F����۩�ֵ�ř��¢va�xع�����\��7a��%OUN�יN��ն���_������Z���qg�����so��Ԥ���[�̇ �v_l�saw��z�3�"�.��8�g���~D=7r��F�J�}(V�Y�x��^
̢3Rc�qt�Z1�=��J�Y?nv�b���<������?��~۶���}����z�^�?��E' ,��ty���G���_~�������o��?�?��a��Jn����k6�M����Ɖ��By��/峩6�[�4$	TF�%+=k������Wm\�|[B���~�n���@-�;��ex&%��j��*`�WgKqJ��Q���z6�4�i�"�?�p��~��H�',\�X>o�Ͻ �a`��,���:���r�y"���섁|e)UKF�<�c2�[��l�Ɩ�x&)[T��<�c���9��=L��h��T�]���Feҭ���W���\�+(\�	҈g�����Lz��g�����O�+��p�2��W�B���J'�+6 �������6�r�g���0�)�K:�� Nf&���� ��I������oAZ�-fV�D-�z?��IC=��-��o'��&[�)Y�v8<Q	���AC?*�f�+o*���c�Z��_J��ݚR{�l9V�T�|�!)`�<�~�E-*�%�g}�r����/������Cݻ���,����#�*��<�%���eZ~��'�r3-�]�˘��0G��IG��R�A�`���a�����6ٕ��?ɽg4�D*>��q���oӺ()��N��Ĩ��#�s=�QV��?r��hm��u�9?�3�99pX+&o�oS���KF��+ɼ9J�Y�S&��񸴽4G����4tT�V�t��1WU�s���0�!�'���9�h_��T�ۈ�$�<Ǩ�yP::4d�F�b-�l(��z�)]�z�!U��,{��)zB�f�Dq�h�V�@|� 6U���V�~N��M�88�>��S�#�t��U�'�]�qƴ L�y	>��y�W�V����ʹWi�Y@�������*�1醰]��w��k�����wŚ��7�V4l���	�~iܛ��J�K��������1ۣ�>̰��nշE�HfYG���#����d��Q�l,��0����=6/���1�"{	d>ؤ���z�9�z�u+�a]v��#}�Ɉ}�Q¡�ڡic�f5�o�'���F�U3ud�>��M��:�/��z?�'�Jk��d�oi�i��+��e�ᾣ��GmJP�����rV�K�g��?'�X��|O���{��߳l�>��~׺�;��rmEa`�6�A�ט�*��}+Vd�����b<=�e��5�(�{�H����n�r]Ud}]���(� k��]����n��[]�
^�<⥐��*�f���i�mG�2G��:��!�>�\����;h�7̽��0��/�{(h0ȰQ��x�oa=���J��r��J��x:��g�%�k�~���\�H�8�Cv��x��ԹT~�7�ˠnM�K���êLz��?�9�.I��]�Ïgԗk�H���8=�wƈD�Y�aVu�-u�����Dc����GY��3�NT�TȧėD|���H�s�Z����SI?�Ƀ��b�(��Ji+S�����D��I3Q�����EBX�5�����^�p8V&~��Nu�[�f����))��-��A��_��^�*)ݥ '�y�_�)��Q�$����������E�cz�JZ��}GEq ~O���<9wc�r��|��*����jlY�s��t��D}դ�r��}�>CZ&�?H'W��d��#���ЗS��q�1S�2�X��{�ۘ�� ���DÞ	;y��R����ow��(	Oz���0Qӱ��m%��3t�ő��=���s��U�������p:&Wq�gٱ����pϽU��0�ʽ�o�X��q�?�_����O����ڿ��߼?������P�^����z�_h�@�k�����O������������_���w�4�֧:Rz&][Z���,�r����@1��%Eu� ��x~���:[w��z���]�?����g���-W�K�U߼�ᰏ�'��^9���
ჭsΛ}7(*��9�����3o��-�k��j�lE�Xa�6ޛ��	������`�Y�i�i2�@�H�H�<�+=�G2vd���<N�N ��]aDh]8�0�@�}�5�e�a%#C�$�^��Z� wo?t�pt<g,T1�'� DR�^��U ��{�Z]A|�V
'��a��N�[�5:�t8�~����6�;H��,#S�x*,�\���{��)Y�'�= ړF_0Ɍ���C�Z�Ţ��T��R�9,��`����{@�2�#��&q@�PD�<�\���9�R�mI[�r���;E����?��r��{�%�Y��}&�
x��������V;�`��ڞ�p�N|R��l��
����[��䄅�\�]�1�9
�4��Z�co�'Y8=`�L����
����%;f�\<sx�����8P�%�{ɠ}i�<��"���C8|�	9P��lW{z�̠����Z�^x$e��6���	�c��u�H����S)��}�������l�<R���	���r%���v�fq���=��dP2���b���@�?��P�t>O:#΂=�"��bM�N�Y���[�;X��4' �/�	�L��0N�ղ'g��%�Ґ����'\/�ң���#`�*�o�OU�8�D�e}.y� �����Ct~�9�ZZ�5��l�F�R�A�"4&=`&Kc� s�������Ռ�'�'�E:+ۥ��5A,�ר����f�}"��db�l_����g�
 W�h�gZ�=��9�_�L�cp��r���WB�~'��c�l�{����˪��^P�z2�N�o���iW��U����v��IJB�5,��F��'�hs����s��Z���2��}I��O�Z���<��@߲ߏ������k����ծ)��U]��-����S��hW�/9�<p����H�xt�~H���\�Uz�"� o��M�v�G$���ks�>y���TG�=*=3��6���R�^��M*O�/�}�ߧ���V��'�U6����W�m٧
��l�_���3�v~�{z���,Ԫ6�h��o���q+�%f�'d-�(���8�߮	?�Dق=w��&�`5Q�j�Bd�Y��HHgqMp��� �|J�G�u���r �2�Rq�ՙ����Y�Y�7dlO�Y*ߊ��Uu�%��V�`T�������_]�ih�S��d���Nr_�i�c[�Z��Z��#�a_viHԭ!��O�+[��:��Y+�mq��|��o��NҵJ��-��S�8���������~r�-u�G[r���t}�E{���hŹ��ɣ+ds껪^��R�p���wi�國.;���L�8�(_��*/
S�}k�<�s}���y����cQ�?��z��-���O]�K`?���1��� OK��6�桡d���d����;$�Hni-Oj��]�Z�&�G�{�b�*�υ^�#��#�&�������MBa�=b9�&��]�ƞ3��]��$~�7J�X7='�3�g�i��?g����*��R�>n1/em�(�J���ݫ.��=Ed�Q�p����z��6���"����w��b�l�?i{���x��z�z�>�.��~�ﴎ����d��9ߵ���a|X�=�t��� O�<%fe�2���7�y����ңF��2A�z��aDN+d�nWk����_{�/��Wt��o?<�O�����N����z�^/]G �w��ݧ���o���gۛ���~ޞV����YW�u8�'A2��+���^����K�7T��4"�S���p�ۻ�xs����7����>]��>�u"��gɬL���]�'ك����<��=��n��?ؗ���?����n(�Yy�o�k�r2�ˮ8��S��@���k��`�aM��2+g��*<��L�N��[�
(��m3��r�q��4
0%c�7K�D�<-A{"�UF����3�dt�q�|�Ҷi�`4�]�N�̖I^]���N|���yx���-E�
�rk��<[�)��hCXs~e�m�|�� ��q�6�r�1}�2Ӛ���ڃ8`\�5���b�Z�4���tkv�=�k%J�㉟�}��Cb9���O��hݝV�Mwď�3����H?'y����j���I�/ֵ�V�ař:S����@���L�+���tT5V�d [s���z145:hړ.!���z������s�:����!�3� �����w3���ASse�K��<8u��	��L�9�s�6oI ߂N1:2�%�`��2;Dse�V��i�0�L���|��ۜ��e%J�X��8��������vt!��MP#�	���l���	�=�{�n3�����V�i-t�g��'9aGr�.��rf��?M�ūf:e H#�C��
<��<�騄.�v���
�2%fgb��m�5hv:�r�Jė���'m��F<z( $=�O:W�zV��N�h�n)�$�&�<ı�{��ؔG�Ҿ���,�B���ܬ���N'�-)g�Թ��f�|(}tҏJ6HI(A��`���s��[я�g���w��["�U�ƽ��ꥠ�$�c�'5�vGr$��]c�|�s��`�u��|˜��F��z�Е�Kʈ�i/t �[�L)��(d)��չ��t�M;��N'~�	�*?G�4A0|L�X׈V�Zkܧ����W���u��la�r�ޟ n��2`�E������_��x֬z<�u��l/���aa��H�~XK���spe�q��F��bs���Ё@O(@.t��CfI/�.�G�S��f�vY+��S�/���,���zo-��6�_�G���WzL�H�ݠͼ_Q݃ys�$s=�hy��-7�6�3U�^�{1)T�+|ɽ�ܮ� ���r C~�Y�~j�E��V̀L���,��5����!rX{�#��A�������w�#�E/���k8�j��z�WT�r��L�X����<E��j���^��̎���9Hg�=\���2���|+�"����?�Ї�#AX�F�j�j�?���qFa�����]�����Z����<z&�?��[b$�W!]vi�U׶�ȹ�4�XS�_'���� d��(k��d)�a�����9������6���r��u��zt=M�>�F�|.�;���v�woU}L@:GN�\�ԗG����ڒ���o0eD	�7u�O��!��3���6-�_W["��Y�"�L4�gF׋9s|��0��+2i�<o���F��HdPE�P2^K��I���e�J;�l��`��s�6�#$ұ��Ş��B��:Z�h3�PӾ�ߎǪ�3�U?��k+2�b5TTIJ�;l��3���8��K�.Uʜ���hX|��~�}m9����7*g��d;��3}!�[}����FWe[��!{�3rW�S/�_�q�=2�=�n��X��m�<*T����#Y~CI�߾�`���O���>���ߴ���>�.���}�፽�<�sY��<�!9����ƽ��
8�ϛ}���~��k���{{{���}�����������ﭵ�X�a��5��I��3	�vISG���,r�&}8�om�nO�����~�Y�|�M�MN���z�^����I ��|�������V�ǿ��6�s����� ˌG~��O`��B`����G<*Ro�A+*ĭ]�9�������~�.���퇟|�>�+����y8۬O�>�0��拓�c����):�����>��+���O����_������{�� ԥy��X�a=z�,��P��� Ԝ���u+x^��&bZN�O�!-�_�p�̊I1�����48����0��薃�qP	*#_ K5�N(^db���͙��Z��i8C���P�J&�c�j����9?�9�s�lmS��Q�xv�<��n.Sg#���8� ��<�k&]�q�^�EU�,��6�Ѥyji����o�:zɜ.Ll5T��$q����R[���
c5o��V_�O����p(������+�x��fe]�gWٷ6���Z@ ��e��A���F�y��Ϫ!��Y=��j'�� P�t��u�,����C��u�G��B�)�r8��p{�=�]3ޑk_(:娎<߭�ñ)8�vx�'�b���0��v�� 5X�{;��,�l1��?r�c|�SR�|��G���|���L�8u_u��<Ŀ� md��.�M��(O=�>Gy'�'QK�\'����H-�w:����}�ǟ1�|S��;���7�Y�㎎8@٬�ك��ؼ͂�:sj+���(�Bl[�y=Z ��N�X@G��>M� ��1���[u��ٚ@��`�<}_��R;ӗ�Ü�)��}�q� ��v�1�9�M�$�t�,�����r%n�3Ϥ9<��a��t�A�J֪�*��x��ao�i�'eB�:�?��(e<���=V�{�W���Z��6�E��>9�o�8k}r�o��YV?ӡ�KzW�L����K��.�d+O�����3Y�O��+�m6��[y��2����|Ip�9} M�T��/�m٩G��M���s�{%��c�#�U���ܞU�V�=P�;�;���&J�[���Yc(s�ў�s�糝��k���	��-���x4ǃlt�=�O-�_�V;��,v��q��d/��zw���>[Lo����^�nq��rw�_�V��+Nv��qIX�6�q������#v��Z�j7�*4V�U�����]GU�e�����v9'r֔��qx��:z���D]��~��g��W�vG�(z�veyFw���?��eM���٦��i/[���w�묿Y�=-:��fyG��������k�G�K��wx�����Kn��q�w������kϕ�i��a��+��mz>l�Y+|�{�?��~^����N�|�i��7 ��Z�d���,2d֤��f�Fc;a��f�v�Y�'i�W�Yd����We��^e�~[`?���V�f��g�;����g[>�-P���A�ASn����>IJ"�:uXR�,;�5ݥ���Bg=��e�6���G^K<�E^��SY۰���P��Y�.u�Y6��g�Y/�?בE���Dp��{��a�S�'Z���¸�k-�Ѧ>C�>t������a�8�8�?�A��7��:R����#ݟ�`����N�fR���Ϣ�xFi3%~��*���ǔ�*RXk�:`<n�e�/׫���﷽��}~}���̾��S����W$h%?��G���}�����-��wn���������=ݿ�n�?|�����/�G�����|�^.��>�E2���9Y������|PA�������y�=|��~�����3�� {H`?_����z�^/^�� f���o�~�~�g������÷�w��||{?(�����=2�%��N#c�~�2 W�r�4%���l���<�3S�z����}j�۟��?�7w����j��lۏ�`��z�sOe�I�m�"\��;���?���c�������[{��{��_ۏ���~��+�Y�������vW�c�����Hʪ�ZP�j�n�KT�A:f��)�O�<�C
]������)���ʳI"[KU��y	��4~q�"{W�ӳ΀��7;He�'д::�L�mzU��ӊ�y�L�U�Z����Sε� B�Y��Q����4_|^ϖ.c�َ?n�WHb �D���R�Az�w�{ ����Ვ��9n��L��<���>n�g��;�_>Ge�����B�lG^S��H�����6�_
/iu��8W}��x��Hy��/�S���/}�d�C3oR�l�S+�1��2��Йtz���l�u���g0rnr�%��g���J����/N#i{x��|�t�
��Ǒ��L��9�������ɏQ9nwX��6:��}�UPZ�ɳ�ٝ��ѫ{e���tht�z�,���i��)�<���?:� ����' $ְ�o�������Y��=U%�[u�Bgq�k��Y�=b$�<O:�Y��*�D��a	m�8-��%pz��$�ן©�ϖ�P1�y���1c�zg;��9ti�p��^�k����`WT�n/^Ym�c�kZ6^�U� �R&Ϲ�v�Q>f�#��c0B CP�T���CԵ���gR1>k�:�H�Hh��(�������&��OE������K\]m��im3��2��KYGUQ��#�<��ջ��բ~����]2�͑G]���̿��Zo�xZ��s9"��̨�o�j���z�7�ʊ��cN�g�'�*vC�u}��#[0�Ki���3�#�?g�<�`�-tIy���a-����)kk���O-�I�׵jQC�]6tz����<��}��J�*�"�|>v}G��w�G�{Z �E.��f�wt�I�ΘC+�,�P��tsY�:�����"�z�JTTڵ�c����7ؔ�@9��\kHn�V=��1�e�d?=�3GQ�?^Ӓ��_�w�"�x�ό��jE�� 1��GV�m*A�蜁;�O����Z� �W4I��Н�!�X}�ڡK��8��.&ߥ��n������%E#���ly�s4��PȤ�C����ӂd�8}n�[u|AԢ�tLQΥ��9V0�\��bw�o��B��a7�xE;�z��=ߞ�����9��H�:��p���WٻV�v�C5��/���&9x��0���>VA�r_�^Ҩ�[xBt�	�K�=(ۭ�]s�Ǒ�/Zl��:+Y���1�j�&�m��M}|F�'�_{A]��/���i�db��YV`��������yg
Ȝ�Ou�ƍQ�Q�=�q�_�W��,��C�і?0e}��������?��@��MZ�t:���(�ċƱ��8>爳���z1�i��PXq���OԵ�sR/N+6��H��ϣ?^�rH�z����ܪ���Y�3P�\.�}�ߔ�z~�<62���T�EZc�)�Wk�Ձy�ܯ�������.����>�_ZA��'������u�f�����7��#�;u��؋2�����;�o�g\�z�����w~�G��O�c0�y�w�������~�u�pW��!k�7H`�7r�ʻþJ�=l�j��R�[{j?o���/~�[���������/�����]��=ڿ���޲���z�^�����'������7��?�����/?|{���rW'�6y6q*w Om�ܘ�2i� w�;嬷o/Y�����{?�~�����o}�~���]����m)�n��.�g:8߾�s��c��<e2
 ���.r�7]�����ތ����|��b?�~j?��@�}a��ݗ��h�g=m����I{����y�irP�1�Bo��;�����5w�=� ��r�O�V���@�Ű/�i�����k/�Z� K5�v�9��Y�n���-��SO�ڎguWC�~�l���C�a�Y�|�����q�� ��u�n 3�8|� D@�yN'�����噾~99N�	�y�N�{���;�7ޟ�+�ƾ �@߾G^��؎s?G{)#��ҽ$�x��h4���Z�9� �Ƴ�=<Фʋ#�d���a����/^�(���.��6�(m�Mv�?����|h���ș�qՠH3������	ZUʈ�K�P�wݳ�l;��i�S�G���`����8+��9�	�X<Us蝴xav��Sk���N@�|�&��ص���43Nk4�����:��<�s��J�I��TMk����~�_���+`�� uhU��%x�z 13��}��E'�X˖�ǿ��&�&��K�����#��g���=Pm���ډ�Ǒ/��	�NKـ�(��Sf9�z����}$�[e9�%>�7̳@������L��1ܫJ`PCI�ɿ��:Z�ˣ�-m�w��rPS@�u��s&>,z2�-�z�9���r������z9x���zT�F0������c�BM{�m�CGk�u)vp��dް�*�k %�vӞ*vE�WI��[+s<[:/��V�}0u�YgkV>�G T������9�r�D��V�hϬ�0�n1�y��lG�*���ht��j��:!��f����f��}�(�^�A)[��)��:�P�G��}3u����%? {�K�o��m��-�+��5�R�򖠤������ڭy�v��Q�a���:�%�$9D�X뒮�c~�������F�ʿ[r=��X}��H������ ^]��7̤M|�ǅ�T6;���+�<ɐ��Cn(���]���|�A��q~7����o�Z��D��X���;����[�դ$���Y굦}��r�тs�++�َ7tZZJ��G���LI�9_�>��H�Z�k�@�oҍ�;$�� z������s��]p�2��,�@�a���*3�j`7�g���2]݋j`�7��T
j`�eL38��\{{��uy�v��bܬ"��kYy��=竇�d�;U.꯹g�a��A�c�K�5�vt�yrO(A�:?���f���ٻ���f�$� ���P9�Wр,x�H��x(��O�<�s����ع�}�u�CT��>�U�u����s�g��9�MqX1���p`Kޚ�V~�~���3{�؄i��^I?>l9��Ar��$q�� q�LY��r�=h�!?���W&Qi�d�������QNh\}���:H[��-L�3% d�0���B�2�[�Lλ�����ޕ��w:��{<��ɰ�������GG�����3?��6q�ۜϑI�	\3>7������`<n{s�����~�����|jo/���.~�*�T���c��:�Yv����[v1Ƀ9v�e�D+������~�������o}����/b���}�?w4��J	��u�?�B�b�G�%>�xj�;�R�o�������/����7��/�������������O�����z�^�o�~�	 K�^���������w��ǧ?�q|�����q��j��
����X2�Cth"�hS~��t�L�<�+>�?�{o�׾�=�����7��H���<�]r'��܊����ӭ.���<�f����  �Ez��g�0�$�F��tkz/vuU�Ud�E2���{��n��gq�������sN��������f��I;'fZ��Z������V׌a D�]u���3]�t�lM"hY��i�7�S_�xR'��ܿsz[ޘn�gw�ϟ�J�{��<���qeW��
�g6p�� 4#X�	f ��$���{�4P(��L�����O���R#�!��2`�_"l��z���&����]����,����Q��BI�3���3ےSC�������
f 0gP����Wi��T�.������ �o,p��pd�ǹ�4F���v�4��O)��g�����
gp��O�﹣�p��`q�1�w��!x`$��LK������V�YQ�%���S�1+�C�q��Ɖx�ݨ�LP|PP��N� YU�U0�J��B)�	1nXQH,�h��⚼�܎;vG�'맟�gm��������*���uy� �)�a�mX/�g�+�ye��h�W���iψg7���p�����w�9H_e{�9��L��{��:~Z=���A�Yz�x�����X����X����[}�N^�#����5���>�e%
&�Y|ey�[$��NS��=Ę�G�H�I6*�CJp!��2�����xd�����>��Fz�Sfg�Uӥ�0'}wEs��� t�
�˼���ɴ���V7�ZP�19d%h�^����x�U:���lu�����o$,�(e|����G�2���H�����/������:�C���0���W��� 3}>�9�R��c3�����L�s�1���s��j����A����� 8������_��U�fݝ0�x�Ӄ�����߷�}.�y�XwJ|pX3��
|�V99�7�F��	�o�M���zڼ���g
]ݵ���)q��i�����H�N��b�~r��x�n��n�k�:�s��)���'"�jr�T4�(Z���<�]���3�k����ݷ�����6M��7�S���v;-	�a|�;��_�_�����,�ì��FL�x{�xD�J�RV��m|$�Y��w�>�b|\k��y�#��<�;ƹ�<�I$t���/8�T��x	5�)ZR��{�j��R�p����}�3�9���m�����_�28/�`zg�M���Vk:����}���эt��h?��W�Zb��Bh��L,�ˏ\g��\�����=�rō��`�����y��B2'���s��^ �Iu^�M��I�]�.J~a��<G@��a�Y��Ps�t�O��ڑۅ��z\�c��,"��f�v�S��89�d{��8�q�t?MS��#l��#�W�c���e�N�Clu��㒰6�O5��$��g�g���F�	ޝ�)���V��S?#�]�1�ڽ}g���N���Uh�<�x$�P�V�dJ���)�ZH[���?�����+s�ɰQB��֭����<��2����jC�����
�������d�7��t� ,Ƒ��x1��~_=/-s�k7������+g�r�TuZN�̵�}�G�jK Xq6�"�n;���gi� h��3tb��Gl��\,�l��d!����[�_�Woܖ�}����g����� ��#>����R�2����Z�.j]N94����ig�O�g�7��=����?���������w�o���X��\up�\_���u}���� �s�y�l�<�����|x������aZX�3���ƀ}�g�N�`0� +K'�-�k_e���rnB`:N���������,�>I���u�u8o����"l61�9�վ���ZB���;m\�uyz)�F�ڊ����@�sUJ��\,%K�ޚ��kn�k���O}$�����5!�ZVWMI�z;���ک/�����ʑ9DV�{$GGn���  ��IDATu����[��iFk��r�)y=CV�� �U~��U�W?�;��d  ��ӱ�8r�jCJ�+��6$V6�Qg��mmw���]jw`��~����5�79k���l����vb��g%*`������Fl�k�'E��	��s[u%Ќ�ٔlv��66:�����Q�v���V��3ӆ|G2�8{�����`�-V]�Q;��k�u�w�T�q���o�VJ�w]��.O*���3ѱPRNhN�6s!)�ʣ�c��V���e������K���XZ��Vj0z�`V�*�C2�r�����Ū�0�b+M3�h�h�F�xt���+���N�Ƴ=8�[�[e�.zȫ�w�[��>�sٰ��F�k�1�`�� �����������,vN�8\���������ev4��G0l��NN������,A/�X�Oi��{��1TCQ8я��S���_�I��L,��;	w��,z	���?ϩA"9�f��oT��~��Lwd����΀6����Ϭڲ��y�/�t�yr$����+,+��P��"9,��6iC������h����V���sTKbT����@+����?8������@'e�v
�F��ӧ"��Y�T�i��h�,�p�V�~�z/�o�L�)�����iϏ��$N�<?Q�����9TqG����N��"Y����'>7��p�c�L(� ļt~��5�x�\���������k⣏�iS��X�Ͷp��N*�_���Ec-:SA���+y��ߓ�+z�Yռѭ���S���~/vn�Ni���������)V�4_�N�H�t�޶�/�P]�Xm��Dܞ�z�u�h\�!.v�-1�.x(�Mk�_�Jq�a�<���|\\��ܑp�>��	s�qTC6�6;� ��(2������<�]���tQ
R��{���q"��,q�M�Sҁc��ϬB���0�A�*���"�=W��4���?�%�!@�?�r��J�(�t�x�12
��Lia�KO�
^�����7I��%�z)����2�*x;㝿��H:(s�$gdZ@��X�>���^� B�����<����愉�?lk�z'5�V���p��S�?�1�CbNV����;��c}2c�6���I%ԧMU�A����P�d��c&V�x�*�䠏X/$����9x��;=�g���ݪ,i���3�hL�H��Z��!�]ή���ݣ �	���h�}��x��Ok��#pP�?ٸ`E����V#x�Ԑ��w���y��%J�T�ݸ_�R���y�%��cНy�D"<�-�B����;] 1,���jƟS��54��1n�GgI�[�=�/;@	�\�<=qK���>���G��gl�^*�e�N}��F�I�`W֮#-�=P��y�7��DgVk�ˮk���,�.A">g%�/
��cu$t�]�N������P3�k*���<;<��~������oG+����o��Tڎ<���퟼2��Dz��/�䁘;��| �n�곟/7����6�lچ=<e}׻��06�s.��tn�MV��8������ś�E,2�NU'UN�o�I�B�U�t7���R�ޱ�'7�;/����=�
p�̗ns���<?J�g���}:ORWĜzQ��+|����{4w���v�%���[�w�G�B޻�T>>�K��}��_���;<-y؃�EW�b���j�xy�xy<p����}r��d:�}~���\ʭO���ܓ���������/=�|X�'��O��dzV.�Z��y)h�)x�Z������d���p��r�e�v����_�.���(��~��¤����*h�nl��{�cP^���f<Xi;���7O\�!�6�֭�}�{Ӛ��=��rk���{�������'��㳩�H�"~ݩ`��X¸�%�H�
�|4:X	`��{]r�vz�yW�I�mꦾ0b	��b8��26�vS(�ti���u�s������cĆN�S>׈�ab�>d�V2��7Q6��V�fɉ��/��)�kI�DYbZ�� ����d��U��Ŵ��M�|�P��F��L^!�[d\�rR�7g��ɸL���)����6I�O߂y���름Rl~So'd�/h7`�m�<c<����8'�����Nt3���0����ĎR�!^EFP��	
}+8�}�����C,A�jӱ�q���}�9Q}����tT���W�V̨�!r��G}%A$D	�ߛ�Vm�^�����o%	�]߀���ln�Mr	�E[#�p������8Pw83���0O�u3�:Խ-�v���5._j�)�J��1��<ʝt\A�$�W�4.Y�#���o�g�S+@���q$����C����w�E�R�7�nx#J��H<���,������6ƖW�����&��|� �lk�Q󙙐��y�W�@!;�����tg��<�0n��(#�Bx�Gh|��&NS��@�4�����A���{Yb�_b���=�L�͡4��XYp!��5�X�b�c�(�ƴA��7�e�����6!���)vm�L��cK<�����!��.���3�{� ��u�uZd^9�8j�K|��1���A��
������V�+{�ٛ���hN��ׇA2���$Z����l���
������]J���d�60|a�b��h�^����K�ƻN�d�`�m��U��Yd;t�?���v�B ��d�h򒹥Ӎ�� =0*��-�x�X���H�!�0�������({�9����n��+_��R�A���d���HHtbMA�~g�@�FOϴ�j�)�6u���bw	�9a*���L��d�﮳�<�3�NI}>�Hw��^��_�׶}`�T��ȟ�w��8��r���@�`�t�C��`M��7G۔�[|Й��)�vx��SKpH4���|\|Vo/E�z��Bp��]�����=�Û� ��s�x�&�<䊫۷���e���w�d�A�����G�y�R�^	��Z�E�Λ���S,�qy���qh]��
�dxǑ��&��/8�5�l�����I>��P
&좚vbk��Y�����W����愋���&�q)���P6���]5�Ŝ��D��n��� �I�Rf��Y2�G}3���o��o|��]�\�-�qG��aG�PDx�+�?�j�y�`��H��}'Y�"����!�{_#�抌~�,�r�]�M����2��S��|�׉	ب�:�m�[�'�;�����FiKG���i�9��������Wnޑ��M�[��Zw���؎� ����0��2�;N:�9�/|��v�c$�L������;/ɍ�r��_ȟ|�||2�c��x��Q��ɱa㲮��6��+�^^^�.+�'R�]�٭z��l)yQ������u}�mח� ���ù��O/��'��gr�\�u�U_N�<s���Օ4��2��0��O�| �����=y��W��ٍE��ph,v��p��XݎV<�T�	o�g�Y�U�Q6tU�\�0���2�m����{��Y�c����׾./?�H���ˣ3�'�J�������>6�u�$Fb��3ά{�eTBYg�"� H8gS�b�q�g�	��
(�y�# ���P 8ٙpTe|�8l�Nʖ9�P�d�����hr���59 �~��LJLxrA2:ҕ��M��J^
(����ط :K�KI�r�{�?����%>�k��y�b�mu�b6Hd��/cq%����UZ��j�Te/��:��Nw|��s���D�pZ���2�VgCq#)#���p��g��L%�G��hp�__8t��&��� �厄�&触 �H���83r�)ۚ�hv�(;��K�pz�kg#�;���aИx��~o���|���J��dА��e��n�;9h���\HC���p��A_/C��Kc���	C�]V w�yǀ��;W��S����e��ޕ�^�/�=?���o�X/��@�:��n9�R�"�����覷���9_��U�2��ko`x����|'�J�%���<J���>��hU; εd�x/[\%��7v�ԕ��sv��\� C��\W��3N�m��S{(��Or�[�O��]ݩ�����8�����2��Q	Gf%�μ$���������q�-��䰋|�K�Y��Т���Y��rgW�xm
>_-����<��IƩ{cNn��W?��r #k0�:��`ׄ1��A}1����wp��V�Qu9A^��u?H���﨡�v\	�Uwpu��j[�J�r��hBfTy�������&KCn�(f�^�&.K��^�YNB5ɨHԍ>oh���x�7w���W����p"s$c�,��&�}��L�h�����U��u]M9چF�V/h|cKP��eY r�zԭj&l�t7��:��#����� �G$�k�o^c>^}e;�?�Y�x���F�ſ '�W��_mG��������L}}���I+�1�*j��²�߷�sc���5�r}�]�[W����e��h��֡��&z�d���3�=�ߨG��*�]�v�Jݔ 5mIX�q��s�װ�^U,��wp�ڲ�w�`{0�I��V_���ێ�'��d���M�)��'�*�r~k���>h�8���b	�;����� !.�mTڅ���*[:��QAj#m��5lg�Y��H�щ���yo쨴���k�"*x�2��,��1����ζo�{UBs
��I:�*#_�6p��Ѭ�z\���N�Un.����y顼u��+'rr�u�uG5�u�.�f��}6�M>(�Q�^�#0
�	��5���=h?>`����T����r��M����Z>X�`*��N>>�i�w�ěj�O�yv��-��9<�z������W.���==��3�V��������/;`�i�����~�����_�������/�|zйLE����d��+���w\��6�1��Ò'K��"�躚��|oe�K�����5Sj��1w'�)7]W�j���5�,3;�!R%:?�~�↡�m%ٳkOW�?�
�u�A��~��|�t�I�O�;�j����WQR*�
���©+O[C�U�ylEyUi�g��%Cwh7F�L.2�����#Y!*R\�Qh吒���׽��N���%a��?�5*M^�@�F�}eR�ǝ��0��g��S��n�8с~�DV����m6(m뷙�Y�O�l�p������ؤ�j��8!�Ze<�3�q���tf8�nźZS̉��a��"�૝���qM��8]�W����v��,,a�m�s����r����sV�{���S�goo,R{��(>�����<(16$��p:��Jm�ޒo�����o�3M�����t;f�����]���D�b<���&�bܷ�&8w���B����kd��7b���+0����SCӂ���@ػ�գW)���me�x~eY4�q��S
?�}�LC��g�N�FC���H����bg.�3m6R�1�bW��N���&8дy#��!c#K�ܶe��0�3��ߣ�+���t�Ӟ;��O4&c{�e�&x%�`{M��Uف�9�:]����'�I�Nz��z��4�F�����MA(ן�?��1O�~������ۼ焢wϕ�1�瘇��h&H^��G4��1���(�q��D�]�d/'��:��Z�:h��y���Jq�__�>m�M:5�g���Ne���6�}�d&ݔ�q���$��ڬ"�F�e�3�8q�Eu�)��Fo�e��.TI� �mq#}4N��6xs`lt�R?�Ćd3J��g^��]�=�{ŘՀ)kL�ؓCk^�QX�+d�h�ôѣ|�ɡ>������x�vl�, �b���u9=��l�p��>��2t:�-�}�z��!��?0}`u ����i}��"o��gD~c l����Gr7��8y���<�a���>Ž�5l�-��v��ӄ��(Ýa���#y��������PG��YǤ�W"��y=�r���u� ��ҘS �}s�d����p_���5�y�� �Λp��i���xG}[�{n�3N';ry�N,�!���:A7�-�J�c=A����!�[�4�����з��Y��]W�����I;!�z	��h,�䷜�o�=�yb(&�GX����u~AP����{��ng>���I��_�S��qn�>�p�.Z���\�L���
���e8'��������H�� k��꒞G��w��s��x��~�Ĺ�@w�8q@���lm��1(v�����^wa؈7e���< �K$bm�$�����]�g�6���Z,�8˭�ȃé|������{r��XN;2d����s=��9'�����	�A�q/>j�;�a��/���<�WmG
4�H��v�b�a)3��t'y��=9��;��T���D>[eߪ��L��N,m6�M�_�;إ �nM�$7�������������Ne�x��O�"�����������}$ oݺ������ON����������3�(�����.1�+0C�6�X���w�ܿ��}��K��+oȝE`�=�>��j�p&���k�dFC$�{dB�X��6�*�-8f��T�]]Ymg�hkm�=�O��S��K�������~"s���GRƫmUH�P'U�U���mU���
�����ɶ�S���C����"z>���je�+>$�]UJJ+QJ�8���K�j�J]R��[��.ֶ��I�FCv��hR�;��gŋp5��50�U[]Q���JhW@����@�p�(;BC���ޞ����78�����@JdB�����1��A�%�z`"��c��GE�A�[�I��%v�����cE�1���{����!�_Ǯ�:;�J8���ͷ�n8W��9ȉQa��5�$ӠsX���T�U��]b:|�f"���$���:���{҆7�w:�t�v@>%�ɠ��=�s_�hX�����c7�Q!Wg��5PkE�#b��8�qp�"O�yQ5��K4sP�xJ%hK�t8� �xe�ƶ���2��2�7z��x¤��/�ɩc�1J���a���bW^@���@ y�����xF�G|0�����i�m?Qw��+�c����nݣ���)pE4�iV�	�#�5 *WUG�2�P���q�$݂�^�08�Yo�pr9RB�A�b[y�s�}��L������}f<���'Y:�hS����s�`H" �����l�U@ z5|E���63}v����X���Z3�`���T
�Qbs������GMߝ���n�Ї"X�D�޵
�ނ��?��6{�hεN+2����a��g�2�C$L�s�����|g�1���|>�f6����vq��Gy2�WM�v�F<��p��0��,�)���\٢~B���]I�D�5�m��l��9;�#p$^K�����f�V@�l��0G�Bs��Nm�N�f��xsi��c�m�|1įɝ\��0�a�sqin�I{��(i���ss&��횏�9�9]J��m���Y�_��f)x�`߱l)R$G���j�MݔP�Q��������LnoW��/Si����z[ݼ��UG�&2�����a.$8�`Q2�]M�g9=:�j9��Խ��̼r�K����M�r�lԱ��A_�� S�.�Az7�7��w�ChU'���l�z�|$��+Ղb?�Ǒ�w/�׷ܯdWu!G�'ʌ����y�}hgS�wR���d����[��1�F80�P�t�G��+�wm/4992@�������L��_u��*>G�M�<���{&�%�6���� a?����Xx��yQ�ŕv|�O��b��$H ���l1�;������M��q�^K��y����ۋ��gN��ATj�o0�o9��c�P�u�<������W�#^�3�~t�5��J8�֫6��-f,���:�������2����q����w`�۱�}.�����}D��c1���ӠWl�z��]�i�X
���w�)g��4���R���ޒ�_���O�g�����*�h'�2�5���m����h0LrX>O�.���/>{x��O��������K�������z���& �H���ٳ�'r�G�y�;�~��;?��W���^�J=�� ��Z*��I@A��A�>[�T:�ng�,���z���U���C���ì]A�δ�ق�&���Y��J�ʝ���ː&H��zu��w�֌DY����3����Z��n#�/�����-���Ԝ8���s
&vت��]���ū�Fe8gg�U9��#�\�`zmk�y��J�O�]"&�!}%�R�{ ���X3d�\M��a�0@�#��$kW��F!W�Aș�A�QÃ�:;E�<f�� �=����Ai�++x���`r�s�0��
�
Y'n�S���޷������
�h�ԑn[�	&6��_�z�B
l�ߑ�?������Վ��dx�S�K�BC	��I-G�T�z��ٔf7 ��`��⃜��"���υ���Ʈ^��)��֖���w�W	�9Ð����<��W�m6r�Omg��Ў�� -��(4C��4!F��|O������B3�ui�M��aH�c��]�8ه �pV3'���8Z�s�={��g/�`�Z�7�a��Vwo2��c3�c������J�;���PN5�ͼ<��j����A.�|�;kp�J�Yf�U1�<� ����h8��Ğ�x��(ds�	$�a�=�f�ʅ](i:)�O� <�
`��,����9Z��c�7��mW��CD�	�B�bvbd��0bO�߻ޗ�buȷ-2��;�d��@;:�����k1�-��i����2����i!ݾҘp����A?sY-�/�ܖ�?�F��_�����d�vU�5Qv�ZH�8&!�(���ڇ2$TY���*5V�$�%���I^��y���j��|�1	`�W�k0�V�{�se�v�	e�#��ܑ��f�2���وT8�W(��~s�]�d� ��;.cj�	 i����f|�p��5�g&��Cާ�������������������K��A� 2�I.in? ��#?#9(ƪZ�5���a���O���i���c1�ܹ�v���;����?R�h?!���m�L�D��s�|/�3�g���I�n)o	�>��v� ��k|[�t�n���o���lʑ��[MZ��h^�H�"!�*X���ߓ������D��TC��H����nA�l��D�K4���g�C�.�-8�}�����D�p#톰C�.�%�K��e�~}�ʸmx?']Řl�w��$�60Ω x��D�� ���]<�nK�B��K6I���7b�����$��3�uw��8��:����-�f�l��ܖ1!Ds�&^�d���h�c������k�=:�e|䄆������W ��qۄH���w�����k�^f�x3��W|,�]Y�����xȥ����8e���(�o�p�PM��p:��E�k�_8 8ҩ))��{5��>��Y��an�|lzr�~̙��ΐ� ����N���vdY&�����kz*���������'ҖE����{������W���;����Go7�iv�[��ƻ���˻YcxŶ���L�� z��ә��շ�~�y��g�4�S+ti:�a��C�2�b�+��2~��NR���wz��7���S�~1���Rd=�(���u}]_/��� ֫>����}��G��O߿�7dQ�.�v���[���@��ו�U~/�ta�7�2��}E���������������YG�s�Ӝ����X������!p���Wkg������*i�g�([��* �ɉ\.�ޜ�|��+2=��_�D.N:^V��N&E
eZ[�`�$T�A�y�J
n�(���Y����%w�B����f'��`�s��l����s��SB:w1i�]I�:b�L
�M���< �Z\IL[�{J��+��Ѡ6lu�d�@�g �37��8���AM��,[R�4�Q��	L�����)�J��{������Ш�l��9�����2UL}w����=e�B�����Q��� �y�|c�K��^'�^�;����:����\F��Zl[<��H�)�g�3V���O�4�2e�/�=5�Lop±p��+F�Z��g���C�F��|�mg�/�Ĕ|�0���4>�1��v�!��E���(�18r
9"z�qdCuy�ϔƨ�y�p����4m�h�U.�V o@/>T�'�] )p
��>=�x���f�P���� ��@��[�z�as	3'(��Wv��E��5g�:�J#x����d*���+�K��P,(m{�;���L�ᗂb��u���r}���� �����O�_��Eu��VGy;ԋ���`�g\�z�ҷ%�!�!�AD?>�@�D���,4~8k�
��؎��~r8�{�s� ��=��ZrnoC%vY��j3�z3��D���g$�U�ߜ�$G8�"p���~��A��H`�_�K	fo�z(�����iK�/+�p�9<����bU���p.���9�}��"�s�D��#�j��W���������
�Ж`��ۛ#���Ӌ�; j�a�p��$�t�%��q[���Oo���9V,	.��us��VAձ�E�:!Q_�1�Ώ�]f��d��@�5�x7�P�G����=�P��W����5#Ѐ��\�[��>n�R�&�'��� x	�8���ۿYy�;yf�ˑ��Agdw?�zL���3�ʎr��1�JG4��⊪3�j��=�9`��Ua�#�����df��"v��σ�ґo/��e�a�V�'��\a����c�歯�b��^b](���e��\\NI>̹Z��� A�<ߩnq�K���.V�I�7Qo�����#I%Ӛ&�6h��n���R}|!c<�8��5�0�A>�>5������ih����vy��� �6g�4O��M�`���R�q=������r���G@�v���� �8�H��������n�WI�z9,�D�l���|x�?�SĀ��	_���0��}��k��T�̋���e�L�bk|������ ��y��GA
������S2��5�	�	����d\d^dSi+�g�Pd#�s�o�U�S*��r�n���}`��잏�AJzi�L�!o6�{�BÃ?�N}^��Yo�Tڶ�Gq��"����G�����#E֭�o,t�J��7���<8�%�k��aY�{�a߆f=�lF��h?�K,@��>� ���1���f���E���-�9N���+=�É�.8yU��o~]������_���s�~�El�щ&�J#���c�\���˽�˘=���Z�e��������k���H ��O�O/����_��7>�G�??>>L��t�[��&6�����+=[�� O���U������_������2���Q� ʙ�Օ-5G�oA�m�MqYb�{
�.��� � S�6��!�M�̍���O���'�(�Rv�e'����QN�"߽�|���|��Cy|X�8�����Y���*�u�Xi�+?�>;(�p��F�¡k�����#hG	e����Z��g�Kzg��P��Id���v\�n��
֢�x���v�l�q�Z-�V��`T�T�Pvs�f�Ѹ�[�'8���6Y�t�7�O��r�T;4�:8���&Ǫ(���R�b�:��!J?�w�n&w֤@q�[��k
mIƤ�8q҉>��?8n��u�"93�1��BF����U&pIƅ{���v�)���Dy�oo�l��v�T��f���8s�ۮ�������y~F�;�~��@�&�d�>�b���@�.U7��;�:o���a��-����lD�z$��1��Cǌ���fd��4���pFL��1���E�nV��0�4���;�c�ޟx	� �E��$s��@]�"p��~�WXr��q��4�GF"Nu��#�2Ȫ�\�,��r}碛8S=�`����uqPB��`�ݍL>�\��q<R��k�'t4�C_UW�x,}<��k�#ʴL�
vOx���T�a�[C���q�p`Q]~Q;�L�E ��u��CDқ-��BT���	�c����	�4�|T:T�c.����{��g��D�~7v�aG�����,ױ7�/����vA�2Ȩ����)識�zݣ�+�m��Lۚ�8���o�1"��_�)�E��.��y��vI��H��L�8�-a��;�Y��&��cG뺥fWw樋�������W��a� �-��_J�R5>̰,����Jc�"z�f;rI��h؍����T,!�h�3(�]�J-�E Ґ�]��,���X���m%��}��q12�k�ґK��k��c��aڡ��s��J�t �X���1�� ���׊��%��o�y�dOA�lcd='�`������I^L[��U�\%)�û��<g��5?g�`~�oF�2l�6`]�L���:~���P ��?A"����SO {1_)���)� *��_s��3%��
8X�*u�Q��=֎�c y�db�}L���N_��ĺL�jP��#.
w��ȗ�g�w������/��{m��4�,�t'�
�^	ߚƼ��p0_�mó�U�cI���7���ˤM�\!�{�������t
Z%ZQ�5�o_�n�]st��[\�D�GżJ�v�7�1�oG(��U1�8�:����G���ಀ�pS<�����5n��B�0Q�Ȧ��8(��3��C�(i��N>��'�Ug�ۈ�v\��S��>���y��8D���i�o��J�Q��w�I)��<�^���,\�����!o���Xؽ�[pB�&ix��s(���S�G���ǣ%�;}C��������j���Ď왵۳+}�Hh��b��"+�o�<MXR�
C?�p"tc�y��K�w�]!�E�����sjsxZ�����x��D~�kߖ��/�X~u�`[@c�=�S��%�-!~Tc:1��B�I����4-�����b:==�Yw}]_�����/5����rqrq������������?����ry(���}�+�ƌI�Z�%t�]F'ˋ��8��|��]��_��V�.z���UXh�.�N�le�	�#99�	�|V(Ek����iX1�[ߘå�Ԟ���3Դ"�,�����W!�ny3_���r�ޒ��=���/������҄�̊1��Q�6��'dS.�'e���V�	X����a/��̠��muV!�.+m�x�@$	�(9W�������F���6`S�e�eVS������ʌAa}��.98,�����3�uQw��	���#��v�Eqč{$�t<�+U�;��Y7M�QBg�ŵ��+�NǱ���p�����{��I�c�N�����;�,���پ�S���c��dӳ�AK	]�s��3��u���j~/�a�Eb+e3������X8W��-�����r�Ì 
Bl���tGx �5p�d$�uð���q�7��� 7Cǜ�/�C�u�^ᘌ�jȀEVS�A2��h�J�]�l�A ��Sp�����$<X���39_����C��N��?S�;КCi�b����Ư��V[�R���3�O#�5��*����f�i�F���r	?�r#���D�+��H�e���c�N�:� VH`U��
��͵���C��9p�+��o�� U�ZC�'���k�t���0�^h���P�;��fA������j5��s�7d�Z�xC�Х]�����A����� ���جj����C G��,�$+��Mn��i������ڢ���C/Pɺqr��,�6��-jcQ���@�����Q79��*��T�jC�W�'���fX"�h�ٗ�2�;��J���c��;;'w�F�X��?M�����%�����vā'FJzާ�~�2��y���ی�?#�����A�b㜂|Җ8���U�����;t�-.g����#Ҟ�}���#RM��y!�LF�h�G�l�s�m��Wn���|��mL�ߑ))XN�����ޮ
n�bL��U�T&�i}k�����]��1�gU��*�V�Ebrz���樨��1�at���gǂ�H�B?��Ԝ��^�k�é1�5���;q�@�;�T_����Ҝ���^`�l���|,�'W�Q��I��" ��iṺ']�s2�j�v�g1}��� ~_Ő�5��]�؁^&���w�m�m�X�L�r�uNz�䜖�,��� c"0h)
+o'~�g��T���ON��6�	�-���S�w5���H��Y�6�C�؇�	_g4�t�x�&:��	�[]�3���~�x���w2} ;Uxr˼��^��ώ��G1d}��,���K	5�a%�~t"vJjF�n��/k�O�Nt��EDܮb��̨�]�D}�]����ѷF�RM�,ģ�B`W
1��<���@�����[�4VaF�a�]�̧#�x���Σ�f�m��ۊǵX��;�;���/����O�.��mgW&�8B> �k�rm�AK�����[(.S�����ȕ���}��t7�풟�)]|G`������G�w��r�h�%�ŎE��I�����֭{r8Z�5�qy��|�,F��"�U]�,ҿ��p(p�
�965�u�	���ϠC�����:N��;�a�Hu=z޼ƞ֘μ�n��7U����u9�������i�O�N����M�i
<'�ó��R�����G����[��?���ܙ�["�:yi������������� ;�xrq�_���Ưn]|��|qO��ԅϦ�6�ߜz�5��N�U~�[˜7������͓I~��c5��|>_3OEI��Mc�Lj[�ծ0���|)�T���n@������H|�xh��sg�;���)���V��>og_P1�Ϻo��fs���ؾ¥-C��q#r��w�-���R�jz�\i�\�8�݉��Xϔ9�a�wa����B�vH(ؖ>g�B���Y��P]�;aՒ�0$��xp��rm��}<�]���$ a������|+�r��'�ƺ�N�%V�X�N�a��2��+�ȑ�����pܚ3�
Ύ��cv�$��s��L�����95�+7@N��Z[�Vf��G`�pwJ��`x��R���Z�/�|�Ane��#јF;��Qܔ�> ���E���k�D%8��T:��H��MK�16�,�|Yf7������e�4=/}xO��Ѝ�H����U����hM����v�V�9T#p4���r�WW�{!�vgCT (�eėy�8��A��y&>���{�g��$��� ���|��ۍ+Њ��w\���+��'��2_r&E��-�l�!���R���>��<��;1~G���ۉz*����^-��U��tG��m���������^(P��M��n8k���J$=��XfK��	s��;pX��<w��U$�D�R��$��$�'��o�ֿ���e7��7�x�d����:���,���{�L�8����Ls��Lv������D��+�Nߘ�]��l[��֭@0�l¨�,���"�T����M"ŃK����2m��U���Cr
��z���S�L>מG���"���:��?���b�ސB���jt�x�ֽ�}����U\e���(������Y�yd��`�w���h�+���aYs��:�ǰz����"���x	_́w)�S�\mwrD2��n���Jz�������9���1[��]Ac &�;h��נ�t�x� �+��Eӡ�5+�e��n�ePׯʤq|��W���𾖟�Ka>�W�Π I|���½`{c�.v�z�����p���}�4Ƹ���ibL2�>/��>��xK������8�\�ty8��6����'�|��s^��.���y��ȉ=�e��>"(��@ض=�����q�D%�_��C��	�\W㿍�63��8���%�� gf
ZB�*}:� HE\����Sbd�|g�2�.�s��@X]��v(L�9$�V�&_�i��L@��l��q}�RP5���X������@�	�m)�=j�Y�>f�7[��5�թ������p�N���#pfc�[ӯ?&�7��(�+�'�Z�'��8d�c�@(��wr�[�q��Fq�Hh.X��i�]�A��E��V���}��#q���fƚ.�z���(���XƲL��$���$��෽��m�~ɎoFv��9Єa��8�tqRw�b	��?���\I����f�v�i�įj�b�m��#6��e���R���7T;�+
�'�@����$?�Ճ���_J��8H��VVS�s$'��!��.5�c��5z�Ow ������b�u��t����q\R+��H��� [Q���Z��&?��[|w�#	z�'�� �����Z	p�P�����j�F@r�6���B&k�u{�S+�$��J�-�v@3�c~��(J��ݲ���E�1�f�w1F-�a>m-�-��Xʼs���{�����u�ͽ���y t�5�z��m�r�K�<��cj|ln��c��zB�R|�]I���eD�$���i���u�gm�b7��G���Vu'Ź��|�l~�S���:V�O/ɳۯɿ��ry�w,����K�+&O�S����ڷ��yn>�:?�������o��WO�>}�������������^�x���u}]_ח]G ���O�>y�كE�?���U��,�f����h���l8i�t.kʘ�ͫ�3�k���o~Un��K9v�
^�ӳ�W%��Gɗf�M�8�N[Yw[��~.ܿ�i)x�Ȑ�UE_>{j��&Q��o-N27��Z��t\d��V�sy�dO���qtǚ�g�ڛo��Ꟶ�]�	j�U@zV�*�޼+߾��|���'��5�a�6]�ҋ���6C��++*�����Ud1��$�v����;q���ֿm����l�Ar'�R��E��F��˫������a�`�xFW��^ϡ�6�y�s��)u�e.4���[g|�"�RV0�:���H���.�c_��F�b΍������İ���ӱqGH�����^��?�g��gS�T�XQ����֌?;�!�3ڌUF{j����up�E=x��|��3Xݠ켑�Q8	�3�`qx���Ɇ�����N/J�W�uD��̸��̸ִra�-'ی|�zQ��	�x�.5��nO�l����Dn�VW�1�h��O�jcY��ΏF�|�!J�l��,��j���/t"s�zxkg�r����c�ϧ��b�D�#�r����
���z֫T���ZN��ca�7�`x���n�
0E�|!��Gc��k���GT��p��=��*',��� J8	tC :��v��ya"�t�����'8��/ׅ��}��.
��@���^R{D�#�Ѝ��#��1
���.�7��ʘ�q�G�ǵ�z��5���L}����Q|�ν�'Ѯ���<ީi2߅>g��à�+z�,�ob�Y�m��:�2#�2����t��D��x5�0}"``�e �uT����1L�S�٬���n�j�;d�o&�k�i�HЕ��<@�˴]e�x�̓�{��A5���9?�#;��Aپ�����lEh�U�X���ҽ��'����;�j#�ϰ��h�
"�J�J� �&��l��!�l9�C���D8�+�[��]��Im�eb��w�%�H����+�{{�����Y胱�8����C��q��RM%:b�.��+�6�meh���$�@��x3op(\���d:^3��r	��9�r)Jũd���� x�愺�9�IpHX����x2��'J��-}c[g�]2�,��jp������T�;���ˢ3��TA�D3�>��;���u� �'����ܓ�Y�:$�f��Z���nz{!��z���}����n�D}�^����{Lg�V;��)q/��y����MJ�=��a�!���j�'^E�V�� ���BAE�����}#��`�f��z�F��AL$��g[t�ɛ�`�5����#>6Ą]��"5�cG>�ߡ+��_��j���D]%�>]�g�v�K)u����s��U��tڮt�i�Ӿk����.������y�+����N%ȁo$�`!���0�n�R��;Wzd�򙀂��w|Be�䤹�^G? �������i t�0lkJv�|��d��z�bt�@�OWi�^_[��#��_?ܔ�����iω���]��o�'S��1�Um_�Nn�;-I�d��I�5�߸Q��]�gP����be��[��zD��ҩ˅f�k���x�\��8�ܬWHc���Vg�+�P|��7��_|.�����y�״|^���+%v�CC�lO�K���7�����w���G���O_��w����u}]_������ZO�x6���k������5�7\�TH����|_g�ޔW�n�a}[̘�Cp6ťb����m�V��.�iZ�9H�N�笖��xz~�x�杋�w.n޸uqrz~yz8]��u���x�O�<էO���<{rx����矞���S���0�/��^��vC�h�e�Ăskk�����q���=]*����'���_|&�mKޣL����1� a݄.+��-�^6��Q)1���0����rȁ�d�г+�A��r��6N�ш�*�Y�Uj0��d�x�Sh����;VlH��[f��u(fT�q�85�����W� RP�+�F8��$�|�h��m���A(��}�`6ж�Ĺ��WS��S`��ƶ�0K�r�s��!�;���������7$����u��ǽ��Y�"��B/T��J�_'��[+�skn�3<O8Cx�>W*;/�g�{�호�s9C�-\m��W���b����㈝�p�q�
����ᆠf��Ȓ[l�����2�ћ�K@�ڿF�������U��eY ;H�pC���J�T���%G�(��B�>a�qd�%��7�����f��~�[��p�<�3�D�����0�d	/�ļ!��n�OC��'~��<�AR?I3�Gg�Trz� r阮�~�hU2|����<X@�3����Hu�#q�ǐϹ��
%�.�̻��]�Esr������9�3�0;/�>�y��[��&
��㌒M�`L��@�N���H����M��[/����r>Zwq��V����*��<,���i|�����^E����F}s�g�_��F�-]�L�	O��N<�{S�U(�H��	�'�������?vĳ�F��ż������r��#�z�8��e��&i�ߋ�A¼�u �v&����{|;�ڹZ����\A"R�5:�w����`��~V����r����9��|�q^1�cPTz6���)�L�J�b�y�!�.�:i��60��9�a�+=�NGllj7��:�_4���u��9��H�{Bcտ��g���1�}���a����4؀:̬���	��`����G{�o�_ Hi��go<uěRb_�i��kg�0�͒v�QI�YM`cl3�06p�B�� ��x%n�x��N�c^�-�~Fe�'a�陵T��
���׽�ۡ��!X���C�^懡�0ݓ�~�t��g���Cpd�C��m�G��)�����E��}u��o�r�����	{�d�nY�%#χ���sr�<�O�(�~ӝ$`y��,G}��9oU�x�"�C}ܿ����p8mǋ��0iYo���	��>׭?v�$��{������.�@�q�P;�jC���OP�Ms	[У�(��>�������I5>ߛ�ą���4���>�����#v�Q/R[4����e����_�#�О�z��:�<,��ϲ5ו�����E�������_/PV�<=_��-7��k��pS��Ƕ[���R0���(|ϵ#����X�������r*�t[N����盷o�۷�ԛ7o��pR��<�^^���<~�X���~��S}��S��|Z�ǧZ�g���}7�w� <T��OC^H��/�a=����T~�ͯˣ��D.��v��v������� $���{VЎ�x��r�t�ȹ��d'��������k{�}$ �w�rq��K_���=�|��J��f���[�R=��kV�w\���ea�*'� 'z!_=�)_��J���]�8^M����Zͅ4��2�y��j3�t��T���ZO/���^��O���o?��ʃ'���}���l)�\d�۪����l��h-��/N�x����O>����?�������ӧ޼��䦔����|�L���~�g�����`�S۾~�{*}��D~p�u���O���YK��G}+ St��9����/�
�Au�2D؀򚼯|�?E�B⪍)�l��I�{q4 +.���J�����@1�x1\�k�H�1#�Vn�[���QL��K+����*�-���+�tS>��F�>�����"���[�5�H��UOAP��+�;~#��6�����b6�)��XF`y�N+�sDw��pZ�4�E�ٙ?*��w|���D����Ql*��dd���ܷ��r���C+���`s�lp$�
�F��{��07v<�t��� ��y,�1Q�\^#�����>�!˒C:9����W�/D�j� ز�m�-v��Ԓpfw7<��75�C�S�|1+�]E�F.���l�x	0z[s�B#Ƚ^Gs�l ���"�������:B��&����s|�~s�j\rJƎ/6v��l˲���6���1�)��7�¢�X�bc��!�}|t��>zҨ���Y�*�ӾJ��!��=SrU�|5��ٓ;t��1$<%G�p���q]O~���F�X�>��t�lKJ�]��X�]1����w�P���J�R<�F��~���35m�	�w#��
����%�d5gUug�l/:G`}C��r� �7G ��&y�*��^��A��rbL/;�z\�c���Ď	�צ+�$E�́�-��	�n"YС׹�������Q	>Re;%$4��y�0FK�0��he��A�eʼ�[D��s.;����9����CK���C�uq�����[��õ�So��UۊA-�u1fq�)r"�;�ӱk}M��΂txi70�۱-^ȸ��ʣ��Sa׍�b\Er ��8�亗8���:�2�k�}D'1��}����b����G����\s�c�Q��૤#��D0D��Gwlml�<�WSw��a����"��۠���yQ�Z����mcZuh��s�J�լ�r�/��=�����g����&��GypM���9nP��$1���R_2?���5�3ؔ�C�+_�xp���As ��Q�0���ӽ���Q�/Z���׋�7��?�^��S�C]i8>.�����uθ�蟚�	�N|[D|�C+�)ӹ��S.���?�:����bdn[w��UT��{�q���y�$^ ��9�M}`�
\�W��Y'#	�D����f�zu�{c�[�s!3�������_�xl\S�����68�
� �_[_��ѐ'�N�4��VM	6!��ޭyd0O��c�ܦ�8�+��v���g���6�<��*��y��ēgN�d�v^����y�ی�k2�mN��~ąX���bT�6�g�;�����E�q�ѧG)'����vi����V:��6զc�}Ӻ��d��YK�9ߺ�j��7�+o���|������ɪ��}�*�����_%��8���/?�Y���I��ÿ����z1���R��0�8��>���>��#*ڮ����uI�26_�qG����/~!��i[��d�Á��
���*�Y��gj�r�*������}��7�ז�ƨ\_���u}�__v@c�g�ٓ�ܼ����ӟ=?��ͥ,|�h6��0��y����,��i��������u3(0b���MU���RKSΧ�s���l��V=9�����O���o}���~�7o����p��_ꤏK9<��x�|����˶����i^:9=;���<{���;_y��=z�����7��?��[�?z�a�Ƿ&�NkdVd���"W�75&��]3^�3�)�؜��[w�/�.?��{RNq���:V���=o͕Ce8S�G�@5%Z�b���"e¶�޿�)v�ƙ���UW��x���oo�&n�暲���i
���*�
_��Yɒ�N�T���7ũ����۠-4>�e����`�b�Il���8x8���-m���h(��_��3��m(C����}
��1)�v,��>T8g1��6����h7|i���- �IP�������錷��1]ll�,i�
M��]��{Ĝ��2��s�7�ƈ�c�'pX8�!�\�C��Tx�u�69V ��U�s�4�f2�����>�=ۉ���0��Ϋ���@��� ��I�	�0�H�/���=���a��Y�;X�y��#\K����"�iOjB%���wgMsRD���pS��G~ �>�
݈�;2�O_��G�ʏ�������(vΣϯ���\~V�q��Am.E���z$�4&�H����s?�A�ˇ�lW���fN0�o�����]�r8��r�t����!�@��J�󯙏`��l��)���`��^�8>��9�����׵��lF:�d�΢��f�������f/b���>���ΓH�X_8ƣ�i>�2�O�C&�Y>[c{�
� �ۼ��`�h}�wM҄�M� 7�4V��#���Ʈ�pFdǠ)p��k�Te��a�|�V�����$;}��'�Q����\��w�8��o������+�x�'���:�˥�wԩ=$�	�a9�ei��V@����沒e�6A�S/�ey���g����������"��>�͏� pذ�|h�� g; !	{�+q�4t�<,QV���SQ⟭>.���n�A�<5�ȏǮ�Y��y JG{z�v�J��n��p$Y'�O*0���	�B|l�35xQ%]���6�C}�&l<wJ���y�,C����L��PB�ไ9������
�@/��U�_cB�Q�"V��n��\ݠN��]s?��_�9 �?����<���n#�?@�\j����V��L	��=�ߪ�q{�����
��
�(QI���zx�a�Fr�v�^(pz	��V�q��{��:���9� �S�H�a��7�H�{����ɚ-,:�CpIu��|%=��@4��y�c�\�����b��ۍO���f��c>�̦�<K����j�zC��z����J1�A������E�m���Ҙ:���P*��_ac�.�T�7��tw~�iS������21��O��2�tx�vs��W�����C�D��ԓYZ�r8�z�*�����ݞ�miӎ�]ʜ,/�/(xxz&�}��ڹ��-�ԋ��BG�}(G�����яr.� �ᬞ�ܩ7oݟ����<��ַ�Í�yy6�E˛�.�+�+�^�,�9!ǩg�,�u~�� �^��_��7ʧ����G?�˳�����i��������u-�jZ�Ikm�z�zI���'�v���9�>�K�������?�H�/���NEk��<�h�m��u�k��ڷ�^��7����?~��ݏ�i�t)}���]_���u}��KM X�rͷ���o����'�~������޻�S��k��ei����������2z��dyv�<��K����]�^ޛ/��zkgfγ��d<���ǖճZ�m�r��r�������G��s-'?^���D���������U�4��5��~����N�Y�q��z<�Z�����w�}����_��?��?��W�?����O�e~~=�����B�,큪#����gۙ5��P�[w�=�@>�|"��=��4�Q�2(�>*�Ԕ�J��l�#�B�j�-^L���F�f��bsψ�J�ol��+�IA7���������l���LN�v�އ��U��[\��};kk�t%�����N&h���'���"��}6|$0��V x�#dX
�����A_�C���c�*+�l�^�v����^�� ~7�q�T^a�H2��wr�Ɯ�nT(�B4J+�2vcN�����h$��HE�����9�W�d�������H���}��J��t���^5��<	>�$f�*���ۖ�W;LG`�3oP@?��0��	���D���n`�A5q�J�����n\M?�C��Nu�*f�VG��2W��;p������yk���|���K��4�������{��iO48Ob�X����b9@��Q'�nx�줗II�Ǭo#�xb�x�ٴ(>_p�yf"��Q��m���o���(袯�W�{������VH&�+�H�YY�:�Zi^���߀�jc Zg���Y��J�ӈ� =^kx��i)d9�����q�)��E#���=X�2F��xD�P��C�{�a����x��ve~C�������ت���yr��w��!���Y�	Fc}�X����Z���X�t)�|�.8����a�o���cU	ϼbx=l+�ǳ'`�~�˒l2�;]��Ir�8(�U��~y�$�rG�5�F��躸Xϡ��Y�AG�Q�y�
���)�6뭳W������PP�99%�k��S`3
�ۚ{�8������ㄹ����~`U� �Rʗ;�c[n��̓;����W�����03bD%� �.B.�'T��$ۿ�)�c$�{�x!P���WDW�P/����Ep9Tg�N|�uB&�vpX9��� B��s�I�.�RUՇ���yʹ�؋qjI׆g�c���${C�oy tn�Հ��~�s7d�z�o�w�G�:G�g6w��܃�Y�c$���U��o行<�Ŏ���do��3�h= "dA��No��E�\$^˻����?D��cl�8��vz��4Ț�y������1l�.�o[ޚ��"�GJ* �MzO�h��J��<��mn׍�מ�QFg�q�<��vx�W�s���"P�u u�a�t~�Hmu��2�- Of��hw�h�9�O�^7���ߔ7X�����o�}[p@�j��-�=���gXC�"���_���B��l\��]��W���g����ӝڷqQ4`��)|T��_G�"���t~Vm������6ȏ&�Χ��*/�w-�B�OWXNp;��f7\I:�K�� ����7�:Uz��kޕ5�Y�t~�[�3�x��0��i��Nt���'�Y��7�&w˩�)��M�k��j��6H\�i	У:L�O� �r���߯����;�������/��e:�K��Le�|��^��3/𮱜�Eci��:�񸼻�q:9�WN�O�޿���_;����7?��_�_^~t&��@�:kU�SgE��V=��d����� ?x�m��ÿ�'7&94�2�Ԗ<z[®�=�Vw�ᆞ]�����G���;��_�]|~&g�r}]_������K?`e���{r������<�ٿ|����ѳ���&RM�� ö5P�{P\�V9�W'�ջ//L�����%h�o9S���=��jl���S+��wrr�N_z�շ���7~�;?�u���L'�<zF�,�|���L,����?Y$���?>!qF��N�f}|rr��Q˯&�����/���~������k��~��|�铏�gw��|�l��"ȯ0�Xh+Ԇj�GWl���7���ɣ��3��Jԧ�M��RZ|uƨ�A�#Zܰ�P<c�����f���4+kI����U�Ho�wnu�m��s gP��Sա��x�06%��+��V����z��I,S��-'	��(�@����I�T �W�k8��x���lFCl{O`��3z�9�>0>��3��;W�"X)�f؆���f'��2X��y��a�'�ʔ�ᶕ�N�իes<g�R�;N,����+���f��ΜBc��#����cL�����5��n|c��� UqC�����o�|v(��#��wV��w�w�"�5nřIN���>�\܎�fP@��5������Z�y[��W�qUF��f��<�y%�8ON��7���+uR���)�he���3]���\�CU��	b�vi�}�g�ʲ1e|;}�3�`����pTw\mr�Gx��4����}5R�>$�D28t��AZ���q_}�ݥ�<�Q1��ר��Eζp�^���ʯ����O�&��hl#98qz`
A�8f����ޛ��\�a�j�;�ܹoOl�9�I���$kr�r�A@� �<��[ AyH !����mB"E��X�EZ$-RT��&{����s��+���o�ߪ�o3/���=����5�Z�Z��+��;^����Ph\ÐL��eʺ&b�l���q"��������栓y�ƳG�;�#�Y����4>���D𐠳`,����bh���x�	U��@��3&��5Ӡ����㲎uYh�\�<�:��4x"{:����SA��G�	�9 ���i��(�
����]�<,�;�7����E�}�o�;h��Q����~?��D\F�w�������Ή�6L'֨�&��I�o$�#v��V5�3�ד\)Hk�@z��$�{=�YK��Yn�"6ѧ�v���`��,���W���jߍ�َ�'�?ޗ���x�����rG��И�/o���vП���k��fDS�����#>F�j�A%A|��'�:x�I|��S��5X�x�A�Mv��N����3o�@HN��o���3�u�D4���6)wL�]�6�8.�V�:�O�t�[o��;�?���uY�Iy!���yCw�mr���<��I��?�����Iw��:IQ�ޣ2p�y^\����Œ-���h�tǰ�2��gLàq�p0o�~����_�A$4�Lܿ�_�6�sp<����M:�u��D�i�A�&��%i�/��=��JT
�8.K\7�l�� �eq|[��3��n�f�ɇ�ǳt��bG��#�C�&M��U� ~Dp➙CEߣ?c��c�n[R��e4��~��wp���}�#��Y_1�=�>��e�t�Q��h�����܌X�>��F��dܞ��*7H�)����*EX?�Ĥ�d �wJ>��eMhU�{[��V�]j��b�'_�}W^���FW���TC+�F��]��S�8��r�&�ӡ}����x�ܹ�|������3����tv~:L���<��k�Im�щf���N��M�S�]�;��̳� ���T�H�峏_��/�p�O����׾��N�o�.�G���.wژ��\�<������^�?��k�UBX�66�U��hiZ�e���t��7~�����8����[���}^7��us�\Ͼ>��z�,/_�~z���������>��믿uZ�ޑ��z�*����h�1׬1��޽/�k�Un���峡�%8M�Yz�Z�8��ٱ+c�n��t���?��o�g����[�
�?�g�\�}g}�ɡ�� ���L�W�P{m�b�}����[Y.d^Mxr&g�_��wR��9^N����-��[�����<yN�����p>�b0prJ�Lxs๳��!�
�ZgZ�����Ͼ'O�ߗ��2Ô��,�ޤt4�F�%�����U�okד� ��jF�0&u��:�ж;��MQ�� �������"G#5�mFeԒ
�T��zA�#�=fd�A��qs��%Ο�cN6��\�1*\�^�s0<uW���A��㎋��"X�]3��k6���&0IL�Ue���0�k<�O�V�I��x.V��1�b�M�/BtQ��6��$�����L��c/C=B�%eM�.�YyP��
G���mg�OB���a��E�>r��!��P�s��xf;�`�E��8w��#Zt����wtVG��e!��O�3�E�t�چS� �,�1q�?�o� ~t�;{f�
�9	W�3���z��B�:�>C��,	�mb����Y7���B01S���<�W̘_(��w���y_n�w�Xq|�;u����~��/U����H-&;��	V���!��I�b�P�iRSi���[ �������iX�0�q������ Bs"�����gt<�)0������n��W���X���(J{�`[��������W�r�$����kr)� �iB�#}Q�d�\�
O;�\�P2�Y<���P��x�K��B��[�o��ݷ�:Wr��F�gsx*]�	��0�_�ֹkO�:�M@w� ?'&|sh߬��%�ؿ���Yv�k����i]�]�������>;qY:�g1���@Sv^�Vߏ<��-�����.���w:��9Y��=}8�e� |^��)oޕQ<�{�7�d��q���Y�p�KX��_�/bB��aͳ�͘�>�In��, ��L��{"x�I�R�8�\�Y���2̿��ߑOԖ�H��!�!�]}W��j$&&�=u!�c��o羝Q�|-8�-��S�"�s����]}����_��/v�fK3�� ����?F �;��$l�2�CC"�H�K����7�l�h_�t�eڳh�ɶ��	�А���.����$|t3�~�����	=���y���{����j<����U�jQ[���4��iE��)������ȕҰ#�¸��f7��<����O,;3��&�擌7��5����m�0���m�2�z��K��p�N=���hTnU��x����9��.성���78mŤ�A�d>&�Y�����
m�����6p�.�w�?%��-ēc��^m����	�� 7��?�k��k��| �6r�·� [�����1w���լO��>i[�}�.ZA�%ҵ���+Y�1��|�`c^
>9Q��0��c�KG
����%�C��b=���MEa�}N"o��+������/�m�Ш������+���Ep��Ӛ���̳����ܻ�����W�ⓧ��ⴶy���k�vJ5K���)����]���X�uW"�����Z�����$K�p8ܹ�o����ңi�����)�r�����)֢�IM�^��|h�<V+4� ~>t�[u������"�}�5�>.Hݰ��k�mgY��uk�����w�Li��᰼�sz���\7��us���I�z�������=~�[y��%�����-@�E����n��鰲��� ?r繕5��U��I�E�����Y��N--K�2ۥ�Mg�������o�+������_���Օq��4�wO��_ӭ��U�&z�'gg��<I��]Y���Y=��y}���Yy�c�x�W�߿������|l���
��P����$ƻh������^{������_}��\�:\�@�]��av��9�t�+F�gi��:�Jrb;+ɔ<'1��&�,	�(Yv�21���E�|l
��oɰd����:��Ş���X1�Y*dT7�(<��g36ųh�LU>3�N�%
 �*��l�#���hB��4.u`���V)�S���۲����ޛ1:��j�s�����9}�x�x�$�W�.�I�:�	z?��W*�cs�³�E�]n;�%�"�BM�c��Wl�?or֨��;�\}nq���n�g�_�)fr���G���p0r�m�2��`T���h���NPMԈӱX��6G&2"�� ��sUzoÎ��$:��Y�f���n�F|1uc��\�р�I �����i<�nl�NorZa�d��`LjU��ʀ���=�� �fW!�[�7gh��R��
*G������[��1LLZר�7�;��q��U��^�Ƴ�K��i�H����Sr�ʝŎ�qZ�J1��$_-Y%����:_�S�)8p2w�JK�S��p��>�M�p�B���@⢁c]Ã��
����!�H�$��d��s�����9�Bp
��8߱W���.K>Q�H��.'�����H�݅�D��4�S}���d!x����8G)H�$&�q��;�����pMtD���݊CS�3��k��l�c�=��;�d� D���qtPr��HL��(�(�w���w��W��iP�~�S�,#����A��-TW.�	����7Kȼ_e�Rf���8�>�����8٬��Dk�Zˬ6��7�N9��h[�ugw�kt�-�H��:.�W���)S�9�4z��ф�w�!)^�e_��"C:Ih���_�x4�܈F<�OA����MG�wXK�Q۠��m�~��>�i�MIe.�'�M�ǹ^"�s4�ш�������6�K�9��ڡ�#_+��ֲx��5[�@��/T� !��\��/��!Ǉ6[[k����Q��#ʃ,�2�Y�������Z�R$�=HK����`#�^-�磂��k3
����Z�G�|'��c�!z\�0�@(��G��o�iCT�`(��VЙi�lZ�]Lpxd[�@
&�s�;c$�bcb{^���\��$�Ϟ��JK�2���=
�v;��`,DV�*7�h�v�;t1�d<�wX���2���H��Þ��&�ka6t���m�=e8��`{xΰ�t�����G)�J��h��o����i~� �gF9`s4\|�6u��<�����g�K`�E���6�d���<1�h�.g;�+S����J?�o9N���g��G�~ׅ�dw�d�>lob���{ʨ��8���zo_y~v�7���ԫW�ϛ�m�_��B"�d�����LSU:�T���?�|�ָΩ�Y�u,�.�R����}.���鳎�}HHe[��G�ѱ¿<^��}�ϒ\��<<�%/߽'��b1�~�$�
��_T$�h����JH����ry�������{���i�����jDթS���R�Ȅ�M=�a�'��`�I �}���ԏ8�Z	:��kߧ9�������,�W����'N����t}�JΫ�M^�@�:����N!74٥���/B�������u�k���n��k^J�9͵6A���{Y�r�⹚��hI�������n���溹�y}�	 ��Ho�����[o�������߽~�����b�ns�ؙ՜��ny5klZy�g�</��cc���kU���w3tj;+�n��6W����~��_z��_����G��Y��v8����h��<O�k[��+G���a�Z"�����l�MX����a�����iz���_���{����9�"�E��9=9��j��e���j�_P]����ʕK;a����|�%�[��+0�&���"�!&�D�<���˒Z�tT�QGXW�'mI�y��|)tMR�V5t�9��G�f|tTD\�zkq%���5;d�6��uq͘�q�#�QuɟE�S�@�����N��9%W��P3�x�]�Y��q���;#��S�,ꮑ
P<5�����S�Î~�pf'Wr	|K�OZ�z4F��.6� :5�$����-��t&����B8J�� CO ��� �V)�Q1F	z,Q0��dkh3�@��b�z��-����%P,9�ؼ����BL��w�*�/E� ���0.�>a���@fH�����X��"g[h0Y̥(~�M��yJ�7�IKZ�}� ��8@%�lI�j̲=�(O��7N@�~�`L��xy'v�`��J0���g�?�0F����)���v�.6�YwEڵ ����8�G�g6F��`$K��<�q,�q�����֗'�4���8�2�D��Q2<P�ጾĂ��(�Շ���!ρo�=�yE���P�?$�Q7,��]��������K�F>�m�k9a8G�Bs��5��ex�䰢w�%����.n3M�=i�O]Hɂ<gѱe]Ә��]��؝��]�wR2�ږ�:Υ�z��Bă����n�?L��.+]��>F�gϫ�`}A�:��{9,��>�0D�3�+|���oI�d��&�3��a�^���5�{R�˫l��n<��R/q,b��w!�{ۓ��b�e�#YF~����NE��j�~�F��xk
<��A��������1Iak�G0�v
/;&�؜�1��aY�ߝa����R0���b�9��'[�lz��)�XdG����3���@���ĭ���0`'�˅�N�&Sh���`�3�$�����N9m#U�i�Zw���9�@�bY���3��3%�����ł�YF�8��{���A���/�����3M��5��N����ӹ/�uO��z�ը_��0ٍ������M���œ(�/)�7V뉗��@oa�d�E�>��Y��I�q�����)Ll�A踖t�Dr�S+�Xi�8;S��n(acg6GE����Q;�\�8o�
z���6wi�`�C�:6 �l���p���*�&M�3~�tg�+�D;k���6��_X��Ť�N"ެ|���/H�a�*��_ӵ�)NFo6�S�W��K���� �F��4�n�a	�n�R��(b�l�4�,J�"q~�x���,�܄@'٣ǌ?��`!�MƟ"��uL*����޵%#1���?}v!����Rq2��$��u�T}����m���W�Z�yA%5�]6#}8^�pk�еl��z�{�Sq�x�M��ܖh���,��h�D7�a󩲌@����뀷�=Ø1�*�#��1G����>�9� ߓ�}���O��: +���A�wF��qz�K�KxE�k�8,�(���x��>����
�,]��R���W��U��G�ݓۧ,�E�.'9UM@�q�np�-�ɃZ2}M��X���|�����<�����p����,mL���SW�N+����`�:N�qN+���i]F��vyZ��ӵ������4]=*��O���+O�߹���~o���jQ]����fIw����Vn�8^�Y��9�4���[����%o<}"�t�g�����:]���������"o�O�k�������|}v~~>�� 7��us���#M (}�����������۟�����_|t.��e9�e���������]� ݅u\��䃗,S9��o� e���[`X�\����Lg������������g���_�r�/j��p8���t��s!���
�yn�������u���Z+k��Otp�����eY���K�~�W�������9/���TN��cP��t�J=e%E������
�[gG�Ľ�����/��+7UV4�C�V��T:�A�
��Ϝԉ�g[�A��)(�0Ng����;-L�PM�@S�|c%�������~�N)8�~��U��LƆ?�kȊW�Ř�M��I����EMu�3���҆�1���k<�>�A�XǇ���4S�A9�����)��%��~�G'���+^�G�w�pa���ߪ|�CSԟ�H��mA[u�����Y�$�@_����$����F ��k�F�l�DQ��"k��2:�DlMAk�NH6n$�iT�ê�IqH�F��e��9��������=����u�� 0�1�������<1�1OY��#���o(O0�	[�V�s0:�k�躄Q?���
,�_0:O�xw�sCd�GJ�48���'v�z7�0�*�lO�!^ő�����GwI��;[����d�U����i�n�h���c �5,����;���B0%�(-h�	H�y��@qpC�S = ���Ì�2�ع��!��E�{!\'ڱ��xiX;�6�rٌS��]˔��A��#9.j�ۭ�
e3���K��<�]Bn�L�Q��`��}��0�=`���)|�Y�;��c{�4�iUA�K
�#$���ߢ*8 �S�������`퉨�>'�����.��hоsJ4������~�3��`G�%�;����Hλ��n�m��k��������Q��wM�3�����w4�g��̾n��9�N�\n��q�p�9�V!��t�G��@ǻꈛ�.8��As���#�:ObL��ew"䈅ޯ��v"1�5p>�m}��l�q��6 5��Y���|���|���߇k�9�ư˳N�y����O��Ph�HV�$Y���G O��V��&]f��3h�G�)C��CIa]#0eǳ��+�J��´����:LZ?����wf��=o�e��R��N�=�ݓ=��xcI�:A���1�Ō�_�Jɐ:�0C
�{��4S xq��D�/��%� �S�I�K�Z#*��	dQV�^ܙ�p"��}������u�G��Q5^;�g�WB蟻_��x�m�,Aߟ���DX^�, ��08B��Q<�-�^�{H�`ɺ�'hO����$o�]�_J��(�|���F^�����;&C�ժ��8kp�ݟP&1�-q׍{?-a&,�E;��v�z�y�+K62{���yH V��	{!i���b������r�)�E��
�h�_,�Z����, �V�q��!�l,��^��Ȼ0�x���=(��he\ȍP�6Zʺf9<ºYX�����/̷��ty&.ͶL�\���l7�uB����8oA%J���/8�c���&t�?���-g2�A����-(��%YwU�?�������Ԓd��]���W��!��-�-�[�����ߘ>|p:���ᰴ�wP-Iw7���k��\����?�\��LX��W��"�q9�I���_���o����k����z�@��IeF�l�Յ<�9g�ߟz�����~�Uh���'�_��s�#j1�r�ϯ�����{���/��O~�G�p����ts�\7�͵{}� *�?��?�����޷��[O���ӫ�V8���k+��
^/5���fu�/]ޑ�3)sy�rUK�]���tAEP���5��b�u��ǿ�K����o�B�k_Ϲ�Y��ҙ��djc����v��Z>f�Ya`�&,�J������t)�������~w���������g_|�[_���?��bJ�E*K���<��Ú)Px����m��i������w�/���|`f[}W�@�4��C��X�N�I�DV\����%��safJ�9y]A�F)$�f�����-�ƻ��(Jh2�ݡ��x��]�����3{�-5��)v�}qP	��h���;��L>�Y����������W4�`��� u����P�(ؙ��C��)Y{Q)�C Tb�FA��p[�s��Aў�Ѩ��c��F��X���HA�`��u:�9�R��L���_�R�@��()�����Jٗͳp��q�� d�2��Ͱ:8<YhEt=�iA�/W7肓������������#πY`$9�K�g<K�3r��m�x5��PfB�n0xܠ-b��B�Ԇ7�����b
��2��P`|Se��iwƂ���|�ߜ7$��l��7V��:L��B5h�2E~i�E�J��A���F;���A.kO'���0cOAYv,���QBz?�	\d��蜰9(́��1��)0:>���4��X��t������p��5��TbӃ�
����6����"A|���`�g�'`NN�p�;2&���^�a-}
'�;8��"n8^���k4�v��y���r��3�:mz$g���dt���f�tЙS�h`������G�]�/x���B�����8q�=�S:®��N�X���")J�3���H�q�Կ���"����lЮ�d]��y'����`�Wg��c=���<6��y����!�UI'@5��X �y.���L$�#=Fװ,q[>w�")����oFb�h��!y��b�t�2ܴ]�β=�d���u���?�oT�"��ֶ{�m N�e�R��ӚI�L��c����Fa���B��(�]�Izd
��AM�W��]�D�-��[� d�'Ȣ>�E��C�eY��9mk��I �~�%��lfF�H��;Tw`z��s�=�r��&�Lce����ȴ��>��C���3V��.!���n�3 ����z�m�$�����`�[�$�nG���M��%�[����h��P�"�a:	�SBcw��f�@��G������5zC��ŋ�Y���Ў�"�n���g�4��e(��vd��A�E�o����^��E)�Q�a��6���3R�U�pT�N�w��>��$;-�p���=�&�r�F*��+x�\�!��}�Gi~]�i�G�C g�IK:N�g��RWC2���%�v,�A�x�|N�E���$1;'��Ӵ�'�v�V�C<�
#��[�_��g�.��Ʈ���t�����Y���t^�`���6���>�dk���U?�@��'����8�I�>��4/v|��e�jT�7�%a�C �-|�~�g���~n����6G;<������K͜��.ժ�i��2ɧ�>/�K�g�6fkS�O��jm�'��w���s˧?������$��4�H|����I��O���̜ 0/鴣Y������;y��*�C��tx��ܾ���~����?�}]���<����	��6\<4~[�̈́tO����ⶼtvG�^>h���g��j��\bNO�(�r}����7_����/�������ԧnߺu���溹n��k��� j����y��,O����++<>]�Ԋ~O5��|�0C�u��P��>}osWoj�B%&0�Jߌ���`�ᦳe:�{����州{�կ�|�G��\e�������V͞���iZ�Բǎ��&[�O �O~r�p:�V�Q�<�k?������7����G��Y�/�i1�t�Z慕�X�N���g�����s�\�*�[v�u;;��ZUi���*�-㽠��+U����U�)�\9�Tq�c��j种Nls2Gɲ���'8��4����Q��v��;�G����'�`k�34SI�;wxr������c.R<����{6}q�F��� �֠7���>�9o�k�{�'��D��B���O�f��w0*�֦����^bF�a�9����IF�!\�Q�x��m�B�l]�� Cz����Ci_<�%�Ә8�6����;3���2���6�X❫L���=��^��2fu}����ۧ�uG��GM
9eZ>V�$��j��vN��ϰ��x*��!��Q&p��1�933J����5�N�x���-ࠗ�7�5®��_�8v�v��n��nc,���`]����O�pK�_�J�R�?���=Zr��YO�z�����Gr�[��P6�� 9�%V1v�d���4���1�>�a��G(���H�<vx}�q$G���q�R�������ȫ��|^i��=�����
�����+а3�W�b+�h����j%^�7Ok��+3�/+�h�Q>� L]s�p�F�`U�	Eu���r����u<�i�y3w�-'������x�N�};�mf�V�h���&����v� b�������Q��������R);�CN���:Y��z��%�VW�&"8�al�(��KDt�+S��ʂ���-_[���� ��ɓ���2̅h'\{2���*�d���Qa�P;�G�^��sAWy�P���86̯�I�FgT6����I��H����ÙϤ�3�L�Z�3�<������PNA -���]Z��(��Yo�[�Cv��I�}�5<��yͲ�b��a���3��'�bl4\��W����t��l]�q���t�/��Ҏ �:N1���t���7�`继i���X�ƒȠ�%_}\Tw�{n��}ۻm�8������F�%�B�@�{~�*�N) �W��o�K��5,�����G�`�l_|X ПqX���1�'��SA?"]q�X����V��ݦ�����;���M�'�O�����
���S���v�Z�ͳ�n�+�a��ߏ<���M�ѵ��`W��c�.#t<aV�1�d������&�IK�T��v.�&q��X��{a|EL����bIN4Gנ3�DI+�ǜ�1n�&�DIV�+�U�0�_���E��hc�o�����_���9��E�TY�����B����_lq�3~'+_D����^_F�S�F`c0�F}�5i:X�W�88�`׉�^��4T�[ь��E۰�L@���t�*o�r���u5�o�7ܫ���qr�ăF�6	;"�'�M�'>�2�N��6�y�D����?�jܠ�GE.�A>v�LVرm�~R����^�k�d:�U����?�3���S��i�j��"&�Mi�?5�_�6u��#����x'	#xG�UeIg����)���\����$Oy�֝;����_��������Nr����s}͚���v��t�
���"����|��o����ĔFۦ3�V�[KZZ����a����X^�����_}��Z����)�-�\7��usɿ��z�x�A>?�Z��p����*
��d��XuE1�n4^���NW��S�Ǖ���ф�f/$�v~�()_^?��'���g���z���v�v<���鿣08b��[�;�˩<=��������*H o�U����)�7��[�o��O��Ͽ�/��?�_�i��S;�,��l1�
���zU�\�I�_�kO��Ӯgu(ByT�;�R����Ea�.��ׄ���q��E��e�D��\�O6��n?gp���A��F�L���劈�7F�D������x��h?^�ӕ3�K4�ǀ��)�����J0���l��Pc!���4o��`a�V�{0����{⻓E�L!��:3�b`���<냖g�;�&S�J�mnc�n��H�)�\w�8�c,IT���0���#�U2䊁���w�a�9�$2d��1o�E����J��/��3�����gi��*��wZ�&@�iT�Ov��#@l�B|#8����;c�����F�D<�y��(2&o"|A��v	����<��wp�sYˢ6C?�B�P}���ġr��?��.�QK��w��a[�p;��9K8�sV�uVL���Hf�q����&��0��oa�TT��ΣG��0�K�b�b�eo�i�5s��3�<+�V�	^�B^�&�o�@���:>F:J(�K���\��b��)�����`�3\��W=�O��NS��i$�傈�&��G߭AAƴ�	Wl�pv�;�^��ו�{_^��$qve���+�{��v�������:;6��Ye�(��>�gNBM\b�����'TN���+��c���wfr�Yk>�ݰ_��'4P � /�ƶ=S�˳Y������/�#�Ơ�X�1X?����Ѱ�go�P|�?mm�?�	)�CO���u�u�[�:J��3��4mR����>d����90_����v�3>��lnf.�Hg]�<��$a���h�U��:Nq(�8^o�jA�ǹ�\Z=�Yg�N2����O;k�p�y��Z��F��5����`L�R�زM�U���zˏ #b�#�1�F|]�f�>`xH�5lm��[����>�K�S��]��8��k��zq�.:�7=Ȇ��8P�9�^ ��U�>�^�V��1���7I�>.o\2���2�8�����`tU�tq}�'W:��%���O��V	���[_�hJ��|��@O��r�.����0^�c���t���	�œs
�+��ҵ���	�a]�����	Tw�7���X�-A�K�\�5����x�~�{̇i�
+�g��Ti"y�{��q$���t_A��R��H)T���lB�E��_/�8�רՉx�"1`�����3"?��R�BC��=p�[�09`e�u���V���F��U0M�]X���:qs����H}�������ɒ�5a�(<�����B2�#
Y)>G�C����-�����;�X4�T}OG#���~�g~�`���}S�CJ�1�x�`{���_Q3�v���٤Y{�j�����q��Zy�q������9�K�k�������W��!:���@�%Ow�?���֝�s�g�[�������-�v���\�C@��>Q��������r����ی��Z�W�4�W���~�g�|��_?��o\��tVN�Ss�t�$�q-h�:	ê�e�*�|qG�Ny�\�AJҭ�����8n��k�kW��w\<|����}�g=;��溹n��K>�����W�{�ӏ����{�{�Σ���u5ЮI�q�:fKϙ�%�^\��騂gj�fF�-��P�]�w�Xϣ�ҡ�MY�;[�����ʯ�~v����p����_����?v�w�x�H���C]��l,�!�Rg���Բu�W��9+�?��?��?��֛oV.~\�~��ԕӶ�rHa��-s���c�)ˋw����[2�1R�\�嚑��p�m�]�ʜ@�7�������o(����l���+Z�?�䱂�Z��ݽ�/W�SP:́ENev���Ӆb�E�/��&hj�I�}��MjEL�s�}tdE#%�ĕA	�P�\���0�*��
8���]���b�/	���+P���y����8�m,~��y��v��E�paH���],���u���U�X>�A��C�ݟs�Z�9ۍ�UaԝW�;�ù��ѳ��Y}�ML~����;h�s�Áʕ�G��`'��d ����)�mK�k��[�~}I�<k-��?�{�,�%�	�#�܈vr0���ͨb<K�����g�j;t��0੨��G�^t�AyxBp0��,~K�qE���Yq(��<9,u�.gėy�9�0� �p��׷��E�-�0�m��2���wpNTƝ6���� �Dl�M�cC�o6�u�P��8���v���$�r��� r����e|	�ݡS��['�6٤��%�$�o�/(��@�IG�O�F�K)���zg����;����)�٥<�@�24���Yq0`��0�`�7f��t0�[/l�A�{8�i�r�'֮h���:�N�����b�{��ɀr�'�,6.��;��C$O�grt^_ �7^M�E
';��Ч����q�
�F}
M�$9�H*~�3z�D�m�d�� �}�O.�Ir0�l�*�3+����4�谫ߐnio'����s1���χW��!�`Ϙ���P�$�й�Mk�e�p����
�,H,+mG�J�&���̗��BG�����Ÿi�3\�<Ԓ���'�M�� ~�w��٢%W�h�v�h&V�˔��"q}\���Ye)*n؛f�<���]s�=o�����]޳���� NC��X�Vf����$Gj���g�x�U���� �dk��`}T���T��y��Ve����v��O�����0l�P$^��%m5ځ#�E� �#W�P�+��7Η��)��?[����
�`�|4#ܳ�Iq��e�e�u�-8��$�a�����w������f{996����k���|�a���)�A�R��+�����8(��=��ݖWe;��Ŗ'�_":��@��']>�+?�h�l��.P�S��[�'���qT��}$��})�2]�]�Ԡ���]F ���7��e^�gi�LA�^��i��F�b�})�4��1�l�w�����
Ƴ�#��aa��K���hG���b�����mp�}!1����V:�$�6����'贑���i�k޶�I!ٳ��,ԗ�s�mR8�mD��ݿ���1��>N��o�ۃ�}��g]G_�����z���'ML>ފ�
�w�(1�Q*���8�9�~�8�򉗞��o��t\�o&���F�����/�R��p�~���?�|��_XV{u�i���-	��VF���7m^��Q���_²���ҥ`�r9�pВW�"�9�ӣ�r��4����?�?���y|<��EZ�S�GpI_ɢ����1�����ߒ��y�i��MU���M?;ɴt�`9=)�E)���/��g�\��&՛�溹n.�>��"���c��أϿ�#����_{����y8�ba���+�Y���sX�x��^uO>9B�l�<�����TX�O9?�5_����_x�)�m^�_N��҅C�&m��2�3Ʈ�tZ�O��껙~�_%ռ���:���C�����O=������NO߿�Be���<+�7�K���ڭ0[�WV1t��\�@���*�d`��
-�f_���R��ၝv�1�6�l����8	w�����}'�9-�H�`�X��?q#c��4BX �aP��*+���/]?�M2����j�B�=��2XH�cgK8�����<��y����KH�C��jOEx�hP���Ѣ�Ó�g��JپW�`�@���7mf\�����Gt�������ԙ�ZvR���hi3����R$��F��w� �j�vDCUD�َ�`3�a��n7i3.wǠh&Q��ƴ���3�t� ;��0^L�<�`�l�  '��q�!`4�O�9��,q�067�w������ ��3rs�h+�g��G���_dw��I�z鿰��C�:�u�W�=�3��`���3��1�9EԒؑ�VqA�����I�Gh�,��w1��k<�
�$�o3�[���"�U.;O-��Q�1g1���G��*Q�0�q�0=�=�n���G�9$����`� �]콥꽛F �Xa�-��Nq���j�B��F�&�W� wb���>�����}ܱ��d��=��?�Y���P	ώ��싈'�6�5�g��ɪ
�j-��w�t�U�<�st�� u1Z�����k��k&���h|k�3b�� h��9ۍ��.���i��X�IϢo�]F6��H�A慜`�Ma=�m�����J�N����$�g����j�oի(���|��O\�[��ubj(�nV�E�lz�K��է���ɿKb�����m^�C�l�C@s���FNf�w��R���11�0|ú	ƅ��ˏ?��'l�!ZQ|�  �p��Gd�}�m�ό�lD�@�)��m4�W �y!�eO��MW�r�&��ae'����$$�pŗ!h�z��h=�)��yN�݅���|1oݵ�m\/��:/ſdz�����B�ͥ�ctk4 މ�j��^�G��w� zl�@�nǣz�J����p(;�`L�v����� A}v�c�X���% �x��~ԗބ� ��zlҵ0}��\�>K\������j��ћ��r>$t�� ���X���[��_�V�ΘN"��i#�؞��wƧH#���a��j�I�X5`� �u��bxΥ'���_�Y�Qށ`����r8O��ӱl>���~��6�_�NB��i_`e�|��0v���9�B��������a�=\J��i8�Ur�9�6CzF�c��"�'�Cس~z�����U����ZQ"���_���X�r�����_��e:�)O�YJ�E�:3�����e���o1��|W���_��g�q<�z�rZJ>��s�����ǯ<|�\���YNWSI��9�ӯG[��ˉ%����.��_^}�q�]K��N��ɡ�˕NӲ�uq�����߾s��r8<�ps�\7�����O X����w����Ͼ���_��������+�)MOʜZ^*�]/��;_���e6��|��w�6�H�pP֥g����>x�������צ|��2����Y0� -B^ϓ��9��+M���)��C*��ue�����AX��Z�G����̏|�����{��뷯���<M��Y�f��&u
�j�I.���:;J���n��]k�1ąu�|^)��s�Ty��0����Ad6���C�`e��FO��x���B�6%hq���3�xN�N;g(�e�zEh��f,p �b���8�ѹ��^��S5hBF��(u�NƵP�M��Pb�Ks��`|R=�؍"^�dg�Ìq5pX,��#)-�"�G��:��Y��ʞ�MV)fL0��gV�U;� ���"Mwp��N���S ��]ܶ~qZg���c���qϞh��Sh��o�Z�W»�s�
����x3Ћ���$9[�M3���\֟$�����v#��Ҟ�e2:g�Q$4$��2,N���p�;�wt��cw-Z�W�f���_�q0a&�,q�(�~DǄ�Q���c'�$��?�C� ^^6w���x-hJ�����A"Q �[r8�o���KV��3p~�7�)��$?E����{�@�b�{��3^��x;�ϊ_�љY
���_�U�(����%&�-td������&ȃ;ug(��1�|%g�W�{���W{cO�F*���qώ�/p�p�G\i	�p�)d��X{w�u�"w?z�"���6�>I�R���w�҂���$zڵ�äJ�K;G7I�Ш�oJP�*a����>B�����|���㽽�"A�~�/h�?��T[6=�b�����d����rA&��u.Nr�pG�_m�0���_j7���Q^���]��w�T��ڱ���F����'C'���_�������;B�w��1Q��1�#=+��fb}0�&��BǺ�e�!���ù�&c���T��g�f�Ș��%m�:��.�6��3�AY��C���x��z��}��WG���yw���J���DkK�ms��M���L�&
h+B���'㱞�|š����ٸ��󕑇�{�S�v-��!���n+8�Q���1(���A��f�c��g�d����6���X�"��XǠ#i�m����,�2�;��e����nķa*�Y���z��>md�ϝy'6#�@�1���#O2ȡA�6�ծ^1�`�a���B��Q��U�"I@����1�q��2�p�$�:
g$���픂Mk�����:�2��@]li���#�ߵ��@Oq�~�|
��'1�v0wk�����[Y?Kj"^r�2���h�n[�T�Gs��F�o���0�%
�\�xab���o4���w�<y��\ ��(����!�����
��
-��>'�U�/J��K_���4����b��Wj�Y
����7�0�	6���}ݚ>'@��/>)�{
��+�;���X�r�`�����m�z4�q���X���(������ DH��̦�t��ܾ��<���%�ê��I�i�P{�~� ?���p|s��h���eAZ��iY�|Zj]�\O�~���4��r�n�����o��\�wV�,0�#L&T�m˥��S���.oKz��
�*�/s� �J��_��������?��!�7��/]\�)�1��溹n��˯�4 ��,Kz������[��o��+_����i��[�j���{� 8D}s�ǒ����>#���.Az<�)�P *���ة�������=}���;o�B�{�2=�^
F��e�Q�?[m�C���	�4������3ym/��N��
�G���>��=��}�$郳��g�p��ô͵����۩R���r��\M���Kl ��MPH���K�B;�pV_���	CQ���G<��H�q�Q��9�M�&k��l��JKa�lqc���,ok�7ߚ5�l��MJ;2�X:�ĔV���GVn������f�W�c�Z����<�ӍSD.0	��E�E�$y�6H����%cE���X�]��%���$(i�?C��}���\8I!��I�����_�4i0��~�&%�f�HX_���D
��,��9a��0-�@�T+S?4g���A������ke����P��|w#�q�Ǆ�ᮨ��c9�t�Îr�ǃ}|y��@. ��J�<�"��z��k���x"��t$�6#�s��u�0S`�`//�X��F�Ԝ�i�]�e4f�g����Q?�f���u��`֝1�!oI>̛�^-�+�PL�NĂ48P0����u���������� w�}	��3�;�|����!1vf�k�(�n{�u�n`��aU٩�t�A�`����&�^y�qo��� �gp^�	`�!�8��2�рS�����+^��$�g��j@�9���U���;�����,_����#�&#�}W��K����\(IYog��xU0����y¹�� �!g�Fh�$o��XO��q���ݰ,�Wݭ�r��8^3ȁH���A0O����B8�sZ�{��y܋����;��;°/��ys�+�� 	���/
xt	�`lF���v�=oSؔ�u��&��p�Μ���&�#�X�<�sdgl�c�;�IѠt#H%�lQYP�pY!C���ɘ���k�}�1��G��Ϊ�#��AЗ��H]i�S�;vu�:o��Ytfg��0|i\�'�r{sAk���8$z������4l�oK�c���e�W$����G7�g�o$_�M@>�K�5���\���-1ݖm��7y*>V�{h�9:H�����hs�,i���o��K|�F\D�wHf�砵��ݘ'<>�Sw/�=+J#�L�&���<��d�}l�Cd%�A�b�ˉ���w���#���hK��ڕ=�y!�7	ӄ��z3~�rO�ݨ��M���4Puݫ���0ځ��v�(�b�b���{��b��h���m}�|C��L�l�OR��j5$̜ws5�<��Ie�	ҫͮ���C�b~��z��:��-�����lH @��=�6Ui|k}Ð��Ɠ����~�>�S/>�d��mii�xk߁I ¿���M�4���K�5�L���t��7V����w����!�ek�dA"� �$]�}J�Ot�nD>�d���f��oN�0S��ч���);˃�
q	����4L�ePHn'z�<%i9x����,��Wtr��,�F���)�gƵ�'8x[�����Ogpc��NYo����;?o��tbԮ�������W��䳟��r~�,5Ir�I9wE��eK�X`��.|��U�X���b랅e�i�������+��;2]<L��s���tu��](���$i��#��A.�I�Z�Ω�w�N+�������>;-gr�w�+?��o�7�1�w���T ��n���^u �$�����;o�o���{W/�N�t5���8}��{��T���4�E(dE��gVU����Jz�4��$z����=|����& �����:c���� fS�懨�}��o&5�~�{��9_�)=y��O?��?���U|�����AUK�5�m�C9�BZ3���r|�*
�� �uS�ŕ;��v�Z\<���r��0��fII��Z�Y��{q�3�W�A=NS�N�e�����f���)����ˢ�35�hJ��Ol��Ex��`%l��iƼ>�;���a1���ߌ�b?>�$f��s��<�&;wD��2:���<���M��|���v��q�vQ��亨�
�A7,0��3;DwK��ʹ�5��Eܑ���|�c��ynx�ϣe�k�����H�9l��#0w�=>VWB뉌�h `
uoD��Χu�Vg���z'*��&���eQ�h1�@vu�
�LE����˘Ao{�⹳�� �D񙣜��.s��n�aǝ�y�g�	4h�y��t��11�Mj7���~i�� �pfG�$1�қ�������?��lp�� $6؝uK7�c������^�a��9�ـ�$��� ��/Z"b���,Gp��~{��h:f3�����ob���RrI!�p�Сt�����ш�a] 8�uǈ�lF[�_{��Pc	k �������lk�GI0�d Qj�r,}'%p϶2"b�Е�ٚ��+��5)_�]��P#�W��L��Y��"^9E�d6|�D��a	4-)!�Lb�C�)�<��'C�d-�)�8$G�a)Hmg������J�^��iL�}K�P�"��x�g����~�s����SsrI���-�x@�+CW.$����v���l��J0%���O�勏U�� {���|a{YCa&
C1|A�y�W�N08�:��F�
�� ?�� �p7g�V��%�r�gb����-7�w�U�c��g��j���E���1Jq3�%���>��^v�=�W�[��wH���]�g�@m��D�VޮP�'w9D�k�2Ϸ�n���|��v}g�ub�)�´�>/��.�WQrƯ�XM�е��\QY^�[f:d��p�U�*
�Oy	�n�������eTá�@�>Omd�?��%!G�J�����u3�Cq��~���~f��������C��2�m-�ﾶwњ���c�v�b�8J����m5��p�-��y��=��<���l���v6�6_��;s`�h�D#~�C��NJ�P'��ͧ���ְ�Pu#K0u�o;��s��E�p oX��+|��6���rl�u�$�|'�������B9�m8�:���T>r��|X�������5ł�f?%�C��la�1zL�e#	��e�l�:��]@�hyӶ5MG1\.���w�w�5 ����'J��v�����~�v�6=6���ڸ��0��;����ԢT�/fб��:������r��J�������0N[[�'O��bɔ����@{����w���[l@i�ӡ���ٟ���E[��r6. ���9����1���|��I[��uf�E���͕��|�-������UwYԮk��p>_��{q.�pR�񺏮ϡ�o�@����|��~�U�k����G>����c xS�Oh�(�x�~aq�:��4٧V���iz���߻�ܣ�^���[��&(m%e�Kb^.*߻�+�����A.�A�kB�7n®��L�sS9/�izz���R��\ǁ���q�\7��us���' 蕦�iz�צ�;����ߒJ�`'R�SŮ�����;�� �r�K�����a7��|���ǫ"�h}潳����g��R��?��O���?�3�{O����f��-��TN������/n]-r�DE�5�S�`|)K�m'P�V�ݞ��+�h�j�\A3�dut&̙�bʣ?�F���V���<��宴���P0���چ����t��E	�7;��S��_G������#�Ae�@�eŞ�
A�3F[b~E��Ď;�����](`�bU\�+���:���d
��N\k&{�璷�W����RLr���@�9�Pܡx��QF��{��S-�bm���}�l�>I�'�pԈ��`��b(�:���[�%�w	s*n��^��p���ٍ03V�T�	eh�c~�F��߆G4.��N�58�F78�^x���F����j��cx��% ��&�+��Q-����jc�g��" ӯ���&P��0�!!l�J	���e��dk��d�&�[ؗ?>�(i����A�y=�e�F�#�e�v�		����]��(<� �p4�;�����9rf�	Y��ODަP��l�$�/�Y�d��'&p�L%�s��j:&sv+�mN���!`�AV�.�aIȇE��#z������{���c!pU��gYK�b�X;����3%�h���]E˔Ѭ�QH�,� ���I1��wDi�f  w���(���q>�sD�՝��L�I�b�������6�t��Ha� ୯�;C#�- �9�0O"1��&�i���pƓͩV�����ڎ�}>�CN[��/2�X|w��QQ8D��ع�	�0�1�8p�l58@�����L�Kǋ�7�(�<��q\��˟;�c'�(3��@Sºw8�0I(��m��|r�~����]	�v��/f8`I�'��w�w���m�MyAn!A���tQE|���:���e����f �^G_O�V����Ei ��G��gaf	}�TE@�E�Ʀƅj$��V��������/��[i������m�dK�S��gߴ��0ƥBO�M��L�e�Cîq��w�մK�
c��H6X0�Ħk���v�b^�-�b���i�7��X����lOA��f��c18�Ŝ���N[��Yk�R����Q��U�?;�`]��dn
����<����$/q޾�I�ˎ~2D+�3�P�:�P���ѹ.]Y }܃�m��6��S��<U����ݺXBJ��79䁹�V����,�R�}�����M�׵��h�|���Ksd��a㺉/	�=�q�;,]<
�x��X�A�u��
���>��k����n+��^�~��#a_�e0�8�m#EZ��ek��k�#�f�����2�Ge���As9�	>�������'�����+̫�+꒨��:��췤O̍x�����dU�
�"���P/��&B�t�<jS��x��
�Ϫ�5�G;d�Aa"=މ����Y+�j�E���n��+}�T0F����U,Iz�g-���P۶���k>��?t���qR�������
�F�����:�:l�pG�x��h�����h��\j�V��z<12��E�=c"b�����IΎ����E�#S/�����#)d�������a=�ؼ�v��_s �6�'�t���W^}����s�t(���b���Q�=�P�9��|P͖��7�4��L�Y��g�ǋy�r5�����j9֣n���溹~���' �=���_������Χ��W���|�6��� �ۜ��/���=$7�+Z%�P2�%2S�_~�姫��*8jfԕ���<���G�)~����2|?�75�Xr��������sϿt��׾7���-��ɔ��c҅���c.V!{����~sJ�d
2v3<��%�*f�BIa��� �*Ky(upB!�h��1�k�k����e�p��\��9����0��8��K	J{�@��&�M3�آ==�ͱ�p���!}�A���+��(sq��,�9[Ȉ�]h�8��rk��mP�G"\��҇�Y��,���mZ99�D��g�!1@}��`Rz�{��ۻe�����q�`���+�v�D~Ș�2�!\7����tM�*�p$�^�N-�ធ;@�a��{�ؿ�i�s�%����A'[v�����`#���J���[t��qTع����O��:M����a�^w1C ڀCeXg~D_�~�8�����Y|��'�hWȱ�
 ���mT�86��n�g�?�8\]-�[$#/��u?�F�7g�^t��ڮ9����x<�8 <&tTK�U���"s9�5�D�1
R��N�+͡������X�og1����ݓ����m�4�q��v<pXc7��d�>� o.1���ީ9_�'6�XMl��>g���w�a<���������4X8��+�~F���R�y���� x"a�����F���H�;+]�aY�8L,Xݏ��u��<'r��k�HDl�08e��6�,�򠕿Niv�4��ŭ�w�Y�9�Y��nwP>�єܝ��@��;ҩL6*�BU�#8�c�PĞc��i4����:����&���c�y���d�EV�A&��xLb���.�ŝ�� a���8���8���?��)��s����5?�Y�>N�c�m �q,ߍ������ï1�g�;Й�(�!�p�þA�1 ������k֝���3��k�X��Cbae�׌�z;8>*���T�5�A=T85��w@��w��oC�,q>�W�
WǾ��R�� �2��N$T"�s��P�q*-�¾V ���/�-67��T�U�p�=�n��x���MH��H����tȠ���)�!&@���M���y���A��n��l�n��\����v�ⶋ�& �pRYO| ��/</���q�D���f0�=����3>�?#M>�ڳa�pc�2��M����= �	��S��v�+��(2&��`+�&t	j?d�5���a�>� ��Y���,�i��Gۀ���*�6a6�x�M�o�s�k�{m��+���00E?���J��P�����v�-9�f �B�?6n`��$*�8���5~$�=x���������
�n�A����V��J�=|��8�E�P����O�Q-�2m��?�H���c<#H]�P�i��#R)�/mƝlӜ����.��|YJH�M�/���R���������n&�}�w� )ڱ '�����Bu�mf�k�J�G�5~񢏿k-aT�[����D-g�4Q�D�D\�����h��� ��{(-��ҷ�g��� 	��9<+޻����2�K;?B�/�4���\I��>���:�Uu��1�yx�$�o��|K����X�ؘ�+�f�j��b����Ƴ>��ξ����޽�{'���q�k��n�������#M (�b~t:����?�ԟ���Ͼ7=yp��i�^���j;���ȩW��+�<?Z�����CMW((��������E�*Ж��~e���e�Hۄ�8�v�sR ��p���Q�|�{+�n	�<��{w^��Y }~���eʖ^��)���_��kV���M�E�f�d;��BUp�3g^�!AF�;Al��ô�x;��Ѧ.6���&���u��4kjW/�_E̙j�Km�.(n�(j�T���d';�}��ƛ�I�)6'7��A^�m�~�d[�V>�Q��$�}C o�S����Z�a3�4+����?��b�0	 ��l��d�F�*�)�,y8���)3�R^� M��u�4�{Υ���%��0��V���攆���ZA:�4���0o��H�ptG{t�WS���0�?3l'׬��5��6��D���A����q$��}��Y�K��xu�i���1\�]i���Ė���c>��V�/�\	;B�m�vT��sT(�*�����-Z��w~u��ϋ,f�&[@��q��K<ۚ� �
ϊ�nH�/�<\�3�p��܉N\�=���s�J��R,L���������Ì�bF%֯9X1��Ju���_��祶��ؑ�qR�l�[��A�E6w�#�$P@͈���U'���UĠ�;��*�x0=���`$*'��@&�#�sx,��%C,%7��P�_WXad����sYy�<�*�����t8�/Db��]g�9�9"b���QQ��m��"�\-�גT5fՇ$��������,ɪ2̟烝?�� 9���z��JQ�����yAe��V�}���8��)�I���5"כ$Q�'�a�)� t�q����6ƍ*��t�4{9���`��"���D5X'Ъ�Sٓ�bkO����b��7���/еh�Y��"%�/;=��::����Qz��tis����Q3Ϸd������K��I(�{T�tL�M��.�cԑ��ƛ��`�G"ܗȓ��9�'�����*�zyr�S�@�гd� C�1��٦��@sp��$��F�~�ĕ�;���KWຜ�wP��Z���o�X�G���g��vvL��Ex"�֟5�td�b��>�x��7iW+�:�zt}�I\�*%b,����.�˅9S����~�7�x�F��C�E��M�1Q�1��з1�w��U��1$:�\�fkC��dUl7�D�$��;M��y�MF�o҅\.�9�n��9�����j4�9�ǁĳ��yOV��DnS�΁4?�)I��m\݆�Ğ^�*��g~��J���2�׷/���4kx�#�p���f..�9��0���gC�s���A�O2:V�P:/�3$_��Qj��i.�	�E	��b�"���L(�f(����!�/�tO�k��Kb��Z��|DQ�ι��}@/Q|[�6L��+u�B� �K�gq�'���ӈ�(�3!yt�%�W�℉���'_w[)�& �	xN������0�{���suÝȃ�-B�B[??���캞�y�ʠ
oDio:��nT@'��GԷP���9�B$�l��W�8��2�&�q�XB���3ʪ�غ���͆
���T���D�"ns%��f��B��#��̯�<cY���&��ӂ�K�<F�"��(c�4�`���̚�;�&���.�tW��F�:�w��C��ЯLVu�v���51�4{����C���]�F���M'Z�ތ�	[��N�ۿ�CB  y�c�B��ȁ�����[�O��b����z��@��{o�'��V�:�t�Ya���T�t�4u<�u�I��� ��T޹�����������������~������;w���]7��us�\�룮 P9�ٟ����������]�)_����_d��O-��vOSTnV�w�{yw��*��8@�p��gk�ْ��g�����U�)5�掌�������;��O�K{�Bm��GA�£�5�y���*��㭋y:�/s;Sin�V!Z�̺$�T,*-���g5j��S��3�#����� t�Z��+�����S�;{K�:�����"L�E�u����Gfb�n=�E�	 ��4+2"D��V��g¸��'���!�����q̙�u���Efd�q�������f��%�yX���ܡn��U]�n��m6,7($�� [6`H0d�Mzl�4��LڰLY�	RS��H6��s�w:g��;3���\�Rz)?�Uu��g�r��9"#1�$�ţu|��̽k\�^:N3�#�1W3���]�PXð��y��y���+����.��S���<G�g��@�����.T�e\mޑ:7�| KZb'j�$���"��q<cm�G	$�67l��JF���@t��N�Ew���@s������Ab�NU֪h�m�{��c|>r�܌�5���Vb<�� z��l8��<�b�V�eIk@+��Aw�Uyg��R�G����m��9a&�i���qZΚ�fbW��J�E�PrY��3�`������k�PY��n���(^F�]r��~*���U�`lV����p�[ �{�U�X�V���R�t�O�O�ʌG�X���zI�1K�8˱��<��J��uA���'�{�ь�	_6"�-eh����0�H~	��x0�r��1Y|���H��ώq�����Q#�����]Dow��:�g�,�Y8Lr�+~`��D��',��p4f����-�gЙʭNqZ��I���i	z�x-���=��/���!�����s� ����|ҍOb
�ǀ߉<�#L���x�d��Ƒ=c� �ޔʳ��?_�.2��8	��E�F���2g�-�G$* �NpR�e咿xqW{�K�$��Qx_�2�e �^�t+1����9�-�/F� yn����:� @���� �]��O^����^��*��:�W꡾~t������fҴ�fЧ�,>�жq����m��7k�e���|��P��B����+���+�$�P���ۇ(Jp�8�IV.'WY��Z�+u�ΎJ"��������;<K�>L�yZ-�.��U�-<8�Z�<x7�[�XAO�vd=pb���cX*����\M�Ph���f�- m)9*�};���}N@	/!�u��	S`��~��z c���7_"A����PI0�d�Ŗ�7��c2E�G�/SB��Y��c���O���.u�f���V͚�e NcΡ���w9z,��V��m �j����K�v��-��0)��
�8�1��6ǬhC�<L���X8~������O��&mW�3�u���$�J��F���5�>a������~���{Nt:�Q��&@4��>�Ͷ�\��Oz����!���;�)�٨V`�k�ϖxt��Ñ|4���(�"�)���"�c=��yt���y��v���D>����Z� ���&��f�ԟ�����m�t#�Q���&�C=��.�u\ϵ�Lc(�6������G���t��nzi���9�G�2����з�F8����.~cޅ���\����vcObӪ�'�c���p�e��G��^KYT{*�ͱ���* �=���KQG&E�w��k϶`�z�iYn·rh�
�jA��mϯ�
��15�i���{��6p���wk9�vy�ts���w>�+���_��;�~����o|����K_��Y����u�_r}�	 ���������̞}��޾gv~�x���E�5�Ul,�4$^c���\׆R_TPـ늂�<�{77G1C(n�����I GW�ۻ���|8�H���E�L?�.��'����xx����R��9�u�Τ,3C���ޕ���q62]m)���%++�b>KDާ"�ǆ��R[)H�����0���Et�p|vA���1f�^X1��$2U�2H1� ���8��f󬥩2�N�T�SKk��)�Q���6�c#&Jꇑ�sd
�i����	1���p�Q�"�橰�27g �pR/%ϣp�a,�;�|�]�!%"L:Z8(
a8�#�@<S#���\��U|:s1(�Փ�k$���C�,E�X8mP�$_p�Y����U6����R@���4A� ~C܎*�a�S
��܎\a����k�h��.x��dv������Ny��N	<W�6���(����׵���cC�e����s�t=`Tؒ����$��`*�8J��}�J��L�8�}-k����	���q<j���3:&	�AB�L.��=�
#�,��oq��-lU'�����7��ư����:!^g<#��mYx�����{s0��;��pכrRI|�%��&X/Y�b�`�O�68�:�՘���ٿ4��%�B��$�8�9�$����Qg~f��k��4���^L�qZe�>�CA ���p>xE���Z���Q6r�ո/	�����vhA��gr.���BO��J��Z���t��a=����a�|��6��Vt/P�����3�kok���P�tx�L�fL���9�,46,h�}�j�q���p��W��6K��t"��~/�I��3;���I鱯��Ƿ:�"P/텃8`���\L"����<b�:p�*e��548.3oٕM��{*��8�A���^B7G�l5�l�|�����0�R�I
��Gя�k3���˯��Q+��y�|����A� h^y��W�z�a�eL�E�XI"�/�A�V�L�kU��Ѷ���@�����<7C`��]�	WJ�n��fLրTS���pQ�p=�_����*�E�)`��������82	繏 ´����+~ZV�&ҫ�����f(t�s)��c�T����9"0{#�d�$٪E��o��v����L�]��@���ի�*�2Fo��֢���؀�26��s�V� �/'�B��wZ��;,��d]^�&���J:���Q52��,�F?��D59���c�H�6f<�d� Ƽ���/If2���>;�+pA+�c��L2�_1�<���5s߸���MH���'��+ݫ=vU�U	���똲��+Y蓞D{��Z-3�m8J�~�ڗ���G��\I6DE�����)�0��zCI�s,��:�Ы�������	L��_$��z�3���
KI�����\�ϕ񂬁��N��1yCHӋ�S�G�	��ڑ�tT�+f��BE7����I���N�z�&'a���ͤ������P�c���J{� �
6��,��u����|�%Y�ck�PpB�ό�́8Y��˜�+������� �h�2�ۅ�i"���X���0�t�x
�����^���D��jе}�~,��B������{}�:�8`�p�Ej��߿���֎��˽�Xon_/7�o}���7��嵇��Yq���u�_q}�	 �����㷎7�psao�ҏ�]�4$����(L;��]�C9h�r�.�+G{sA�{��h��/w���J�����v��xv��dzL��D�[2s"�^�D.�����˶�a�v1�[��Ÿ�S��!6Bd͡�y���(^K0�i �Ұ�b��J�'̨�h��k�/�ɩ�c�C@�jP�w������gI��U�s#lT�we���	'�R�5@��[X�45Q�11��к:`�ʹ��@P��߂�	�k<�+u�¹j�5��\���n��1��o�y���R5�⊋:���:��ꤐ&��4K�';���o(�R��綰��������k���Wh�Z�p����珣�*g���G*,�wg(�k�0J��Tv��=�Q�̅g�^�I�h�߭�!JT*���J�d0讖���@|�Ns��s�`� 0�CcH�Sl �m�M�^Tep���b=��J$(��d���i�]a b��C|�8���\����րI)�{j���8�D��&�V�g |�r�u �H[t�X����ԁ�@B�Q�縗���F�xI�t)y�H�C/��Y�|��G�ℶ��j؁|G��H�}�ϛTm ^NhP}f&i�lt \%������<�����tA��Ԅ˱���8L*�_�K��:�b�.��G$���:�O�Y�[�#���L6�,x��"����2~���\���0��?}�Q/H��RW¯=�u>jC�Z��>��ݢ��v��1��N�p�`����@M}Yt"��7f�z?cN�>��T����;ʕ�.A���qȋ�3���=���U�x�ώ�p~]���gݙ��&�F��J&�zT+s�Q�s[���;h�
��x�p��
����0�/�S��4�ߑ�[%�M�1d�H�7!R�o����ν`ږ����3���c��-J�\-��K6��|-x���YWȰݘ�Y����gp��xIt�5�ڼ��?ڟ聺P�#׫#j�O�x���+�>�&�%���R�q<��Bg2��I����-<ߩ��j�L~�q�	�h��@���T���� x�e���Ӟ�84�|-A1��Q7�����Ug 4d$�X��X�	��B���9%�x5(����.�a/m.t��
��sI��P���vsny�O�ā�0+�o�L�\�Q�	�`U\8}��g�'������6� ��1���-�8�O5Y'�K��7�U-�TB?�1*_(�!�|H�uf��)�?��N��,c;5s�zDe�c	���
�k�Ak٧�|a/P�?��J2e/U���:MrOX _����xU�A�����-�c��SҀ�Jxw��-�N�
O����m�4.����u2lsU��ψ�n�����Y採�����*�&�������ǗK�(֬���:�C`^��fH��/�7Cz�bN�	��3}����ϲ�P\�P��.���k[B7�������W�Ǜ�mA_%�>���}fW���:7#ϋ����**&��?�:`���j��t!�m<��#�~6�te�}@��|qi\>��k�Lhp�<q��#����\�_Q��=����j�zG|�6&�b�x��h�)2Y��<_��t��~_� Ķz(�K����m�߱�� �ڱ~��ӏGZ\65�A���fC���8Q��ʃ�[o|~��O|%��u�_��+�O=�b�ׯ|�'ϟ}����Ϗ�/��`ֳ�;�� �&�.%$I递�l�B�>xz7/��|��l����ߍ�@�#�G�)�S���~�V`N  �U�3�k�
�,��u9��ڡ1C���9.NWW���-��q���F%n�d8U�9�>��p���@C�7�Ѐ�n��w�U�ƾX���S♡�㈦0�"P'n�Y+M��\���Q�.�b�t��Ju�z��p׌ a�ř�fj �nc�xZbI�N&��
 c*R�g�<�"��� ���uN5t$�m�&6�&��k[$�7�Aུ��`���8>�N�O�$χvc�;���8�4:���4�ͨ�->�D�kB+>t��9z�H!h���Ǝ2��XuPN��S�?�N�_I��w��;�^�D1	����Tݩ��
�`b	��[��N�T1���<��'�۶���XO��\I�-�g�-�a�c
��\}�Vc^����#+x�v%!;Ф�_e[��E��g�����jpO�Ap����g L�g�c�ӧ gU�T�~��û�S}L��Tm%���R3���)�,<0�q���(Wh2h8V�"��N�by�1�|�d���J��d�3��S���n��(m��,V����J���4�ZA�3O�y�Ly���X�=�Z<�p�絏F���X��"r���n�m���y���⨂7A_�9����(�i��4���ck�k�K����0��\�|�L���_ݐ�I�:E�6x���ՠJB.����8��\�{R�$L`@]|��Y7P�|��j���z���h:�2�Uqϡ��l�eMp�x��x��0*.��MY�1U�I�!���1tovȍ2�a�x��;�*O֝���3�� .m����}P��ߐ�fĽ�u��W�y���>�s���~��W�J�h@ �ݨ���u�Y<�\�R�&���8�1X	f��c���Z_�k2l�@]	'���x��n D N��ܡ�Od�,{8������� '(��ɜ���_m	�a1/ڴ������H8�l��?��=�!0AK�8v�Nc;t)�{��Q?����2]���t����'�?�8�jr��)�`����tX�-J����8���a��o�� �2m��A��d��}Y�sS7:W��2��qyΦ��^��X	"x�_��c�����*�4��o�/p!!�Lf=1<�]��R��qF:6��W�Q�;��<c:B�Z{"Cֲ�B��A�?1���jG�B21�W�SY���ZF����Z2�J�#;Dw�X�M��;Ah������]�+�+�|d1����"ɂ�I�ye]�o��W�&��<�Yֆ��ypך����K��Ʉ��`����W����eE�.*[�zl4�iR*��%��S���c��D���|��Xc��>�Bi�d+*�,�{��~���o�G�:U}�iM���"��Ba���S��6ܿ黣��##ⲑ�"R1��?�X�J��w2G�'�O__�1���&��$�mO��XQt��6>N��=�,���胔y�sT�:M�>_P �d�q�q���s��<nt;l�̘�H��z�ʞ0P���ų�/OTٝ�vcN��D�|��� �^���l�F{�UF�����+vn�>=�
^cԁ��vd\%��t��+\๽v����]o�'�z�h}�ݟ������_���u��� �w�y��T�'?��������{q����s��V�u���k�XN���|ar��:,C	�R��� �6�/�,��^kkY�]���r��|�4��"�\l?�xӘ������$�B P����c�,�~�gNP�m�<ߊ�n�Z�q;��틧�jwKUn���f��{k�a-���k��Q�	�v�B0wq0�*2#�1�	巢T�1:��"�	�۳(�x�vH��C�&pWܷ����1*�s[��N���C.b;EL�NC(�=p%'�n�*J ڨ�o(�CY(�����8^��4�}VpL\�СI�i	���j ���H)p���,0Ɨb8�K�p�4���#Dێ%5-ƿ��e��v��&�@Q�>�k��1Yo�!�4ShxFB��$���e@ f�eYR/�>֫�����c�t���5����ѝ�q$g>��Vc7�ɸd�kM��8�~���GW���+�7�}r��u
gnp��d;�#�:���,���ݜ>�/�� �:=����#��q%��;�t@�k��+��7���8�#4f�����<�k�Ј)��� �$&F�'���p�#><�^�"�9!���/h��)T���n��>�R�\��L)��^�`t|-ń��\|�W0+!.$�޺�W����r�|�
$;�Cw9���ټ,�؝y�}�m�x���`,.�tHNz�ė6����p ��
�-Fg�L��i��vfؓjͥ��{�Q�s{see
��N���N c̋x�j:Vw2��s�JC�ޝ�Ĺ��׋� ���e�%X#�s���oTs ��`��v���O�3ҭ$��YiW/8��#p�W�|t#}�	����4x_���Ƀ�W��!�F���[!��^.9z]D���ѷAd�ү�i$�X��y0�`�-)�w��T�S�L}V�	�Y����'MNc����|��jhy(�!�Ϡ߂���mVA���sŔ�!��3�u;F*/��[�I>�$�!7��M&�p�p�z���۱�Y�8B@so�]��m�V�("կ�/z;����|H� ��K�ͤ�ۡ:�j�x�u���/�o�R�����#9�?�XDsz����x�����&x���	��
�O[�C����1��E�~8B"L����&}�>z�2��E�X9r�I�H]n��*��Mb���'�{��e���+�wTr�o���u<��zÆD=Cp\��h�Α|�����"!U�F4»�
����8���Ʈ��r;�`�+�*	nK��|d�X���SgtAR!�N��e�.�.�zt�q�;�<��F���T緵�:�73>��4�,ǐ������&�=���Z�<��Cb7�?�����J�d�2���\��$Q��	���نu�� )2d���x��L�}�ɵ�+3nW������%a�����j���=j��k���9�/C8�A��|a�#�U@��u�\����|y_q������2�R`V���;��v~�s�v��H��v`g�m<�/J���I
�=�
��ClJ�gK����<�R>n�����T�t�V���&���䷋-D	<���e|U�,�q��L�Y����ӛ��_�y���괿�s2+�����{_�₤�|�p��Q���M1��*�X]��u�gL``U�/V;��
���\LZVvV����vw���;]�}�+.(����|#�����������]}��N�]S��)���3�� `�KT�d���6/��2�	�T���P7�9/���e9�K=_��w�-}b���������y�p���R����^���n��÷����} �����f/������gO�<��x<~� _���u�_��t}�	 ]<|�|��������������/o���rZ��Z6glp�Q0]x�i�B�����Q�r��9^~��my�ɇ����������x�p�&��Yb�wc���'M��o.L�% �M��ޮ%d����_z�ǋ�v�ֻ�O>��YA�>�2�(��v��̸J%�ɽXOvWƹ1��:ډr��4�O�����"J���)q~��I5���Ii�G���/?+��{�l'iK������c��T���� G���gxZc���xm�N��Ayu(;p��_�<���M)h��Y��'|�C�r�0=�aS�4�LD��F5tSZ�\�c���p�EV�Y8�tW�[����b`.��XY�Jx�"A��1�a�R�����c�W�Wk�`��g�&����4��!�]���N�0��~W�B��+��ƺ`� �y aAK���B_�;�L����V���i�t�,�ω�� �ɤ#��u(�%2�YuD�8Qd�$�a�=�Op��N��΂� ����4��`�c:��gc������Qv|�1�'�ugq�����1�ݙ�[�+p2��-Nz5v%�M���Ⱥ y�_��1;t��� �3x�VV}�B�`�}8���`MC��@�h��Ҧs�"��i��q��?E��᜔�	/�R*O:V`,e8�*�ȋ\@�$��=�bwRl�v*��\n�UL�Db�����O��k������p� A1��'O�ũb��;c�&�c�c�ݐˋg�o���g�'N���y�&:��F��V�`Ц�Wdj}�`��ղ� ��<�@IN��D���w37��t�"�i�׃kѽ��>��z���qE_ܭD��b��2���[9��D>��2��?��r���%�8Ԭ8��zD�bs���l��k�������O@�����`�����A�����$�d/��E��羆R����|�P��,]
��d��o
����������u�8d��l[}��e㝊�|��ߐX,���b�p=FP֜��?/�d��[�7`�!))��D$D����я�8�/e 9±�,�®�\��oEΔ�PaO&+Q�PAA��	�Er8����I@?�ܕgB�E��u��.ԓs\GK�V#�Ǥ���݆���'�%��N���'�V�=f\X���',:�x��s��J���u����3��sڒ-c� ��nA�YpG
�.fÖXp�r���� ���*�*���1^���j)(��F�[��/�-�ZO�6�W��W�/"��&t]��O�ʨĄ1`�;�\��W>�	��v�C���qq�(��}��=�y Β��k���Do��4��{j�p�����ɻ����E�'���Yճ�4 Ίr>�GM���s�e��qMu��~����1�Y���%�4��8�
G� lҷ�ZJ4�!:渷��,&r����.�)򔺉��2��kW��,���Q�"7���x���a�m\��
���z�&��|l�Pm��fʑI�&0,��Q�I�:�އ8�����_�q���څ�6���F��<~��h�=D��$gA�V�����A7eDr�W��,��c�Gm9�Fhg���s>/Ǚ�(�tL���x�[�P����=*�����"x�'(Ԓ�7D{��%H_�\��Ab�SK�c�!{�G>���W��Я(:��9����a�R��+HV?A�Z�".�ֳ�.?2�e9�H�P[�Z?֩���ɞ>��8�rt$�W��d��h���"�+n«w��J �mК�D@��!��㦏���V���q�C�n� _�&V%�S}����eș�m,Νξ�N����=�yr�o~��<��O~��c)=:��٣G��_���u�ק� �2�:�~a?<>����o��'��[{�����?#I����X�"�g>�.ۤZ��>����ɐ�M9����}������l[yR�����c �\�u��L���E�\g�t-���%��������������=�����m^��b8��Yͭ,܁]n-��n�o��p���j(?���a�/�<��M�TU��s����k�>�S  ��IDAT8��	�@�|5���Q��ѳ��ln�s�`�ʧ^[(ScF%}������.8�Y�K����9�k��ۍ0�^�J�RhQ�"sF#�YLC�uJ9��8	��>Ъ`�1U࣭q���l�&�r�XrlT\�����������ٶ9� �u �Ї�ȝ*�J9a��R�)M©V�~#��5�.�jQ��p��VΡ����*�u��~��=��{��wxu�8��B�0h�c/§hH�`07�SK>�n�"� ��3�+��x�������ZG;0Y���loߑR=�ZM�|.���Sύ��b�V��>J����l|���g�3���qW���	�\�t�ȚB��YYG:�-pv� �m��2*�p����̍4Ч:���+��hȃ&�.�w��Ay~�p��!eB�pڄ�g|�]IK��ŲS�"}�,(�υf�(�s���Dӛ;K���rc���r���2_!ﮑ�D��{��N���2�*�:��H��:���:�z���J:���b���
ǘ��h���(އ<��O{������0�jIFc�����2�����<$����Zp>��[*�W�Vf�\X�s���5�R'i@ǕbJ\��T�,�!��ܬ��c�w�t����]G�3�'Wa�����R�/zv�W���k1��C�8�p�c������B��nJx�ۃ��I�u?��o���VW�K'�e���Y�ꃵ'�D~��Q�k�B�qē�Pe�c<����	L�F�����x��$"��@c���I8�ˈS���K�!�8-Y�Rcު��\Eac1y������nr��*�"�#ncH��衱l��#݇No	Τ��\d�0߬1>���D���s���L�s��ܪHp0�PAd>���7L�G �\b��#*�H�ۈ�.y-B�pK��<|�W踄~�T�$�0[f�4��3�\T�Fa��6粃ݬ���ݖx$�5�?��	�9���C�~[B��5`���̃�:0;^�4U�q9���;dH��e_9��v�fG���t�u�x�e3�J�-쇁J�R�7���3��y�����a;Ǹ�6я�3b>&���Ȃa�h�7u�8:� �rKu1�K��k�7X�.���y@w�Q�6[U�H��(_�l\Ӏu�i�l^�h�M;(�d��S�)��|�|H�[x��q�=��>*���	?�l����/�e.6O"�dc��6��aIi����ץυbn\��r�<�j�]=�M�6�0q�i�vhh��0TK�y���~��q�&��({���J8O�o$��nF]&f�6(/�D'wRu(�M!C�=ʦ��>T�{A��?�NWe�8՛��8]~�#�T��ۀ,ı�����r{���w/Kiq�Vwi��Y��9v��"��E�ύ!�g����������%:\P⦖�������p����G��ac,�`8R�8\�u��w=ab��y��8fEǺ�a}��[/�ͯ��on��g>�'O^ZlV�������z}� ̓ n�?8��7������ك�
�/�F�LXFڗ��8,v�Q���8�9��a�Z-˷�����>�����x|�|��x��Rc�g��}0������E6�����y��.p�����x�̓���?zx{��A��.������&��8�S��M��v�	 ���u+����:�ʅ%��;�8p֯�"�G�:-�zr:�U��f�jp89��� PE��X��"x��1�N���PS���"�%'�YS��I(?i��vc����]��s� �b�C���P2�7S	BU�^����+i�f�2q���(쪼�V�߳�Š���<�kN�t&���j���F`H?�O��0�p\,r�A8H	G�� \�Ъ�s��a�]����U�j	�ɀ�2�,3�_���0F�B�auX� o(�<j.�c�t����GY�4L���6������lj�������H����<��� �C��"]֠������q��!U1[�nZSu�Lc��ZZpzs��F��׼� ���g���KI�؈�+��xDc,��X����@k̓��`5�{K�y�h	Ҥ!��XL/���\��QA���-�/:�ɿ|>8ך�Ԙt7T�p��| ��F�
X9�,\��T��,�VOL���\���\�D����yS��_�r�AZ��qL���-�����+%��2����&9W�?��#HΛ�w-���G/	t*�o5��m�� �������ί"��JxbG����c�|�48Dn&�!��f���X=q+�J{whŁ�s��M��X�7�.�ޯ~�,w�n�g,�T������������Lu��[7�Q��\@�<Z��*����r����+4�V&�HǷ�)E~�ϋ�1�u�c��~jwdM"A0�q��ɦ�@7���5�ަ�M��q�;����m��c�8�";����a�*��(w_5�@�o�G�?�׼���
�i�}%<4���:s���wQY�p�D�j*�zp2��n�8'���@y��_;��R��`;dl1]���\ך��`cB�_G��9���;�Y��`��:���}��"<<�T�}�s@	rV�&�� ��=*r��9�)��q��-�M��<.�X���t�e��P�3����?�S���D�f�Jߝ	R��A�:j��[J�rujw�)�&���Ì�=���������h���z'����\�y	N^�Wy�i^J�����Kz<@0��^)r�/fZ��@���$օUJ�Nw�'=e�n�k;z�V��2�?L�.��8��'��ð�yH8�<�mr�0U�Z2睽��<Cc��V C�c�� 8��������d*�{�T�hc�H�˶�¶:��T德[��#Y.1&�Ր+�d�w;�|c�bJ^qd��n��H�� 3����f�x.��H�pj!�'�g�7�:ք�q�q������{�q�eA+�0\?l�j�9��pL���W��V��2��'�V-li̫�>�V8�≴=�ry�����v���1�ho�{�7��z���Y��o�K��O���f-0����n4	`���r5 ��	 �"	@��+�vk���@j��\�ܛ�|~��~��VO��7Eax���ri�|����N-� ���Av�r�G;�\Ϗ<|~³��x�c�+1���u�_r}�	 -W�O���o?����ӏۛm��*���㟖 �K�_�z���ܸ�G�lCP8��ȋ}TO?y���������˲}�����Ǟ���4v8��Z2�x���~�Z��~C�>��8 A2�A@�1�^��/B��w��/�ެ�U ���<ä9����.���e�w�!|r��;���]�ݙؕ��TJ��=݁32ՏO!��,٨kQ�b�OY����櫌m�Ӎ��R��\q��`�Q�����ss�.P���ew�TdW��h�ʮx�]	߼Q���;�D�u����^�h�Q�֠$��`���F�s8�By��{�c8�	��h��aUԽW��R�7$j.G��m�seÁ;�Y�2��v��$i<z�C�?��l���f^����P���)��I	iI�:��	#�q�����Sc7u�xA�0��9CP���=����(��Q� �@�?_�]����U�6#-���>j�g��8�����H��W��.���N�BX���](AM#e��1"�;gw�x��xe`�M/W�Ї��߸��Z���f�犀�;��3+܂�I;R�>�_cM�'灛�����\O4���@.��No��Xc,W~��'�R f��P4�}���ܛٴ3�����"ڀS}V��z'dV�̇"���wF�\F�:��Y#�3�96�c���'gD��!���<���uP�4���Z㘓%`�󹱎�=)���A_�+�ȳq&��KL������|��e!4�Ę�p�.�->���[����P[Xm$;���ܾ��f^'$}R�Z�Z$N9��6�����k�\	y�k6R����rC��i��.��<�;%�m1��:A��������F �5�����6if���%Y�)�N�l�y�&�D�A����x�I�J8aC�2�
�;�p�:��C�1�.JI8������j�àӦ�Qy`�b�V3́{
]�t�z�Ob+F3��D䣲z2�0��Ļt���7��k�aH����L���L�5V8o���[^�8�F���rM�c���*]K�q�謻�^T�c��!�q�k?r�(����Ȱ��J·2����#qDU�$�Ï@�X���(7�cGu>�-l���g�>��#b�=�r���FT�O�X��Xv�iTG�%�9+�r���8�d�;�����NُJA�hޅ���u	<��gw���i�/�����Mx����ծc(OD��[ȲƆ��H�	�G^E|1盕�D{�k2�	�t�`c�n0C����$��{N�Wh��|�f�`��h_x��.5*iʃ7:t��?�e[cFU0�wK�DR�o�dB	x'�YE���y���?՛�<
D����H���:\F�G_q��3*U�n���ia���h4�����pל޼��+l�����~��տVN��w���c>v �X�=�����9I ��?���2tg�<�53�e�0�xA5p�S�,K-�I�x��H$��A�I��dN1G�b����>�M8��A��'���h&���d����6�Iണ�28�Eu���_Gg��Bت&<���p��R��B��A��a҉8����obܢ#UK:�8�@I�W�#Qj��&}A�э,�CUb�$V�D������m��J�x�ds�t��i�z����G����S_�K}�X�vxtj���]�n�<��M�A,4πW)];�1�`�bӗ����?�������˰�]L�'=`_S��2-��*Q���e��ȄF�+��e���͏:���
��֛���7v�f��u�_����SO h�[|����������n_���8�C:��np��]��������[K�ZB�C����6[;����������~��_��o|��(�9.7�;�죛��ձ1y$ ���á���PF:�bQ�N��$ <7�& ��xQ\$���x�<{�ѓ�}�O��.e��4[���P��0��B?}��������Nh�Jɂ��a�QAr���m �Y�m,TR����\��F�A�;��&�\��,�ee5��Q a�Vîb�J����T�%�ϒ<N u���XY��@ʲձ�(cԼ&��guJ�����y�T�,�ە)韆�[�NAQ�e��j(�b���q�@���qJ�b���b	m���r�+�3X���9H`���q��J:��n�R|}G�@�� K�u,C|�i�6M�<�:o	F�8�H����E��,p⮄�����(x��g�Bc��s�s�f~"2i'��%�"PW|g�	�%���T�+z�=�.x�gU�%^B#5h ���a�ZN���U���_�|:��e�IVb]bgA�aNICE�F'���;��5�d�u��p-*q��'�>���yY�(����opdg�m�6��¾ ��[�=Z���D'�:T��1��0�Y~�H�g�s�QuS�	v���|6c@�8���o�Jx�� :�av��:dn��6v��x�Ƌ�ڄ3����x��p҆,ӆ�Ͳ7�SF��o�%X���8�y��j(hy�99�����X��N��.8ݠ$�Q6�>�$���B�d��5�/E��P�>1:I;��?���b���v���W�e�:���u�����R����<6Ii�[�ڄ����
�
@��5�k�;/�S��6	��<7�YE���5&lEAa6��N+�I�`�]r �F���}2�+����)��n��,e\"0�̀s�w��#��Y~/  y''.��n���FȌf�6��H��Hr�'d��"r6�W��*��R��v#�W����n��w�V*�V.�4��a.�vUNt�	��WK���'&^�hk��������R�Ȥ��,X�:��>ϴF�x��"h�E@p��q&�׼�Íh�v�tL��	�)���Ůd���3�:�B9Y<)q�����֩U*�ʐ�V^x��%�@��פ�,Y�ݚ
m�o��9j[Bg�s�)��L���_@r_�n�)�ka7D5 m�,賀�$��:�G���$�
עm���Q*��I��X�J}h��U�yԒ���lP� �L/�:���g��3�����'L�^��&[,�
~��84H��}@��-XSa���%�re�y U~i3�k�n&UN��~�W���=����Rwq��5]�m��5�f�c���u���	8��χ�[b�%��H��'vM��?����(�5�$�Y�'&[<�2�A�U��	Ҫ�	���y�ш�k�c{e!�`2G�2䵔#H�#�����m�v�N��
�o�"v��p\�y)jǫja��b���z�.	=��\v	h��>,��K,i�1�rH����5_/��û�mB�*#� ���G+�ɮ	XHv�&
�m�K�D��#���P{V�=`=����A���xmGoU;��|�[���O.}�ԋ�S)<�SV-�|M Άx�l�
Q@F��.�'cj����_�����Q��'��oz��:�̩�.���.,Ώm�7Gg�
w�i-�{r@;L�������������~�ڹ<���}�������ק� PGjj+���?��_�����?����g�=��y��n� wWhF����{//����K{�^�8(���3AY?��^oO�Ow���v���������G��|��?+���e�8 �@0�]��A�_�k��� G0��"	��h%�v!���"�4��o'�&0^��7켾��?��7_���Q���zޖ�#�ƾs�0���0 ���j	4A���mvS�L�R―����U�lTы`mv�� e-Y�2 QEi�vE��)��N�4�Pr�늌���qg�8-u�XI�i�1�����E��P0���u�Iq���&���@�@W$+���ndV�l���F����Df���EQ����|B��/�3���s@[��� �,QF%��	j�
�(UXG7f�����g���F��g�'#�Z�S��0���ն4i��G)��� 1<�����^�]P���h�rH2�,a$_�7&���q%���R���p�Ď���Y�_�ÿt�1�p�@�{��db�?�~�*3�;�]�+��k��N2Gއ2?_<�s�}�B�$�8CpBoapV��d�93�W�����G"p�/70��
:y���S��!\������9��G��`�dAQ�ǭn��q3.p9&ܖ>9w.¯�=�s�Ga'kV���MG������ٽ���c�L��>�Jr��҈�#��,�P$9ёⴺ�$vR�O���q8�_/Ox��e�D�޵�T�*#A�����I�w�.���l�eg��~D�`<�`���0J�<I�+�7\��8������D> (�&}'��;�å�G/�>�u�D�*j�nK�D����i�f~��B���n�c�gC��
�w{����9�O�=�(a�w3O��EQ?�냏!�%�i���C��	�cI�/�Kxڃ�A�f�̰���.���dD�Q�%d	*j�Z��l�n�9�?
�m���F߹�G����	�x�פ�W]�rc.�-hk�vtx�#�.��e���N=�c�5�NK)�A�4�DG����g1�H�<��B��]�c�y�hkҁ1&�L�h#��$��#����ˁ%ω���N(0v�� ���:���*Lc�uϤ7E`�	IVL�\�ER��L��|��}�i�B�"M����!�c�AXJ*U�S��|>hw���Wc�F�F��E��1ꜮN�a灛�$��i1�����K�G.��X�~�ë�6䮮Q�a�ȧOԱi�G��M���4�|�h��t�F�%�	<,��pq�)��hdz;v	+�y��'?J���rr���<}R��S�9�3�ou#H�>��#pl|�K;��>^t/v���]�I�	�L�FqL8P�Y�h���'��y;P�-�XyD���(��������mVJ�q���K=Ou�	Ѭa�*��:�.X+�H�J��z:��R�	&����>x�;��"r��a_���~0Ǐ���|����7����v��_i��j�aR����mۤ礿�:��+�mFn�f{�lw4	گk�W���������]����$Q� �c�lcs��VK�/}Ф��в�{%���S�U}��s^7�s�	�+ϲo��ܹ��G��=;������ϵ'��8ʄ6�UY�:�G=�������|�/�;����_4�r�PMV�r��P��,�u�����T�,`ݪ>?"�z����ww����o����a}�tww3�Q-�ˍ{�<�_鵪�/��9���;?��ڹ���W��m y���������������/����>�����^{���깔��������Ӯ И�����������xR�vk��l-%��JZm%���؄F�"@~��#���Gvw^����0M���R7�'t��Nϖۗˣo�����_���8��/
������1%@�����R��"s��v�_�=�|~i#	�ֿ?�|��0��Bi�?k]�:�O�}�����/��f�nn��p8ŧQu%��=a��!�<���;-C�m�_�<�^K��ݡg,r�o�"�QUL����<�AMC����B���ٕ���1�蛶���w���K��N���wo�e��<C���r�(֝�I٧!\�}��ER��X�Q�A���Q�~5c������X#n���<��+��,��:|������� ��y,p�d%|2@�ʪG 4��1��R� V��P�W��N��xB���^���E,��{�S�1Qz���Zái�F��u�ٷ	^4v@�B�f�,�ə!^��9kGOX�R��T:��Xrdx����[�5���'d����P���k� 3 m�Q.���ŝ)ju��N�{>�v�=��`$tP��%�9�ɡn��F���ü��%���OɊ�������[\&;<	����X)2�l�N��=��
x�g����k�]�_]���^�i�����.���x#~�mT�I���4���_�T���>T�u�Z���aN0��a�xkO^d2��N�(m_��.?�]v�涺�~�q��z�:��_�6�����z";�y�	>o��b���3t���H|�G��|����|��s���D�Lw�b<;>}m�����e��{�4θF^��d]���ީ������.D�5�̓��*E�a>Σ�ܙ��d Mi��<��ҌA����qT`t޿G"DU��������/Yo���ǣ�V+�N|�N�����Iu#$��SY8��e������F"��ʌG�a.��cwzv��|G}��,���pW=ԛZV��I/��^���.P(��D�ca'�L��aօ�V���x1��C�B���?��Ky>�������U��V��$����\�2��D�_����&�|�ꋣm|�n��d<�F�i&��ׇ8��V�#|�R�CQ��� 9A��X�'t��q���eR_{��qt؍�ٮp�g;NW�r%��*s>qݾ@`DiJ<zk4H��w%�w���u����qx"/������A(�<Z��>�d�����9�?z�3�~���j���H�o��kK�Հ��_Jz!�iM' ���5y�8&� <�Z�&`�WVt $��J�2D�f�ę"�_�U 	�ܜ�S��1�
3�����R��|���4�#ʧ`�l5�2���PN��6�C�!���tjKk8�G�DBq
�)2����8�D�O>�
x��'�Y< 9���֐ �;�w�;�W����e�����#��`��^ٯ]EP��@���w���|w���e,yZU�#Dk$�l8�_6�������JTM���	/�/h[���8͠�^;�P��Gb@��-�'�0덪kQ���x�!�;|�o��I4>Y��>�-����w�Uo�`�_�_RyMJ�M��K�#����&+v����e��>�w=����`��'q�Hbp:,k� �z[~�7���S_��ʛǷk�Y\�f�� �F�(&R�o�����*ת�7&�xO?���m7u�����w���?|��?��g����U:6�#OD8?���ǖ@si����Kw?>=���
��T�rZh��6���7���}�Ư������s?��׾���2������ק� �C{�ۿ�O^޾��j�������*�]�/`FJ�݌̖��`?��{vC5`�B!�~aH���mg񹟛���>�������?~�K_����̓�m�dY��I ���G�[�����.���ϣ	�G�N� �O;6 U 4  P [�[;w`;�~���el�������{��������R��f�0x�>��6ҋl��x�%�	g�\4���I���aL���Ē\��%�ͨ�P�)��	0+�eVN�\u��31�㜬2��q�*�+��Jgؙ%Ei�_�%�^�Ġ�8�G�ĝ3�U�k��f��C�I�ݼ���]�Q�����e[P�������Q,��9�dd������6>/mT]���V&�`W_]��R\�]b��*���q�L~v�}�X#:�~x(᙭�>�?�~@�p�0��~uh�s�f�7�w?�¨�8}HA�\���(��Q���v;���I%B�W����}��"AH�`�����o�J�$�E�(%���:'>���m��Z.:��"�`DI�ㆆ1n�����=y��������͠��(��Ef�J�r�9*���4v1�I#������Y��8��{�v$�C�y��D?�0ֱ�nr"��9֧�������:n!ab�$���*� K6'�ˣr���h���"�����������u�͖鎴����N��9��T�[hpO�+�J�<��� �Nc���nl+��c#�w�2�y�é�m�k{J� ���M@U�,x���幬A�_eY�Ѳ�#������`�K��1	~�� 	��,�x@��
�7%ڃ�U��b_��#QC��݌� �@�	�t^C+V�r���"�eφ�F���"����Hv(�yX�Ow�ę��n�ag��اb>���z2����*�,�'N�}���Ωݏ
���r��8�E_��M���U�Vv�wN��q��[�mF�Y�e�is��F��`~��I�-�"�ɭ����ح�0�S���j���K�B�>w�
��Ҵ~�)4I_�i��e�w"�S��!�bR�/Z�Ih��x�� ǃd�1�Q.v��f�����$!����
g���2��%��=E�
8PC�Y��A����s�l<hn�h��tǷ.O	��� 0>���� <>s0�{���R:���2��H�)1�6���<y���2�u��jR��׆�@�ϒ�#� 9�����]:�Q!X�Q����"�?��۶H� ��h���1�عN&��R�b|;��IF���g{�����6���c&k1�\��H��0�	1)�\�N���3�}�))�X������NK���Z9���|�P1��mlT8�[�~���Y��gi׶���'U=_qE 5>U���p�)}���>�Å�,�`�c�.*l�0�yV%}`�Y��2�bΐF��H�p��rE��C�7�#����:ٚ��.��N]��0!B?���㥣c�W]yD[�k�g��R`w�4:f��*��V�#p��㝬cm��굤;mQ�%ڰ�*ݖPvU"`��L��W����<�a�W��ű
�SG�~?`�ML�
H�-ڄҴ�c��X=�_�r��x���xw���O>�/���=���'3m�/���Q	���5�b��Z�������7��w?����c��;�>���r���앨�<Mt��hm�~��lw�m���R���~����K��;��Vo?cum���_=	o��2�e�<f�f�������nZ��O�����^^f:��m^=��]uT?c�ީ�����q+���{��t:=~���}��u�_���' ���ߛo?>o������ai�hn�v������ο��&�����NO��؃��ˍ�x�nl�C7��R��(�����VN=p�|�7�'7O?X���������7�ڗϥ|r<^,���|��
C �0K��-��EԸհm�[e��aQ	 	 CS��g�a �rs��Ѻ�?����?��������gm���w7-_�\�τ�֝�S�'ݡ���v����~���wO�{�����]�[A�`�Qep8��n������qpVW1"7Q\i���m*m��R�p�m.�j^��Y��HA�����3����q��*�T����:��[E������Ǯ=8q&e���O�p�r��F�j�G�Y�1�a�B��mv%U��˸q�*��
��s��[G����0�"����0O	�O��aW�Po6G�(]��HF�'�c�ẆY��jPV]�t{���t�U�!���s= 4�q��c�8Q�A��n�ˁ�>��
��{u48���;bT ��
A!�vL�pd��i$������2��$�N��x\a����\֪�a�D�1X9bH�!�]��k�N��(Ơ��F��X9�83����>��V�����N�3�b��\$I8ށg�����|���@ܘV�mLIZƳ^8�Ҏ�jS�>v��%>Ơk�W5`��<����� x�c�A�m-�L�ǅ�����Bw�p�!�6�[x��@��
:�,h�a�k�H�ټX�&fi�*����5��t�W �#��>���.tV����3����{����'��3�
��>�~�r��QxBJ����]�/�i�o�|hu��퀵wGU���R��<,<��� �Ǖm�9�s�7	��ٰv�+���H~��)�i,�� ob�W�Pu&�a�@w�B�Wog���^H%U)�5��O�k�C{]���.�;�G�	�Á_�z����U�jVùI�>��A� �ۈ����b�u�Q�$��Nȕ��gPK�j���6Ε�\��(C.��`�B��%*��`�1��w|����\�:܇C�v:�%�Ϫ,�Ɇ�u]P螈���J�~�5]�
��C.�&���I5x̠)?:I�<�kBh�ǱIޢ�≗��-=�/J���j�Kr�7Pw��\��ص�������@LK�Ρ}��p�/��Q�"ȅ��
�QF���D���Pͮ�����Hdٌ;��0�;��\t��e �4t{A����>F�7��(��\v�5Tb+�����<q�|�*͊a�~���5?��o�K��V��_�0��6+N�%��Τ'�S��!b~"o��H�h�,�<�� |)�b,�{�e����qT�� �-��)�G��¡��)L���l^���	�hC�,��2�g������5��*U����z�Q��S�3���z�&
S.�6��R����@?�:�|��qL(���~���_�
�7@���Ѓ�JP��L/U�=�F�C�]|HuzG�D	��O���R�~��r	�ؘ�v���5�D�W��A3�b����IȐ��Cg���ĝ��� �J�	�x;cM���)ƙhBnP/���x���G��%�<gqZ��J�&�^>�_(� ���y���
��|e�G��qՋ�q�qa�&����5��|=����ͦ�nu�=|~c�ʁr���!q�v��d��Uh�l��es��ru�@����o�u��96�;-xK�d1�8nn����@�a;E�
u4�-v��B�z��O��<���9%A������Xo�?׷�m3%�FI�esY���C5���x��gD�W[��z�g�;{��M�74=�%��.o^���Q�.-!����8d@�+ʳ��~�ח�~�k���y�r���Ͼ�8�P��$����z���#����}��CM��byyA��ˀN�����z��?�������w�^�~j�G�������v,7��Υ��e�7���\��g�վ{��^�K���|�]��8F�(k;~o�����������ϔ��z��������u�O;����;�_����~��^<�������Ӄc\�nsY5�Ӈ�PnX��M8�k_��O_>׾��܍���ͥ{c���E�r(���o�֯��ş���K_�]k����C��|>�$��X/"��m٠M4���"P�]���^u��Q��﹀iB��_��?SI������[u=�{w����?�{���}��u=��car���8��BE�eŕ��n/��}l/�㬘��P���̸erXj�� �m�7QVˠ(Ƴ��`���3WV��3�Ъ�P�����:�J��;v�����{��d܋'�>59D�PU`���_5>�Bb��	I��S�D���1��m�3��y\�G$��Ϋl�Q;]Tʳ[-�J����y�n�V���PN	ތ;�X�s���	KN�\f���n��*Y
��aiz��ZƎ�"K{I����^���ц��:`���1l��"Ϩ�����S�HW���	�+�1�]�d�0�" �h5��Иw����w7K\뾭�aLwFZ���i��s!�4���B%|�+%%�������@.��FX�sï�J�Iӥ�~���+���y��AS�7�s|؄'Ѳ~�59T�{N^�KO<�Is��D��䏐a��ݐD&0P"��ֶ�oׂ�9'��T�ByX�� (�^�:�zX�B'Lg����q���A������| x��.�$|�`�L
��p�Q{��-#�-�q�.��WBp�	0��s��qj��;�!&I�,����
�i8��-�o�����kiU�6�mA��>�\&�/���gǗ9)ib��/�_1�Q$�z�x�ӆ����5�Du,V���w��������0�!t�YOLs�^���Y�@J��j8�|0�o��`A}{�~��>#�aT�q�@�rǐ;17���8LJ��L�"�hĤ�A�7���oK�x������S��L~;:�u��v��!����/H����N�j����f��T2���^�6GO6\����9'tW!��ŨfE]��GE��1J-�RV֧Kv�_���p�v��_ѓ� yx�m?���IEn�<��N����!�=&1�_�1WE�p�u�y˰��ɹ~�����Nu��U����sC[+�)���5d�r�^��!�u�H���\�)�q�f�E4��J��q ?%��܈��e����̘\�X�<�Bm�}���X��0X��$λ,F�I������>���
�����̎Dm�	wJ�	f=������ɀmT��B��>�1W�b!�������]z�,c��z�$QP� R��4 ��X���P��^tLz����F��A�`%�"�:����N����I�..�O��Rd���N�T��[I�W�����/�<d�|�O\٧|�XJ�7�
��A�!������4`��>ͧ��̜& �`d���ſ�H�D��t-��V1��8+�Da�G��QQ�nd�A��?Y#���N�A��&;�m[t�k��=��|9���>�c�,6K�8󆖑kVx�d���쪄��%�E��P'��X^o��'�w?��O�潿.s6���4�#���o R���Ηj��t ���������,���֓66���Ҿ��c����g���m���cǸa�|�݋˖����t����O�W����u�8l�P��>w'�9�JP�¢���(�`�Fm1���-�r鼶���u��u�����3����������ݾu�����f��j�(C��ͪ�%�/����٩�%ڔ��4Ӑ������ ֛�����׿�W^���w?>�O���N����������' \~�������7�����?��?��S�g��Ƒ*���D�Eֿs��>Z���xQ�������d�x�e�����Z��i��������{���wn�����M)ϬI����jkk����$L�v�Z�L�R��+Hh��� 	 �[�����]�uO�v�Ȑ'���s������o��w����[��x\���͜Bu��k����gs��%G|T���?����:L)`v���3`��$�Pa��Y5�P���}+T��JA1�,j�q�29Y>b���]� R���ug�A��C��a�e����a��5��''_RWR=�\g�D�+K(�x9��]F�典K��LJ�8�ԑ&�>9}��@��.�����;�6vF�`��B�k&m��P�d�%��h8꥔C�I%��/���}��KODpՊ8�b��+�m�w�W�=v	��``�#Qw^U���$"���
F��Q:��U�(��s���������_B[�~jN�'940/�5� K'N�:� ��(��3��	8���(c^ �Xv�\�g�P�@45�Sc&�9� }W�w$���l�m�[u��A9
�/xQ��W�p��9�*?���h�q�y��}VUqg'��Qy+�U��ħ����0�j�u�\/�� ;���݀I�����	<���cR�����88��J�:�ҹw�b��NNY8Dc��B�>ם��C�+4X_���e��9Y�B�ѽGz	I%K/|h�De�J&�]y�8��A�=�^��x��/�X#�0ƀc<�Z/X[��29�9j ����υ�X��~ڍ�Y絬�W��m˻��5��g�N������k�+x^�~�nJ˲���{v!j�g�r��b������m̿1���0/�;T�412���|�#��B0���j|
�W���ۛsV�p���!:=��-Sųk�\1+% ���kO��^�/��ev�;�"����څz���4V�~G�ӟ`�D�+��׹f�!�?��ER0F��u���>��>p��x�r���Iֻ���N�We��~ʲ�,�g�@�,����*5B�֐��l�1��z�wl�=�\L���H��J����q��A���LИ^g� �r�*l��:9k�/�䲅~�+ex[��2��k�?��;d!��H]�b�O	�5E.�&|E�R4�i��Ѫ��=���L�;���A_L���AM	�e��*!�y�n��6���&,*��N��4�'�+��d�M�w��J����%�|�_F��g�y����+c�g��2;��]Mz��6��ޯ�ʳlWT|�/�]+rC��@����W�'�Ao�G��U>�i�X�GJ�l (:�[���c6+ UQf{�G�&،}�hw�v:+����PMh��$�xM�ER���,]7�������"�T�>��t~�N�]� ��D!�_��t�5�v�Q���뚒�Gw[~���񼼼�ڿ��w���'�ͫ4vJ
_���<	�����S9l�,��p���ן��x1\�s�|��Z"E�1іep������*S�"�k/���"��v6;�ϗ	ܽ�����������m}�����������hȐ�o���zq:i��f���d?�{aw�(�?��A�ll���z��H7��n�7�Ϳ��~`v��2��:��u�_��_p��� �.ˣ������W}������/n��_�CMΓք��~����ew�{�����g��/�om�u��D�3�>"�3�ZI���x��ǯ����w�����tz|Z�/�u}����&��f�y���?���ԫ�Ul�H"�Њ!���؀d�8 @`�x�A�̒I��,�؃��2��(�⸁��D5I�,YU��z���������ַַ�9�ʤ4�?���{��w�����k��n㪗k�O�>������͕a_h&�������D�� � K"u�\z�ϲ�[�{	Z���X�z���}��_������yyxs>l�-w���@i��O5l�V�������R�}�V�y�ah�(Ճ^��Y�tOO<�Ҫx\	�7�2�qֳ��ټ{�)�5�|!�KH�"'[���P�TW)�xB����
�at���G��2��E+Z�>�a/���2�ƕN^O3VW�T=������,K{0w<������'��{E�N�����ԧ��>�Ϋx�h�֪�T3�������!���StŜ�ͦ��&�4�!jA�Ο����)-+g_�c�e�LOV�1a�K��!)�9Ia6!m'�.���x3�j&M�_�u�}�C�&�C�]�V.ᤝ�S�A�#�I�A}ǚ:hː@F%���{�㏧�58�Nػl�X�v�H�6�x��F|����S�eT����6��;��$��p�y�x;wj�Q�6��'�_�d`(F�D3d�'c�r�%g$~�
 ���L|T](��tR_��;?�r��	��U\�ٌNlyKpѽ�.��#�9�7?:pv^�H���A���H�Q�0��u�@��`�W��$�IC����	�\s��@Zd�W���rl��ѯ�3%�`>�[66����<�;hW4��Ĳ8L2��&��,�Ե�JG�N^����{���=�=��#~��?&�����HI{`+B���RUB'�9�T���%5�E8΢�:�k���eWR�/'詊�����0n�[���uk����l�J�˧,�^Dxo�nw��@}�+  8���i%���U�)�e��"���W!cH�����%�� G���uB/�h�X�p�����dUd���9b=��yW��K0��b��nM�:6�x޾.�?
@�,\�b�f�����Fr�섣��J�X���p��k���K�$ϘkT�`�>��z��:���'�_Ҩδ �?]'��˜�D\�����fy��U�mZ�5uf���8�-��?ZoF��	Нr�wq�2� /4�mY�~c��� a$&�^�4f�E�*4��N@�$�<䙟�4:�˵b�#>�إ���<�W� �����Z��7�����B�=�mN@
�l�5��)��nI� ���������h{���#]����?Ę �b��~�d���>��;H��>$��N��Hc_l��O�_N�I�-��S�!�5�%����	��W�%�J�k�0��_�PL�t�e��&����rAP�i�~���I�;��Q��o w�!\�l:��$A	�2�3H��%tA�a��l�ScC���*��1.�E�<�d�C��\��&���ְ^`?/��A���r�T�V�9m�)�a,�^�_�5��O�a�&-�́Q�[]��&��~D��WL^��E�6�)�c	��_JU���ܨ�8�9G,��~:��z����C;�Gxw,��P���"}��i��O�c��~`�'������Sr��wɵڰ:��k6��w;�d%w�<���,7������!�u������۵E�ʲ��<-gu����_���������T�y��eS-���̓'�@��vp�U0+m��$�v���y���0�òܔ���Ï��ܯ�������׮��s���Y-S��*�nU�X+_�kҪڋm��������z���՟�I���<E���U�Qn=�o����G7Χ���oݺ�XrB��s�\?����& �b��my�����x���/|�����y�i�7?�����i
�ރ�E׿w�C��;���	Q���nn���I���&V�]�������/���o�����S�m�jR��i"�ֿ��?���Bz��@�J�� �04�DO��BrK`�-��󹴫;O/���o��k���7^^�r{�zz�L���,)�*�c��)~��Y޾�Q/C�u ��	�2����X#mz��*,��cr��ae�M�OZ<��b�U)T�+�uJ�x��C�����`^|ҝ��Pr��O��Q�Ja�'�w���߇���hX�A(���X)�>�6��o�P6O:}�_����h���o�N\8�����5�� ���B�2��I���-���{&�| ˆ=����q�����p�:j8��sX���S��h+vR`�	�1�;��Ltc�a���!	'�)�̌����^��MBa��:򪗬��aw�ބ���H8 x����.D�pjf5��?�%�dQ��
H��ʾ�5qY;A�=~w(#�h^Xx��#�V����O=08[�Uc����0N]�=���1_Hm�����W�PNcek+y�9�c!Z·��x�36%�b�Z���0I�߀�����|��K����I2��#@��"�D39��-t�	C~p���[����V�*�CE���_eK�W���M��*�'��x��x�}p^\�Cf�υ�b'�qgr�x�8��/v2���"��N���,��y�d�H�m���?���9�����僷O�Z��s�Y�>M�c�@1ه��<�ĢN�>�����@{�����r3����Y�:21nA�t�/Σ����A��b��@��%1[F� ThXJ�c�_�c?1����#�G��恲��-��%�������x�&��$!�֗�c��#��rGbٔp@�Ǆ��ŀmI�F���7��>�45u�BX�5K��X�Uo|�D�O�,��H����N}�/�넰ox�x%��t�̨�.�́=��
Y|ȼ�xH�/�`�8m�ZQ|.�m[F1�sge�8�����D����&�ܟ~l��w���1ܳ���yk�g��#�|�}%�:B�C@��G��D�����'����_�ؕ�A�&�j�p#1��9��G�����~���0g�@d�_�-�4i��?t��$6���:�"<�����DO�V�59m��Y���tƝ��<)$:ǥ9q��|�N��Y*�9��[�s��S<�9t�J�S@'B̬����$_�ݠM�9���y��3W�/B��(S����׻�ô���
��}kOz��j�[���y��l޷����#��}��[�g1��H��
�~���[5�3�S#H&��%d�r�?�mɤ;c�����|ΥXG%YŽG�IL4dfL۫��7��Lk,��\1�#�c�h�d�y}�׊���{�Wl,���p�$s���k�(^�Wwmh�ʑ" qy�^^�y�:����O�!%��fR&�|��hc�*��ɪ�v�L���4��}c�M���AD'����ǫ���b��GC/�k�����i\�������]�7|$_|�%����{"� 8�c������Kiӣ�7��Ϸ�|�+_m�v��k�j�inI*M��oX�_�و�<�c�R���,������Í��a�x���/�������}��g����/T���#YPv���/�����|��]�������nS�i��Ar��M�ު�����O^y��w�J�;M��C������s�\?���+ �g��s�{��ʒ>}��j�r��M�b�vٖ��Z4�sn߯�|����3����\}o[����	)�])ٜc[6�&@zP{�?�6�x����^�W��?���V�y���־���Ѵ2ԕ�^��=��:�U$oA��������	&*��aYVTΖe������ս�~���7~���������2/��xn-UH��y5����u�9����w���>��(�Rk1I�z�v����X�Ξ.D�@̆��cj��,�,s�9J�B��&�JqX� "�5�Q�vÓJۑ�S
�i��/rp)[6�l����T�b=�d��\�Y�ա�c�Gx(�b�aѕ�%GP
&ۆ#6�P1��Pi05�x���l�=Pa�wrdZd�{���NOD���d3ZK(���Q8ۼ9�)?mJ|��wpEBN�CSo4���yl�ii>2��^;��[(�	�1#�������ǒ�.���G����q\+�?K��`�pN	D{X��u��~��,i�GH򹤠B��O�y2�|��]�� w{��� 
ܥ��q#���G�l%��H��D{�YI%���mUڋ�4����,1�@���	�:>N�C	�b��hs��8��BF��!����ޥq
Y�ν��yw�и��גv���8?�i�恝�ω�Ёq
��g���|`�&JO��D��u�x��i	L?d����	8yOj��O�`�ؐ���m.���4L�>�#q�������
�l�����d �R��y���x>��3hY$J�x2� �P-0�m��+@n1m��@�X�� O)ء%p��P_��Ӎt���NΙ�0�]�za},4�pa�nI���>����{��5�n�8�lڌ�:�n8a�u�b&}�Q��|��T�S�w+�c5�1`��c������S�q.s�~-��C��FŁ$'H~���|��_�g�z���]H����[ȸ�(�3���K2��JO�t�$@|�r,K/���31��yy�s��a�#�d�@�
4W��+V�I?�ʵ��,��;�����:~	��[��G��k��X;��XK��Q��v��[ C�9�D���A��*%Š��JG$?�J����6m�5�>>�u�_σ��g�<���	���K�;�a�5�&�5p0)>��yz�������<���J�ڭ�q�K���do����p��Nr�N�l�N/��=�8��C�?�co|���8n����fa\�}�V����'���K���9�����X�H��2���"�%�?H��xc)��#�ւ�Q�G+kV�[0�/d��m��.W��s�?�1`�7����!k�n<�7����Uk���&3P���!i㥃?��=
��>7���1�'�y�m|@|G��^w��~���u����l:�A.��d%�����?L�A纗ڦ�ʗ�گx$>ٸ���Fr�t�LS�'8��)�a�S$ߪ�w)�����6�����1�ڃ�,�#�d���X�/��U���	�W�x� �u�D��-(w��V�{��F�c��!?G��>G�Ǆ&b<��!$���� ��\�64O^�'�1c{�(����2�X��xtL��cK{��U<�,�[�=9l�콎�����D~��cy�Wd2�������W8�~�vs;P�i�,e><\���~�W�o9�ȗ�ߩ����Tf=��:�Lv�!-N.���b<����f��l�j��r�r������Ʋ�o^�/�|��_���ʓo�|9?zi�7��ME�5�X�/d��KR��x��Ѣt?M�>�����߮��G?N����n���Ԫ����k�lr�������~���$�⣏v����?���ô�=�|\��g��\�W��nN�]���X��~"_~p_^�������ֺj�+^کe5��h���rx���������/��/�G7��3e>{����իU ,�T/]����ߍu^��T�L1Ӟ����l���~9�\�v{8�py�����?��������y~r�~���z�DK���4���)��u��dm�ͻo��6���~$�y� ���k
#�($�1��X(�*U��)�@7���d�yj��Б��'f��Z~�]�lB�@D%0t؃���J(��������mn��!��l��@6���WĝáES�rP���v�8�3�u,�e}���l9�M�ֱK�7�8�i;(-�J1��L�A��VR�adP	6�8\��D�欼�&x@��� ���e�:��򪑠!��ǡka��.¡���N;ƌ!6�b����W�Y��ɢ86�
�ë������j���C��ְw'�>����0	��N��&�8�
�$c'�+�<����`�_�Gy3�0tE��%h&u��52���!ˑ�����v�r�gӘB<h|��wM�8W�N7�����Oyt����`����|�<Fo�nc}^)P~��|����ۑ�	_��ΏA?&?�Y��w�����zrY���{��9K\y�����2����AF�~Pd��S��Nl��>cH�d<9�)��� 1R:��м`.��A#8�{�#��$��i-9�IB��:��u� @]���B�T�ǻ^P�@cr08&��8��`��)~����&*<�C
��O$t���'qw���(.f�VX7`�M� +î�]u�rBdK�7f�%PN$�i_��I��>���NG\�|�A߀~���4!"�b�4ˤW�/� �	�j��+��T��#�ͻ��Q)��2���I���b�[��9�XG�=���r�pݔ{�� f��/��or�r.�V�*W��U5���@�R�vN\����uiY.���]�:y��N��e��9�lx8��Sþ�h��]l5�.󼡇�� �`�	B�߽���]�ѐ�d;^�#iʾB�%��>��N��s�u`^��(��@]�'<�	���s�����D�aSl>P-r���2%�>~�a��~��y��u.��?��$M�c|ѓ�"�����Ӯ�����,6���"���l&v$��p�76�@s?�aq��h�}�a����w�'���
Z[K�ER�tD0uе��䓊��{#KT��4$t��#x'�����#;x8|�y�R�Z�0Nr؇��
�m��K��7��"�5�R���&��������^�[�4�i���XF��g1�uZ.?m�]�������v ��B>�v̏�p�=n�4������+�:^t.�$:8A��+Cր.Bg��I��sH�<�h׃���):��c��G���gYc�+��0W't�h_^1��t����c�;��� ت����T���� aa�
)
c�=���g1ܓA>�hw�<�����M}dY�!��s�^,���E���}$;?���.\[s�/:_�lZa��n��Z��-~�&��!�}Xy#���+��� $�i��.��7�<p������w?|_���+��USZ��?���5�!��z�ڔWeW.e:�M���_)��n�K��/�ŭ;2��_�:��ZrK�f��ג��~����g=��~�vz�6����adn����|1/����7�{��_�W����t9?�=/�E��>��LS�?�}m������:�~��Vj���%/�nӮ�����qp�m�a��վʽGʃ��Ϟ�����OHqU��ͺ~������ϧ� �T3���;����~�����_��d7������/���8QǼ��E�+�8U��Up��ҋ2�cWϷ�+-��r��b.��LJ��^�U �vu)�ᓋ��������������K�/��{����i�ޟv��e��<��4����g�:&�����b��*���7K[����/]]>z���~�?�Ư�Y.�ݪ�ӋY��َW�iޢ�.2��Ȝ;����a�}�D~��<�2sӠfs��B�O�<]{;�v�@얄��v�b�S��JϹ9����w\Fg8)�'�v��n_�q���ؕ2�G���ԫ�^S�mSzŌw� h�Q.,9�`ç�qwx�d���`��־z���h)��W�C������H���tN)YF/����>����pҟ�`P�X EK������՜���-���c$��]�3�B4�ϩm���P/;�~�d��D���/�jɧ�����0��I��J-�K��9au�U�z�/>y�:�v`<�rdk[�@T3����{�����>��m�d�'<,%�'y��C�e����������$��q���h���-#��i]�8,�p>h4F_��5,�}�%�����
#�>gWn�i����q��L������NN�(��[�%Rz�Z��ý�Wjk5�̻/�y��p�m�n�H@L���!'���0�C緩�)䅃E�k��;���q)��#';J�z��EI���A g�W�Mq�=i1���pRY�HācL�e�e��ޢ�ֹ<z8��*D�;�y!���W�|�E����x�@�/����Y���e7�}��z����;�Pi!;��ӎ�C)U$
�붐�/�YEt����(�%*)��Z��+�}��g[�8����9?+�!2K�AU
�Iޣ�2N�Fpm����Ő2�q���ر�#8��sT	4��6��<E���Ї�qeD$��y�!P7DZvLbΣcZ~41�g׻%�����g>���g��tx���X�@�]�(a��]>-�q�\G�<���dX�'����:�{����h ��T�
W�	����d��Y|��	  �����}�U��%�w�9Q�Cse(���;{	�L,��`4���0�,���<rh��[�2�p9������4�&�JzU8�(��Ĳm��H���@>�4�㨳�H��3�1�П�=�lf��Z-��c��Ӡ��:�c�8R���掸�?H�}��,ԁ���z0��l�H��3t�ܛ�$/Nc�����X^&�0dR�wH0x�5�7���c���F��rܸ��I=���x$�V��8���hɐ��uN ��'ػؕ�"��"Q!8��(�~O�Y�@�Z��
E~�O�uӋ��u$�8	�|n���o푃��4�f��&�%K��p��s\���쯏x��I�I�b^-�!��I��U�m����o}�2.T7[�b87��N9|V�{O!��'pI���H����ԦZ��.����=I~5[��G�\������c$����u�u܁!��_��X��~��$|*�-���a��	=���4
4��F���J���ޘȫ���X���k��+��r/�e���v�~��|%���]��?���Ԅ�m��*�A��=�� ~>� ���i�*a�ޓ:ݨ?|��w�}�����~�K�����M[���][a�N�;z�u�~��l�E�r����j�G�-�`��խe������n��~���~��ۻvyS�����|ř�����K�xծ���Am���s�o�ߛ�ܓ�w��¯�v&M��Z��Aa*�<�X��</eӡ-�����������߽usw��..�]����s�\?����Ӯ �����������W_~ W/\�\��e�δ)9{U�/FuϊZJ������wߒ��ϫ�iՕC�>w�myV�i��.`g5閫�e�w������<��o��կ��?���y����ޛ��R�'k�+姽4!4[KX����:�U�ܹ\����w�|�3����|��7�o�����@��k�vh���=���E� K�j�+?z�˷�}G��<��0M/�Q�k[�g@I�Na%DBQ���F��2bΩ��ﴷG����g9�|b'4��B��Cg���ы�@���]�}��1*ŒOt����N
������E�K���n8Ðt�S -0�	�[s��+�x6�X�� xE�B���1C�{�S�斍8�H2�pT�����DN�P�[�V�	��c�R�6��	'͌�[�]��˙�`_�>X�!m�(�[� ��+��6H��f����&"���qP���|��,�D�w��-�N�nP��-�w�4AIg��O�-;�`�o�7��8��-�&Sf8V�ά����`�D��I�,��(a' ��X*���hX	:NKд8ޙ%���d��$5��2(���`/7�� �V���m7�J�TKԙ�*������u>R�k~��$+۝�d�'�mӖ|Fy�������mA�i(�EkKDLw��Q����81!�����p�3E0�puQ��J�a�4�C�qHd�U�gC[�m?��g����@yJh
%�@Q��v[W_�4Kt,�$��S��fL_
�Q����z8v)m5�|��Ob�G�������������ז`�Wؘ#TK���� xn �l��F¤I�"q%��G����izl	�x	m�53�8OFB�0���hX^D�����B�:�b�j������&V�q��\װ�
|�Y�!�9:�u]tl�BIh#��'ܠ�d�Wϰ'��뷤%��8�O%������N��+~�oB����%v���WV�D[�.��I�_��������$끰��qa>E ����C��=W��V��$���I����|�ԯ���D��r���&]�����^m�/d%�N���Ce���A{E���y��aS��Х��1ۑ�^y�vBMO�϶��q��Nb��ೱ�����I���q�|��t�i巄�HV�+4��ʩuRR�_@ܳ�}ѓ�8[��X��#%�8*\��"IQ�Q�-w�<���̟�+�{��"#�[��']Ǳ�\��p��5��|��*8b-йu9��|�D�������/�7p�Hv�X�����N#�+d��}�|5�zqU�֠;2�ʕւCV'��&�I&&*^.| �o:�Ӄ$D$�;��08�Y@�²5HN;l$����U�I�`��8��D����-��b�#��1la��L�OD��aH?�Iƺ�IW1I�3�A(F��@�	�?�X���/�

=տ ƅ����w�4�����-�h~+�eS�S�䅽a|ՊKS�>�>����"�`�Ղ��ۍO���L����Ru�5������U��?�h⇒Z*q]��I�#���͒�$���4$ZE����+e1g� �d�N���$xk�w�Vm4�O�ã(Ǘ���X�����h�`�0��(��F;o��@�#������b�Jw�7N�F��«���l�M�H�n��4�ߚ�}2���Z�V��As����ځL�<\���1�Ս�϶���A%��>�8g�ʄ����i�ył�I}N���I^�j��|c��hj�{�W�"/���0=�J���^��$4;p��p��,�����dt(��\�7�Y��w>W�����_��O..n�:m���~���l͏�m�o�r�%������ɣ����o�~��z���Ƿo�����:촅��<�e�c��m��d =%Ď��ym�/��a�?����͝\�`�b�'ĵ�yq��egw�­�[��G�����?���w��+���o�zuKj8��s�\?��3�O=��w��_�מ{<]��o�_��psZ����a�+$�^���?¢��Ж��ȃ]�����싯��ݴ
���E��d�&`�V��s��/�-�1֥���̇�J��l����{�ۿ�����y������|��+�?�y���7..w����4wU�X�tL�r8{��ɭ�?y?z᭷���Çw����V[��U��6�ǲ�7������m�9��@�!�~��J�MfT�+��Br���{�~"ߙobV���֊� �Tq��H>����(a�)�p�Sĺ��Ȅ�E�\�����p
�4��r.�hkv� b.�-7,�V%��b撄fc�4��3Oj���Fu�Ӎn��c�4r&Ap#��f��Vw����]�5]LQ����pP� �0J<��Z� r�����@��2n���ʞFP;�a��[Yw��Q�m������L}�\�"�i�{�z����Ia���"����o󁮮�#9��H���0�O���Z��V�iYP��z�ꆁمp1�f���Co����0E�mUL5���]`��Qj�=�-�%���fp �k�y#E�`���`:�ѝ�Z
���	��mn<53�`d+�S�nF���i3��'u.k��0�zI���|��BP$�c�9���Lw<8j �>8	ǣÛ�%�������	�����*#�Ǣ�%8����wEv�ˎz8)w����1޽I��[jq���(�f �BX��W�+a��;�+̏��*p��Ck��E|�&+��'$��X���n!���9�:�o��k�
�{S�۔�����i��ʥ��@5��+��;l8�n�Ga�>��
<N�<^O�w��(@v ��
~ ��\"`�G�Vvo� �{!��㝕��i�EݦjA.YZ�Ti#����Dhv����B8(��{q�9�eٔ�R煒Ȁy����INx�8n�E�'#.�������N������8�j����� �JfJcs!��Z	���d�&�J8�
��Nԝ������	>Z��jb{�����i��Vë�����u����Z��dG��ѲX��=8�f]ԉizE1�39��K���=lq
}���!3�Ӱ:�_�|)!���q��H���T��H	9� R��m#�d4�"�����<��) ���^�NN�+�; V,9�TB���u��N�89G�hKؗT��f��.dt���
���ڤ�_���P�����c����64�z��f�,�Wu4/M����tlM��7׉ϊ�M��:����� %��\��t�/$N�K��B���(2u�Ȧ����M�����bƷ�m�.s�)�]���I>�D�)%�^s��f�M�+)��.<���P�����������`%�^��\���㉮���j�mZo����l���$�Ә�,�v��"�j� ( \�ݲѽ9�� ;�����f\�����D������E�dH��@�!i�i9�h�C��b���@�R��;�h0��'?���W�L��)-������q!m�i�����`����LW��讃�vD���h���>��g� {S�����S�{�i��K*���ɟy�`��3�5��a�d�6)1H'���8������3�-&�`��
��{]Q�c����mhg��ZO�n�!e8܂�ЛM>��鎗3���#�\��iA�����>�n.2����<�o�!t�jҠ���Zr�8�/���L��/-�}W2->���:�H�5�@I�U��5��(x��.�2�����NV(`�����1]$Ѣ`��f��m�>H]} ����O�v�f�H6�̔T��`֠��hqލ-�uK������!�H�ǭiR�iK���?v6�}/o�)�������%���șl��`�y�q����6�y���6�;le���?_��G��n�dz�P��7�7^x}��g>;��̗��_x~>?�1��_��4�+�粝	�rX��l���W��'���9{�\ܽ������R�m��=��[��uO6�oQ�����F#��eR�����w���U�Y]Ʌ|��ʛ�vr�;�پ��p��|,x2�^m����\֫��g�<����~��W_{対���`mYJa��~�������SO ���G��]���\�[��ۘy�[��Z��Q56�0ʊ
۹�1]��E~���_��]�rsEd36ٴ)~�fl4��t�ɲ����n�e�W���a���n.�_����W�~�K���o<����[O������t�vg=�lӰ.��NWO��]�n>}|�f���=�і���v�8Em�P�P�4�ɜ�ұ]oew�ʵ��x����û=��rٯk^B�0��Џ�Y�aD�"�����$������;�� gL����M)��(gZ�,V�ؒ1h�-6 �%���R������c���/m�9 ��P�`<U�8g8`����+�9��TCB�dp#� ���io���dK_�q,��E���lX��}8/\P"�IgQ�?By��DUN�x�6����?t84��=�;V��a�����Y����2V�p��-0i�}�p�����|���]����T7���phAQo��l���>8L�D�%c���L��#���ߺ�|�;}���.� �{Ӆ�e�_���Nᄮ5@�$��Lq���8��-XV�S�;Ƙ���WuH�[�Sw�Ų���5'IT� y���N�M}�U��T�na�2�7��j�o��e!���Rҽ��1��A�x����g
���h�,�0�hn������e?mm��/BF�����X����e8M���p�$�xek��7��'A0�����<�Ͱ�ɒPJ	:������%��û8�dSIN��7w2l�w���u��7(�	�>r�I�C�A��m��,�S��$=�G�x2K���¸}_f<Y����\/�u�8EӅ�C8�KjK'�����H� ��|�̃�#��Z�ұ�ݱ�N���[$d����@�_u_C�h�OZ��	�!�/�LP�R��Opf���A�6dr_	�(��5F?5݀u�����!'O^)�g5���\e�'4f�:�D ���-|�!���ڝ�,����B��=� o"�t����(f�]�z�G�ޚ���)zJ'st�gY��}��k��d~�8>��o����y~�CקWN @u���� �+�:&tDg��"=�[g�I�#��`XI|,����~]�\��eѸ1Z����=�Ԗ��h�h���m�Ziv�9�2�-��s?�?М��[W'p9V�	�-������|a�=���92�C	v����M�-�>MTΫw�8�J0�{���,���+%��'y�S2��)	��|r���<TP�y�@a��������*I_�]*^1U�y
��+X�k�|D�~ѡǏ��\� ���#���-$��TU�+$c�?X�A��HҞ�}[|ݒ{x{�R�r"� �7K�W�ϑ� ��>N��y�[�=���-�=��v��y=��Z�O�i� Â\�
f�؟L�����W��~��0_�8*�W�҇+��=X��4��^>�~#�`h�ɸ��<�Aߚ'�sJ,��I�Hz_h/<�GB�R5�X���b+8(���5tCd��� ��Xmk�c����K�y�<d���@K�}?~�c� d����� |�ˈH�`�m41�\N��͒t�օ���6�1|b�U�m	>^Ձ��uq�?��f`ܾ��(������H��s|xMO�� ��{i������^�Ϸ��o��X�y���^����UΖ��&����}�0ж��?�m�:u��/�<�e���>�>�䭥������r~�����\��l��/�t���ؼ����=~r_=�pj�G�y�:�b8�|X�^�ڬ�5T#���	u�H�WOo��-��>z9��~����Oȟ|��\����l��V�_,�ǭ0���[ۍ��e�s�1/��;�o���$�A�~�����9z>����*������_~����ǲ�\�h�M=��+f�ܻ=Ōj�-�-�	�|�}�"߻z$������W?�2�Y�v���th.&s���X-of'(�����	�-浔��v!e^{}r��p��ã�y�en���4QU�a��"d���Z�˴�����V� 糫��v�6+�z"D�m�nˈ�N��� ��F�˃��o�}S�.O�h��8���)�I�1%�4���Jo�j�d����J���dV!�C�f��__�<��HĆN�t�q�V�V��° L�̝D��㢹b��=0�v�����1(hJXܷ+���f�p>������<��Љd��֐��
m(�0=W��0b$^�;^�q���Yǉ�S�L��\��'���"��N8����T�:l��S	x�1���t��ýEVvֱCi?�,��	fc��v"`�37����P�H8�|�r����ؔ}O�0#${A�~��
������{ߠg���|�=h܏�!���m�;��A�e%�8�����=�-���H��ru")��� ��њ�����h�	W(���I��βw���)�xZNʊwN��>GbW-5�[�hZ"W!��Ō��>8mҋ�$�:�~��s��iM%��< ��fw�W����Z���f�Y�i� )4W�E��$�e')��sqR6��HhZ{E%�s|��֙��ދ�*gy�{jn�51A�O߃
�E�NȈpk�S���m����i�NqzG�s��ϊ��AΓ�����e���M�,I�I^�o�Q�r�%Y&������!A�E�	C^^�x��G%����� ��	�(��;B|w6#0�$�+���{���^Q�h���5F(��y�@뾖�y�*G!��#�9��)��f9G�'�#����#���e��?'��:'h�:���l�80/H}eF:@�,�J���s�Z��`�W�<��ueo�ŵm����'!��7儒�|+���8��.�~�ǯN��Ǟ���1�nG]y�Y?��	�t���@�q8A��rű���>���Z$�[���B�/��%���].ۼq�r!]S��H=xQh�K�nE[��ٌ�=�[ů�p�9���()���H6��Z�?����D�4`�Jr?𢯪�s��tD��Z�&���)%ɊQ't>4����brת!�4g.�o6��~ �MG+CV:N<� K󎕶<n��\�8f���<H1\)�ょg[N�0]�5&�%�h2%��p�I|^��)��U��[!|mG�������TQ��kI��B�a�w����?pea Z�2����Q�5x��W1 ��>�$C����BWHɯ���}���=�$j/-�:m�S@N��^��E������Y�m���V%�����+��#��/܀.�wx%�K$�k�qz�hyE��E'*6Я�52��]F5q7H?�<.�V���X+]�wz�k+t�F���E�j'�F�V��N�u��� G��ħ��	��e�ZB��~��k��,�d�x�Rz�%�l���7tcz�s���J�llģy��_��C}��Z~u���W�'h�̶_����A(�n����J��S��6��~X�Y�&�`R�rx�}���w>�����M�ɳ��K�*Co��'4�j��[���p8(z�M��Ci��+.SmWS=<ݵ�u�"8m��r;H�I]_��Yg:�VLY�|�������y��i�Z�Bכ�+�@��+B�罊���V�`R�=�����yC�,��w�����m����y3��VI�ܴ̚����e�y����?wy�,Wr*����~��뇞O=@^}�+�?��k�����}���|��'�u�3��8�C������@ةv%Ov;��'�ʝ�n�Wn� �v��sl�ƜϚxyBwT�]��2�+3���W�l�$��_v�p����UkSՄD�&\	1��e6��kw&[e���b63
�ȉ�]���dc�^2�
�?��}�����d"�+	G�$N������P�C�8V��)��7ג�X��X8р>��_���ϰf("b�-Hx�B�>��M�0�@���a d5�@!����5r��Ӽ�X㑶��3E2��O�^���9l�� ��'8b����tw'��)�odFp����$�>���M$�p�����ў7q�V��C�c�΁2�9`.4�q��0�߇50�؁����d��1�{l/���k"��&���+7�%!s1��Od�Qߖp��F��0����ݍ���i�T�s]�>�D��2�{ka�b�G���C���+M����K2��u�O�;G��EU{_�:2��C:����wMw�cN�j�3��O�[N;� 0��=���y�#1�{N�Y�4z���.�f�Kr�+�<e3M�z��N�ˑ,�u 	��S�<�Ś�(jp�c���&[�}>��89��Oԙ�������Uq(���l_?ͺ�9��@U<C2NC�>z�r��wÙ8�:��4�{�C�e
p/�,���`$='�;��W���R��4���%�`�5W������^�g�w�x���mPO$D9�>�!�i���8�7i^�-R�	Zj(ӗI���)O�1�8b�c���Ok������d4�~m�F7q7�	4�x�P�9�	~��l�~����3#��
�[�O�t"��{�{�%���Ǹ������~�@Tq]����۬��Y}�����m�  ��vP��z<5$IF���a~Π���±����Ҹ���w�r=�E�Zy;\䷾��b��$�"�����^R����"p����i>���IȲM�����|$.����tN�LI�ğ�gI��VջȄOP��꼭lqf_�]�	}N�pz��!aBr�"O*A_US^ܑ��ż#�7������
�n�8�f�,���Jǣ�0��^��ڕ%%(p�Ƒ.�b.��_r��j\���J�����!�[�
trP��p�4~$BY�,� A���3�$ۊj����9�>��7ps/�Q�%�nnCt�y��r��x���'�: �~J���.�_�7^��X��h���ЫP��E�Β�2�Nz��'�[��K^�mN�m�w�B�ׅ�`�f��Ȯ�L<�ԚG8��y��K����k	V�˩D0�Ů72=g[��=����$���;&��jZ�,��x�۹�` =�m���
>��ߩE��c!�ٻ�E�ߐ���������'-�~�#Z�c
��������&s9 �X�'�`��S'J��8���*�2^z_��u�<$!*�e�/���ҁyl�%����uЅ�o� ���U���`��%���O�j�� 8�GA5��r�Te����<J|?���i��}�p\�?�8<h�%-�Y����p���Uy8��pT���ǆ�V���B��*�y�b��\؋�4W�h%��0��{���w>�����O�K�\;{��o��[��^���L�QöWeڪF���e_沝�l�!Ϻo~谇���v[T���}-4>�^}9�L&�L��斸C:B��]��y���>?<�������W}�[�����6�)lR�f��"Q�m}�+`.�v0�L�������<�/���~���,gg�E������~��g>�~����y���������|���?q�X^����5�s^.0�3�i��^�ie���"�V���oOv?�3��v_̖0PM���ާen~��#(�et5��es�ue�ٗ=@3hwZ��M0��M�b�s�f��U�=a�AG�3OJb����5�3��:7ᾲ����޻+�����jF�[��c8���4��I�qFn8#[u7�5T�%��(�V�N������MHq���āB��c%����S����"xц�h���0H(˸��<;x��BW�Ĝ��ƛ�y��kWȘ�'e��Hy�5x�|)�����	�A�=����+�Վ~��&��a}�T�p��8�}Q���!CxX|cb��9����(�lu�p�@a�xK��ˉ$���B�����)�pUXя��6|mdD7�}L���+Ծir������~�o�����=6�J����N�#)���&X�s$��Na�"Į�@���R-P$"�D>&��0EM��eA�#_8�0�|�O��9��!��anl��S4�� �>*o�h]}�ƶ2j�.�*�x��+��-3.M\"8������9��n��v����}q$/�^z�b��o� �Y���#����a����w��s��� ��$9�y��kYr�<���]��#h���:W���}�]�O,"q �<b��y�%����c�S�O���-9���}1��LX�#n�<��<�y�H*uHAA��Y%zkq�Xl���S	j�� gI�z�v�]g���L�á��~� !���6��'Nt��N�J)iM�����I�9���	�m-�R���ȮP�a<";���l�Wo2es���BJlY���,����Kp��J�0I�Gr�6����6��E�)y����tV�3K�_�ƃ��;�E<9)9��]���g�}1|H�"��t
f��%�o�iO�N��q
��xB
���Z6V[R\��ʛ���\�|�o�'*�mG�S	<fӪ�p��#���b0�H�߿��J�W[/t0���j�D�uG�^i|	��СNԺ=��}\��i?k¶�����A7�w}�*�������J���5K���o�	4�ߐ<Ux@���bNI�մ���N�0q�����K|mI���n�N���p/t#���0�:�~S�ߢB��Q��Z� �d�ec1����5_Cq\*¸��>���M���\D� %��7$�\=��oS��� ��5������f���J`J��\�@N��O	঄�y�'=R�d�a9�[���u��l�`ss�EƠ���ğ��HާV2.8m0+�8I �[�S�{��p��Y�s"z��jG�&I+�"�V��|��L�}��^n2��8���a�ҏS&����3N�lt���-W���b �N��9�W������@��K�r�ֱ
�3��ڱ>�>j���Qy^+=#����t{����c�Q5�Yp��Y��aӣ�����`�e�q0'MZ�}6�;Y/'>i��*���j�eb��^�`���ׄ��$�-,o{s�W�א��a��萄�CǋӾ�}�#��Va_I�q��6I�U�J�>.�R�]l=x��Cjl%�f_����wH�l�Ϙ�L���W��j���^�_�|g�X~��/~���b����J�^�����|j���Xu�_\�B+,˪�1o��Ԋ �ԓ�%�tg���/�̠i�^(	�ô�Zu��Z�e��|�M��Ӈ�n��g_϶�[�FL���?Ha2s^�x��������ǯ��������7.��ؗ��)���s�\?�|�	 ���6O��赗?���7��7����˃�\.�ڦ٘�(<<��r��֬d�2�ye�����V�{�~�����Go��/~U�ʹl��4��o�+�OBP��-�UY����"�n.�����ѩG�]��E�����
�{]� ۻt�3�	����۫���*�M�<Y_ܟ��+�P>++�X)�����p"ZPd±�	�?%!��.}$����.�c�ǎ-�"TԕrS������lTvh�����?Ŕ�'7�Ի�oPBi��9X|�(ѿ9��%_ڇ�A�dq�O��L�r_pĪ�_F�^�mV2yާ��l�5�#���r�@|��}6�L��lv�i���h����\���SN�F�N-�f�Lap�{�˛��9��l��� A6����+�Ё����k�6��;B��<0��,�Q����f��ϸ�w-�'�c��(�J�y������$�j�W����6��/��X!v�� k�G7U:�y[�I�G���JȀtC>�b�6�p�в$�'�c�sD(�5b,3l��)���܍���n@�E{8JЧ'�QIN�%5���lX�ޯ��_O�(h4����r^s �a}�rco�;x!��ݡ���Y	A�Hh���P�Y��G����:�#�S������<��m�d$������<^@Ōt	�Nkqv����
���p���bwN�ћO(�4�����3GGq4 ����C�LM��B��PЏ�ٜF�����^�w��U��=r{Ob(�{AĠqT*`���{��\��:�� !�c�r,���V���������]�z�d��3�@�5,!k�OHo���,Gzd�	4-�	w��T��`��?�o�$�6����_qӼeN�z��"���`Ρf|��1�)�|%�!q�����+�ǵ��3&?0N:��_�X?�,T�n��������S��v0���N�������1v�C�#D�a�\���<0�Y^v�@W�#b��^꟨H ��۶HH�DG�E����lԐ��=�=����e�e��t]b�{��~�����Xk��ɤ�ƫ(��i^��K�4�@�0%p���fB A �>���-�w�)佟n�=�.d�_oO�!T���= ]��U�4=��}�}{����0M�G '�kO�g^a�t�j�o\�
������0
��Oq:dK!8����5�����:[�<�wI�.���� o���"A�F�.��~	���OK�1a��I���q����SqM�l��l��u	k��7dD�U�{�!�7Ȃ�=��6�I��
�0��ͤ����_B��ݍ�`_0p,�W80V4D�bh�'�AJ����@K�V�j�D�s�J.�W$��n��IgzD�jt����d�`y}�UI�&tU7�V��&��|��!��@��e�Q�ur}ԭk��5��tI�j�=X륱��?��3|������h�z�9�:���r��r5��v`%;��t�P�vX�A��T���7��՜6㕀5���w�a�o!�~xe�v���;6h�k`9![#��Zb�]�0߬>)Љ���7d�e�1U�;=Ia�4���>%��տ���/V��*v��o������y���QΊ�-S���X횭w��U�J��Z�������� ?�~�*g&�y���>�>������MF[%��m�IL����O~,�,���d�Fӓ_���υO��J֥W����+�3����������_?�/��S�����~��?���+ ��r}�6���/��;7�����*V��*�����@�O{9�C�`��߃h���Io'���$o�/�_��m���E�0���E]UkYH�[$��
�jx+��ɘ���U"�F5J񃉏.3��[1V�f�x��v�~���c�����\�<TMB�B�NVz��8�|d��B�fjl(��x��׸}�%r��ɪ����E0�R�`�y��FK�������D���uxV-��1��2f���up@� =+���p�l�o�}�s�>��I���)Æ�͌^��x�a�dGS���=h�`����?}�}�QF�ȉ#)�(I�Y�Wϊv�ʫ��Sdu�������k�mx�XGӄ�F�4[2d�y0�L����XOq�M'·&�1��	��z�Lk�6E ��H�w:	R�j��m	�v��dz�}�����ufk��lЅJGf��1M`�X�d�KsF ]����_�ryԧ�=9Ȑlw�C�� ^��������(��$�/�Z���)�փ�d�.�Z,`՛�x^�+ίH���>/≺>s\.3���N�NoG�nP�eW˲F2�/"e��F��cC�H/W�&�=��Ew%�x'��%�s�H��S�bG����-��Á7�P��6gP#��.B���Hz�S�� ǯ��pl��^�Sg�o{�U6�8�ͱ�o����t�
���� b/9�
}
���%��
ȑͯ������J4�y�(��'&dS��$�Ɗ�W�}IL;\��!�H�v>c	���KH`�G<�'D��I#Z���d��$N#_N��:,�G���)�\��Z.f�����_��B�XbK��P���|(gԙL8�ڰ]$+y�2��Ao�6�αD����Ӊ��%�������ര�ln�;�a��vݵ�ݫ�˓�pʖK�Z��1�t>��Pr�&��aR��1�7P1d[@W'F��q���Sgh��2(�2�a �D����-��E:� ��+�Dƿ��Z<aQ��F�WA&��b0;u�h�$��M�^�02�0t�2�,CO��_f��@g�� x�|��6:��|k9�@�iJO9��ۓt� e1��S=փG\B��^�d������d��љ�%6��W�T���}~ĉ�?��Q��n�"���.����#��&ۃ�p�������4��>[�*_'�s`����T8&�p�����'��i!z�s�_]�)����p�*�!1!%d�x���J~�����7�A_�9�r����n�!��I�T-�/�g1Y�y\Ψ�Fs�>�S��}�x��ܳ����CIa��� wb��R�.+����b�rޠ�HF�1��&�I��wp�w�P����T�=�I�j�MIp�N�r'|��<������0�����y�˫���|�����n����*	e������<;3<i�CSo��)'KT�m�J�Z�sJW� �=���F�,��u�%I�<���m�O�h�� t>���_QR��y�7�ō%�G��О�5Hm�Tdީ:!�A���c�/�gix���0���S�W�Ԡ�X��{�D�Of�Ak'�Te��~��<X���ߓ�0˟�]_�q��e"t�1Z����w
F��,Jw�>���>��v������ծ�(�S�%�H$��{���9
n<Z�����u^O���u�C���ޒ��<�#�8KZ�U3��b0�����u�����;�_z���_{o)�U_E��S(q�\?����ϟI����l�w��|���vxnj�L3�\q;R�\�߫��&=VԦ�ڂ��/w�+���������|��BJ/�����&�����¼���E
ש�ѯ��3�F���sˡs��皙��o�q�W�ل�v��~����'��?��ܝru�[�v!N��e~O��QF�sT��Ka�ll�=B`�G�0��=V&�@;R(�B:�d��!�������
�*�ڼo����;�`�Y�X��} S9�m�(��4 �PLPdl�y`'�]�%x`Q�O��F����e$ՒX���0,}��X��:�$<�c�����F���ߟi��'j��Fֹ�a�e�o�ic����z8y�t��b��h¼�"M�N� k,%��H(���].���ɨ@?|�<���p:����u��p�o�����){�b�
k�������N�Zi�a�p�KT�p��|�����U�66`�����W�˵m�A5s0U��H�^{ּ#��'��{��?�o��p
��1��~Q
??���gLb�>h> ���Qf�p�@���\�A���d.'�!)�S�7�|:�c\�ACv��p����6�u $=�K��Hd��}T��wop�96���H�GݝRPnq	5<�$��g[y�b�i.���|-k�N�TX����!�I{BR�|�Ю�?�T���C�κ�%��z¡	�)�eH��pz�˾w��"�o
�b�����i�뾇�q�^��j�|�7��Di���O캎���\�>�˽���~1�$<���?�?
��=���aR����"%~�,p<���F�b�?��c��!p=�Y��W'�8�	�����(/I#9}q�IvTw�P-�Qָ�ܖ9:Bp+d3�m~ط�e�D��7����2��9��-ư\b(�D0�h�n�[?ˉ��p����&��(���^�,�B&�8�	�1��W�t�j�K�Ѱѭ&���AE��;�2����G<��:=�^\a�,C�.{-�m��x��1D"����W�>Y��`��W��bG�8�� G�����^�8����d��O��.KK��.�[J��u%�-!N�[q��;ۚ8��״�S��"M��.^�6P�Vj���Hv�ˮ�/~���J;�Y���U�ڨˠE�lWpt�.&K\'eI�ЙH�~�Z	� ��y�����h�?:�N�'��k@sM%6�� �[B���S��$�g�B��P�ʂ��6cvӂZ�t�aN�,�WJ�� 9�k���\��Vi�����e��\]�h�Y��'�1�H��'�dh�/��E:�]X'�}�\�B��u���vM�eU�W�go�u�f�J�K���	�B=�,���ڷw����٫]1ĳ�ߥ =��/�P1H>�6y�k�>}g=�� 8����x��:�`��Kld��P=�O�G� o�0�཮�+@1��8��.�4�|`\��]��xˬ8:���HS���Z؎�J��ag��d�w���	�4�
PNrZJ�������²����"�b>��n���l�/�Ͻ:��bo�|��	�m,><�q��	�H�p���&�o=�T}I�_�?���������G���O��X�3��[�g=	SO�k�?���(z��j&쭞��%b7���oFFwR]o���T�2 \�س�[�[2A�ą�����]���ߕ[��������(/�Z�}�~0w{_H
?ۦumw�k��]�+�.kkW�������~~��& 4�t�b}�>}��}뛟�����k�L�ҬɘlBJJ��k�!r�i�7�	�����w�^����P~��?#��}G�*�7��_j��V����l��e��}�Y�	5������,�ʇr�,!�m��g�V�7�i����_>����]�[ro��98�yM������e����Ĵtx9'�S��u
�2Ɋ=;�-�/p���
'�#���
Uj*�U,���IYw�Q��l,��6����i�ƃD�EvN�pq��������b5�<�,����zЭ�U떋J���%2�Pf�66��c��R"{�X����� 1�#ü1��0) ŷ;M�|���'j�*x)^n,t���Q{��I�y���w�g7�\n���<���輋�n�nwv`VzJr��%�&���f
9�6��9ɬ?ޣ��!|��1�Z9���8\��	Y�ۅ��`N��1��9�����'W>M�hVx->Y/�x��hUe�-��϶o��݁i;u���x�9ۊU}�s{���]n�]��n	� EK8
��gq��oA�bN@��wQZc[Q��>����%_����r"L�>�3���ZyD�~}��+'0t\�s�\n!��?!?i����h�� |#̡Z�8),Ȇ#�!xh,�w�@^��Gv`mA�Ҋ]/SH�c�p�t����OфBW�8��=VW�(W�;�p�=ӹM�3�,��a���X��G��o
�ib�&��G���8p�������pW��dU��.K�yO���p��kz?���ై9���Y�B�&8XE���.�,Y�UD+%��`�C(�"��,���%���X��ARa��.�pנ��ICO1O�=���58�c�����+y�x��"�+=�gk�[L�h���8�B��pP"Nc��*=�W$���䌥�%їˤ�&�:��ːM�9�����=��v.���@⌚��Nq�&x�/Q���{;�$�8�%��Cf���nQv�`z<��I)L���7q����.N��C~# ��<e��m ĵBd�-!�|�d#�n��˹f�`����M���+&�P\�4:�!��a&�{es�Ҟ&YPp�OMe���b9,Ƈ��'qG=l��X5l	1��u4��z`��xl��* ���d[A���������zT��3�����P�eG!�@�ϟtk��`�)��h(��Ag!�c���$��2�(�M�J�Gp�w�jI�G
8�>v��W����W� ]���OҎc����T�1q�b��奥գ1U�P���u�QЕ��!�]lKTHJJ��m�x	Y�06�a�'�6��v�'�2~S"��%�ŕ��/��(�dx��R���|�+��l�P�Kl6��c��w�aGt@�oM>�P�-�p5��8#V����?����s�/dJz�؞�m�=W%�j{�'2�r8
 >�d7y&��cM7o�]�>���ػ������Vyg�|0O���m�7�w�O(Frz�MW��ʪf+�9{2��f����	T2<w|q\
��s��$�	�'�	^j�B:7�.�CK��{�>�a�H����]�xm��/]�P�ߕ�XWa�8��w�!���vZ\��!ǈ��#�,>�BSi��d:���%�WP�~�p�.�ఠ��|3���,�E�c%
��/��\�#BDҖ��H����q����vMm��r679����l�?������~N�_�qMX�]�Wg���Ħ�����}Sb|���:>����҈~�?���ё�y�
.��~%����Z�q�T=χ�o���|�����$��|�S$5�~�����,�\l����+���}t8�����z��rgk��ߟ_\\�������~����YT ����ֿ�ڿ��?�����|���}����ۿA�b-�Wf�����޻�ږ$YB�Ͻ��gFFGfde���*
�[�j��nh��S�����3`� 	�3��g���[H%h�*uvYdgfdfd|_��=g�s�͖�2?'�Q����x��s���nnn�����D�q�ʱϝ���/�_|t[�o��O��������??i�pW�:�63!�Nm�0v�c��vA;u@g���˵[�©ms�Sg,�`��`d�o`�ܟ}s0��8�������g��O>�'�]����C�l�:�h�v�&��
�h]b��#.��A��A]0
�ǿ��������� h�@@��>�:L�	�#��8����3��'���4�xw�y.6��lw��ctЅ��V�+4��n$=�RG2K��MVچ�?w�������f���1 �Dz,��e$� � ��ỷ<5yNa %��v�s;Ȱs�Mt�3�f�d��	@�gޯ��bV�XC��GcEp�/}_��<&zf�+�uj+v��`�Ϗ��$Q��R��>C��>�B��Ҋ�#�×40���=3ȅ`��$~Nl�Q�@�Ԉ-� h�*p��Om��I�N�,�Lf������'�,��:'�S�vF/@��#��_)8���
ͩAF�n�*%	�9��e<�F8\�r�*�c� �W��x��1x�3�L�!s��!�H���Z�6�-�]<�T�Q/G`X�ڜ�|��6���R�|d��'��w?A�ο)�>�Ya����!�Ս9i^�V��w<�m��iN�e����+@zL�1�#ϑNffg�"��w��[��j��9��5	KiFz�D������h!�����=v]�{��_�6�}�,xd���h������#�q�'�Zף��;2 G�ԍ�汮�X�b��X��ж	�=W���z�[neT<��s/��
����U� ;�l���	k�ie��Z`���*5��2�n���.�J���A����ރ5�D�%�$�# ������I�i�Y�W���@�h�����u	�aη:�vtX��^M�;)th�H������7���G.UM���~�#c)O���\G^���:f�賠%�����zWb�s�IO�#�ʸ33B��Zd��Ŗ��5�����fC $;��Vt�av��?�S���+��,���f|���J]p�a�QOJ`�&q�Q�SS�o-��R[�Z�>���к��ۦw#�
��*HΫp�n���m�W�r�|a�Ӣ
�@
Ƹ��z���t��\���
�B�ⵋ%��AI��_�n+BP#	��k�W�ln$a��l�2�u���Z����}��s,�.C+��_b\Ͳĺ��I����d?���7�\rT'�{].Ƃ?],Fx��Cz<�Y�Mݹ�l�D�B�3�d�jt{bEW[<����j��wt���#�8I�H$}Y�.���Nu�(~�&@�����}P�VA:�nr?�i���hy���^2i`�ձ�g1�&{Xy��S�铍_2�e��޽�V$�X�m�콋�H�@��ß�^l�:�ߦW�G�i79���]��/��"F%H�X�a�b��k`��%>
�un�vB���7[4��t���i�2��@�u�/���ֽ�}�k���=��+�j�<X��a�"P],	Nqa�E��7(Eߚ��v�[�O���1��-�X���2��BJ�;��-_�1�X���0V�ynKk<���5��O�d���������cz�O���?C�O���#�|>C<�9���
G��a�!�����]��h��������^Tp�w�C��+l�r�m�q��H�ڇ�W�����F��Ogb���M(,R�+6+&\i�.��"~�J>�M��f�$$ڔ��|�O�A^�͏�Ԓ�rs���"�{�D�}��z�yKn�q�q̑U<�� E]�6�RQ�yȂ}b���(����(ُ��������UQ&A6K8賺b+'i�]������X���|��0�=�z�U�8��Y�g���6r��ǈ/X��8�z���g����?{�?�w������o?~����o�=ȹ:u��������� ��:<�������7��/ޖ�|.��j�e��#[uw�d`��}`�;z��6w�}�^��,\�Χ?��/��?���,p_�$��<�>�h�"��9��� ��Y�% \ų���\p����̣	���j��Ͻ�3\��ԓlg��ٙ?����O>��7"��Y��?k��4�F\�NWs�9���T7C�z�'}(�n�M�oL�nĕ��39��YO�	��R�p�Vxzc=L��L&.�;"��\\\���;�Dp�;�"P�'�N3�T+M%�Џ �%$d���v��k�r	�h'#e�Znt?�j�{xn�Qx����'ZG��(7ж��^ǀ{�^�;��/�.>��6!�;���/:/�����o�s^#0�Fi�4�#��I�H޻�S���9�Ð+�����q�A�1���搭[�ׂ'0z��QK5Њ�v��]��z��"lw���x/uP0e�;�Z��żڍ���W��W�PV�I"��AEv`7��{L(�������I�����l�?��֩���>����{���,������<�/���x�����>;��q��k��Cs��]�0�1n�LP���DA��ِI*k��C����V�UiГNNw8��$n�\�k� -��b�����`��:}�������i{=��J�����q�����+V�4�Y�m|�.ҝ����J±��Eл�B����d�=�rM���ۜa]��eC9m\�L���V���mZO�W�|�c���^�ꀿ�Zw�z�X�F��ɹB�en��6��s)�/t��{�ċ~�P��Kz,�)�WjW�I�a��(ڝ�¼k�y��d���W~�6؉ï�ғG�b.A{d��p�D4��ԗ�W"��Sp)a���:#����$�KT��$ӈǕ��"�H&�}���
�F�X"9ωwty^��n�c���?�Naǈ��50DeY.�i~����Vi�6�������$�]^�ׂ��~��q'�컞sޤwZ�����@�Q���%M�ڡ��rD_��!��̩:b�f҅�ͱ�Uʲ�˺�g���r|-��[E@�_���i�[�����Ǭ(f�`/y�1N�S.�L�}ͮ����6�V���g��㒖�U��v�sw�u1�� l��m`�*=imQ�}Щ�цƭ��1LK��EfM�<yi�Z�s�� ��n"��	1=` �~l���O
ތ�'-v|T�	��`����;�|u��cU?��u
�,�y��� ��L�1��'�5��;"�]�M;��X�ϊ��p���L������&��K����K��H��-�W>t?�y��r�1u)(#��狝���3��f��!�}t����m���h AJ�$�V��CbX^%��xu̓�b�2ߴTQm[���?�ү@���Z0�����w�J�ڼ6w�>��+$_m).Cj��5�{���Y��l��EWZe���!éﬣ��C��s���6A$���i
؆dń��W�}$�:*�$�î ��
��	G�Xg9�0q;�]���!�fLk�8�2��cr��k~G��6�F.�	��x��U�ĕN�����;��k����_�cCg����G/�ʋ"���o<zSN�$�F���b?��f2a����%�	J��bS��ݼ������_O%��w��Ա^�"w���`�q{5��?k/�����6�s��'��o�3>nl�i[dsJh)��mTG9n��>��}y������/���7���}��~q����~*9�s�_�����7� ��YV����Y{����;��!�7���rF�����n6f�s��,�f�h(�Q"�ii��A�?z��|�'����^�����-�%��9R�Fy��03];�z��
�
�q.�;L=%*�[�r��>�� �#3|d���S�##��ϏO�����姯����*�F6��Ω���'�Ur<����f%�kY�����)FL�B���
� ��������s��-ޫ����i!z& �	dd��E��)a;���c�(Ol��(��D����HH�}�Ē��x��RF���ei�礄�ھt:��[vh3J�S�L��c�_h^�ᐑ��j<�'�á
&���/�E3ͣ`��a��]P�t)��7Yp���a���~��'4n�N����A�Zܨ��$�ﻓ�w��tg'���m���&������:�A)}mC龡���:Y ����J�nl����8G�T�����{�᜝[A5s�����7t��Zا������ő��gT[轑�q�����Gh�(:����;2c���{���m�e38��Ҝ��+P�� �7��ѺY�Y�]r�
��[�h�i~����ۉ����ɴr�
��b2��2-�n�F(V��8�1i��Z�za�P��
����8=�mu��Z��RJ
�EP�dْ����Q��Ti�նk���y���_�+���D�!İ��w�r`��<�9��/��
�o��>��C˘��S���5����3��%7��*�U��'���'�!�[���%;��y~]�\�.��9�G���⑂s�}�2�_�5X0}�uI��DNI���]1�Ǜ��R�c0��!~.�V�_�O��M\Љ{�CκeL�6:d�1�����VC@��a.�V�	��7�'p �J�w�_S6�=�/x'͐}�:7wU���=�@e^:՗[��ೡN����WN]k.�I����c��1F���^��ه�]�W���{G�}$c]���3� ;��ƭ���n�����-��!X�`�q?/>���J[��?F�`�WJ��sP�&�9�۲N�E���U�ּ�N�du��Fs�ڔ8TF,|���+� ����q���Kۍ�V��V�1����'�Mm�:�L���6�6�w�B���+�"�[���:J	�]u(օ���)��4J>« с�DE*�ߓ�D�p-�-�n�I�~�%��6w���(I��%�{m��Nwa�O�������#q[})�2��q�a�\�,�Z��I�v���g�l��T�]�0~�G?�����	;;�6� ;V�>��QLr�`n{]Et
�c �#�a��dRʎ�k�G�d�l	�(�N�JW�M�˥�T���4K��R�$���R���;\�����ԏ�"0Ɨ�QP��im���]Ij�k|.��cm�Z'w�M��S�����|��ٶ��[��i����ꆕ����:���A�9�K������7j�G��kp�>R:ǡ/I7��@~�n�茕 n�!�؂d&q�v��SIg��b,D?_��u�z����d�I�����Ϻ��(`��Q.;
|`4>k[�v��XV�1]:Eg�Pe0S��8��MQI��A��u�ŧ��|�]��7�%o�iu��p8��˃�v�M�Z"d��:�9�J���_���N��V����Пz�b'9�rq?I{y�����/>��듟���ߟD�V�f����ͅ>�vF�	��d�I��n��G�w:�r,/n��O�y�������'�~���8����_���u}���P?��|��gg�ogK��v,�0������T֒2���&�O:���f;�g�W�g��rB����[��&O~�c����@~�������e�Gp}���d;w�v�p��m�)��kjX�����s�Q�(h�a}�hF��6�;Gٗ'���_~*?|��|~V&�æ
���i���v��o �]dir�;$�E���@r&�r��4�@����!�����?}�|�$K[\�h�'��sF�(�@�\�%�g|Յ2ŧ��fl\��0�� 5�]V-^��hLkP���ߵSq�%,�_$�F���	��VK��&#�_|���qtb��K�$�˻J�?w
��������egQ7��$��ܽ���܈F��x~Ԕ�p&�W���!���q�A=�Σ^O'>�-6���#O���)\&�t|M.���+����,���ȱ�F�䳢��"X�]����WG ^���0���qy������v|����ϣ_p��#������ϖ��YN�����)(>!'�v��P�L`�Jȧ�[�=V'���g�6�ݰ0@� ���>w�!]��"�7�A�Py��LȮ��c^��:�t�s�}�E����JꂱW��7ˈ�>�y����I~�5l���r�
�楎q$`~�{3� ��D!��7�Qb�~�2�
���]�1X�u�r�:Z�P���.K�x~��	��|�t��c�X/�N���K<�Ax0J��^|�a�G_s���S����`\E>�6>�0O�.=9�9��I6���,#�\0���?9`Nk�����+�_�w�%x-+�p�A�����������V� ���06Kj���1��nf�K	iZ5���-X�K>a���\�eق+ˤ�?�-\��y���R�L�0��Y��L���a).�}-�m�=<��0����7��A�k <c����o컙� ��.WE�H�x�Lڤ#+���4��vQ(�b����y�z���}����_��6Ӌ1&�[l���Y;�K���nMfYH_J:���Z��4[�e���.�
a�����!G&0���0;�{�A/��T����1֢NY7#Nޕ��9�#�{�e>��l��|6�<Qv2>b��U/��$��1o:Hwu�j��a��ٞ��DI����90�M�L:@D8�2�ߛ�y_ƕxDb�.���Mئ��T�	b^�����2�����G�}��=B��CO3=���U����/�k;c��p�R�V�����Ja�=�A>�]��<�����챵�C �:q���e�u���q�w�&�Y��U��l�3Dj:r���}�{7���hrm-0mϯ�E���� �w�R�TO5SĎx	����o3i|��]�4~�R�MQ#���=��|�M:0�Λ�K�W[�]�Q7�����'э�m� �q�H	an��Y�M���N��~�&�va�8�|BX���'�r�������+�k���/8��}��lS�G�����ڷ}�#�i��;?09�t�V"1���:�B`��+=|�ƛ>��a�l|Rx����T��_��*�Ue�Q?c7�C�;�6�5�s8q@qS�N�ꉉ��Eqd���:��z���.�D�c`�ܻ�����%p_?���	YH���<c���͙1:]��"t�%^m�8G"�N�ȘRwQ[z�ι���m��/������~W޿y$��>�?n���.����'N�����@��Q��(vR=�~+�&Ƶ�c�c}�P��$϶.���*����W#���L���1U���X��&X���8��m.d�a�����X������o><��@�|���������� �{������������_}��e�{q:����T����@D�pm���̷!@MɌ# NS ��>K���$w�|�ه���~)�{�&�>��g�|k��SZz��2�=�RAQ�3��s��`oi
|��ษ��'�`4�/ύ���K�??��|��δ(2��j�2�X��˭�c���:.�T(�l�kz�>�Ds�dt���>R<�:)� �30l%���M��.2@��I���E����ڟ"�svK%��쀳;BP	���p��hM�СG���a�e��Y�xJ�3]q��t���l���ƑW�х3XG;��o��ݬL���v3Vx^\�bA��Gŉ�(zJ��1��Nz!�A������{<o5E�
}�~�����2$�D�>^s�z�=��4}'�Oܠ���%��Qz y�O�m+$ñ��*(J%���ԂXݼZ��QJ��bǕ�N_�;;�����E`���跍�u8I��B8��׶�1Nv��>)O�a/��C�8o*��<�$Z�n�=;���ɘ������3��iV�PP�P���3L��@�KJ�P�#f��Ӭ$~�Ȑ��E�MF��Qc>աg<��m1�e���e$S*��hi�
�_r�3�/�,F<8�">��-*ݫ\Q����rU(�sf�}B�V�n$'���ud��0^�]���0�y�C��v���kf�O,�m�i�ר�㲯���}��p����m�i����7u8�����;����`T�-�=�P�296�J^����Mޭ������XkUzjzI>�:&��W�e�?]r�.��y��<�k�_~��ݖ ��as���Ҩ}Z�h;8=vri�Ɓr6ѹ�DgO ��������мK�9G߁1()�F��&+	��D>��)x:m\���9K�M{7�n�\�ݘ����
���7b���t�/p�:6n�ay\D���*�� ?-i�q<q�1��>>��w�^]���|Ϟ��i��B'��w���T�b7h�Ω�1Y4��H�%�W��[�"66�Ҿ�^�g�2�3�dd��G�K����R����\C���a�������\C"F�y	Y�I�X���L<\�lY�$\Cr6J��-M���98�ݹ�є�"��@,9�<��_��8 od:"W���W:��^n⢘|�s^��a	8o��AIz=]�g1g������tV��e�?�Q�.Y����+� ��)��}��D>������*=��B/�]߱��I���c�8W=������K���[z���J!3�Y��Qk��m��/��0t6c��a�W�@�Ꜧ
��d��#&�Ơc��(�N����Xr!����$*i�����&�W����%���P�R)Dx���k�T]T��<��c��spl�5Y*���X׾H�^�<���N�l+M�L鰲��l��B�Q�1��]���I|���ZҤ�BS�'��I��L��[��m��G�������_ٌR$�0g,������:�n������>޻�/��.����}��OՎ)�4 jk�u?n�&�K[����}�c֨O�fU��A�"����.�}��,�뛵3x���Z�m�J�Fi�#�6YX�b��IY>$�����Ik_�,0g�d���~#�{y�=?=�x�������d2�mj܉ƛ���}߼�M��i���3���[ޔ������(7�7ӓe�5e
U����Nr ke�N�k@?w-1�A��n���v����d{~���f�?��C���?���&/�z�vϹ��ٗ��t3lGsy�q2-�-J#�{L7|����c�� �pܿ9l��v|���o�����Y�_�{G���������� �D;��~��_��?������G?{�⃻[�Ǧ����$���s��B� �xB;3yi�������f��.���_�ozyS�?��|��5�K���|��5�ُ�g�b����|����^���Pb��|�C�����PC�?�M>|�T~��G��Yr?�o��4F8����t�C5�S��j�-�E�]�Y0�|<�u�}�
tA�Ԇ������{P�3~/U@�e8�t�g�]��u��� 7��s�`�>�>��z�/2���ٶ�t�f@�~d� �9��ݚu�?0�w�@L���L����s��5�#��.�K�X&��ڝW��DK�D���s[��g|�s��4�w��\��hِa�~�h�9���;զ�Ks��%�Y��0rVF.Ż��-���oC߃]��x~���vqc�û!p[�]n���d���cL��Rl�+�5@[հ�}|, h3[z��k:��%�}T���&�ϕ�J��3������5G_���xg\c�������T��#�.���"�X�0&�����0�Y��J;�e�Z��;���?���4���^#�Op,�s:;���n�}��+�t_;ڵ��4=]M�&�ż�9�I]�t�����MN-��t�z1�G�c���2�W�>5��b
v�/�󼇮�Hu\ky,�˽$]��qv�FZ
�p�p���>v:H8�msIi8�h�z�{���h���S��?����1�]�]��<��\O^Λ=<)a`#+94�/8P�* ���㽝�%��X����9��_��,}��L���>o
���ɲc��s��eb֠���|�w��X*� �Ӷ6}�8�y��f�EHN=�:Ŏ�Á����>sބ(�r�.��d�����m���3z�`�6?s��_��9��ڎ'�	�VCܶ���u�f���CGW2�ٷڸ���A�,�yKpf6���l���e�C���5`�t s���|u�~����>������]�1�#jjI�Y�I����F.���� -�0�փ1��+�o�����-�����=���T����[�8�{�f�_��P.�*� ��RBbW��$��P�T�@
��k}OG��^��ݲ�wEVM=vЂ����%�~�uƴ�%�m#���Y�&��K��3�=�2s7y��	�i�t�U:d*����Ծ����	I��=-$�!C��{��Bx7�AqY�����Y�%�>��,xh=�'������Z�sд��!|\4F|w˅|��#���Э�XRx��w'�?�>y}���:�^/fI�||��8�w���q�D�7Sp�����bO��<�g�Wp[�w����%1��3��d3Ξ�{%*>�X#��
q�����;�J����kϏ<Xt��4͢�d�@.����~��)��=��
�h,��-�m%h{1t�ք�������ۭ��Vld^nн�S?'��6���=��R�ՎCJ�%>�n*F��-�=�}��Ί�x�F��ג����j�t�x��$h��s�uՄ�EmL��o�@�&�󥧘]Ӂo��B�c�v�[�%
NLl��t4�=��������`]�L`s֚� ���Q���p}o�����ɏ&��T�������1�1�瞤H2~R�`���4'V!��"�37[g���1��+���'�����_�_7�s|�$=1凭i)2�'�a����,����|�T��7ޑ?���Ƀ����CCB�I��S��v�V�d9$�N_��e�c�D�6�Fѻ]������?����_������Am4�S���u����66�ʬD��8�l���х�i7���sZC{�o�~{��_{���;���o����۶}&��])e��������, �rx�ٿ��҇�w���~����?<��~�m⨼Z=�~���z	����QQ>ߦe{k��r=����Q&�n�o6���|���[�&���;�ߑom����Og�0�'9��-β�'�a�"�MAN �m�<�g�������/��g��Y����6��r����(�%V�f��UY��]e�Rpk����D�4E�IY+}%��*5�B�.���a�PPOA.w|S�@�>���E�d���'�����2���f����;��'����x)ŝ&s>�%4t���鋀N��Yѧ`�	1��<h�I߆���7n=�&�]�΂�L \����Q��i���P���fI��&����A#�N�u������W��M��j(b�km��S�� ��(.��g�I���� ��3�q�e�Ǿ�����r]����Ov0��E��B����ɩDk��r��l�%8�����2@��G3��wiJ.;஝�N���%f�<��wd���4cىF�����x����t�-D���dO���Ȗ��
��+_ٹGt��v~`1��p���;�V�NC�H!�|��#�}yctl���^�82�ϫ��h�.@!�Cc�8Éj�_�i�%��p]�9�ʜ���ZZ�|6"͠͹�!�r���9Ь����t`��}����e,��W��:.��zff� ���Z�:O^�{]�����y��ݨ����Y�^s�r; ��W�q��}�,�#�n��à�����$���im�c�L�3rc����X�q��@�c;i�*�q�O>6�b�@4_�(�u� �B�޶+x���M�v;~�� g%���P"�����s�rp]Kz�P��
3XܚWЄ��'���&���P�|�1�ck�C��谷�a�?�E���� �=
<_0V��K����2W+8C���ٚ ��%�=�Kj����mr�wu��SND�.)xA�p@+}�8�x��l���&��j�N�(��=�u���e*��d�װ`H�X�?Z�c�a0��Jk���r9�t���+�-��l� ��Ʌڍy��A	T����F��t:�v*���&i-�|���+0/��������ڬ�@{�o���G����|��^��y�J��oƊ�d5�rp�a/;oA��\����,�;K��?F�s u�h���կs$�Y+"�a��	�bi�8���Y*�>'�*Qp�љ�_�}�s�E����:/=�s�yX���Y�Y�bb����>�pn�Ҳ̀ ��:��N^�Y�q������j��>��N<+1β�7fm䣣BF��@�z�RA7�����x>@�$���<�hNOȷ<~��I�tl4Q[o���v�Ӎ��^���?R���������Q5��(
�P��e��H��m!`*�z��od"�b���YL�{�V'���X_=�IQ~O���,��Վ�T��G��h���m�;
m�Af��a
����H�j��b�Ðc�B::Fb��z)�?PA��(O�ҙ��-�8��r���z����k�pmnv�c.������>^g�U�s2VN.�
`:����E�N��8:@�I�xwV��,��{]�t����6�AWvZ�,��&*�D��6` p�K {�[�W�l)��4��c��j�9���_�{����C�uջX6��<��%�Wꌘk���ƿ/����l�<}�����cy��#�����wn_��{�[����a��*籩ӎ� ��67����$�ɹg[~%��t�_�x,��/����<=�s�L~�t׿o��b
t��#Œ=�PK�r��K�0#�$��nd��t������ۯ���y���z���C�����������F �«s��{��ko����[��������Nw�t�r��������j�>F� *�D�L��^*ا��x�`;lr׏��,�����O���V���[�����͛��Ǉ��]�-[Vk|�~4�jL��L[���W��o}r<�Ǐ��'����v����ߍc
�:��nkR���v��2B��<�b@g��ʟ2�/�������²0�$��s�虲�G�9Rz�`�)���;��x@��!``��AߍƑ����0�����b�A?9+}1j�N�8�h�+,F*��X/	@P�;�c`5�A�qͣ.��v�C��-fm-�;��(x��IT g��]�?���oZs����pT��e����6�b� "�N�=h%��9�5�g��]ƅ~ߝ>�⤺��9�o٢�qO�*�K���aX�6 y��/?�yX�B8Hg�5v��n%��� ��;�KoW��S����\s.+ݚ;_xwa:�m[������5���;b���8w\�A�rY�%�IU4�������f㌏a�<��jT������wG��cYiy����15�v���Up��;t��Ҏ��?G�#���,S��G�܁���uf�����4.��;�DB���Y�g���,+�Jǃ`ײ�&o�ʼ��>��;H�r�'�J4�U�oQ	�'!����J<S�y�u7�l����Χy^���3~��S�F��3�f��T�::o��Ԯ��\砧�hɊD��&/:x��J�H$JZ�5J�b�&t�K�@aM�,�@#��c�n�H6��(�R��fRX�AM�	�R��;�b�d���x!d�*�\��8�e�ǺB�V诼.l�����F�G��T�]��j�2�(�?�������p�U�%&��?��K:^�~�{:��(f����q4F��1s������k�sr�B5`\$nM�nEe����zX�?b���E�+�LL݃Gi��F��N/�� ��)�R��%�A�����o��J��5P���e��#��l�"��&\7{&��Xp�Kal��y ���Q����ةB��z9��H��☟"n�bκW��g�1.��la^"� װ��B�)p �U"����=��&ґ'y�dRA�\��L�)�>gL���'녞�1|�*�<��#�	����:Db��ny�.���0��c��2�*S7`Z�l	�@��H������+G�%�\G�:^�u� ��\ǳӆ��־w�.�%�k0o��>PNN�$e��J��O��= $e���z��0��S�$�z¡؈�(�`����#;�������`���%�l��Z�Kj�.�D�V��=��$�~��`�d_J�8;��^��,k�LҚ6�(K����VY��������?������\�%>����<0˴���c�.ֺ�1���,bYj�o�ֆ`�񳣊a1_��	|�Cf�%y�X.-�x��>Ђ���v�)�7*��kh�yޱ���6��ni�\�yYi�~�/F�����g���ta���ɼ����hO2&�Z������w�:m����^���>w-�b:R�=I{8]bmY"ӂ#!&tK3=�հ�A��6h�m��� b��f�?a�����;?�ɶ�iR!�;�!��E��g�f���P�?��u��,X��YO;���&��v�� ���\�=޻	0�'G)�r��~�Ϟ��ϟ?�7��|��#�֣G���Cy��h���I�8���UL�M�Ϫ��󟣒���I�x�\>{�D>�{%O�$/��]5����f�\kr����*�2�n��o`
_���a	�ɢ����s�_m�a}��_�g��_l[�y}P�1������������+ ���������~�����/�?���S�����co ����WWF=�����W=L�禥�4 ������r:��s��Q~��y������|�P���7������|�ͦ;�q�����������x!O���4Kל�&��C�(����v��n�����@U1�?q%g)	�ta��@A4����e���&���P��H���� ��f?��?`&�朠sz����q�:2���	�G� �q��7":	��bǍ{i�>���))Q�V��E�ܝ�۾�*�Zt�{��tn/0��$�  9�Q��ԩ,0@	�x�[����%�%x�+�¾w�~@�m��n}h�f�]����L�P���h]��_{�p�C�?�C�dDѶ����m:?v٩�[�� ��v%�?8 �B1pxu�!�pRt�]�>>�����3�g��fC���Y�-�w8[���vB?0���=V|��B8���pc� ����ae}i>�59��ݻ"�.��������{Z.r�XJ�4A�RT� ��,2[\�Q��߸����Qj:&�X&-�p*_��A�˔�ځ�Ye��A$�� O��\h��AZ��t�~���Qb%~�ޡٓ���8}4��*<8ݻ��F<�w��.d�cep�a�Z+����~��ww���t�v�e�-�5��y0˂����%7�x�P�)ˊ�i�k�қ&'Qlh���hI$b��^�q����ec̿9Ez�����+���K$ʉ��x�U��LH�o���N�B�Z�r~7��]~��q�a��P�ɳ?r�݄-�ʉkE��y��*O�͉Wc,�pP&tB�򌘣v�C�]�br�Aڵhf:Hw,�ڪHF�ܚگ� `��Q�r�ZQ��3FC��τ����m�6�򄥋�k�E�f�R{�SPqɬ���g�|��C�Ѐ]@��L��~9��������H'ĸA[�A� ����dZDēe���ݪeY_N�_���8�c����ώWM��X��s�r9�%�_�Q8�"L�xG���{�\�6`.�Q2wFU�ߨ��_O�HsNa�K�����2u?��$P$a������{H���f�R�0ݦ܏EH}� ������#���<-�7!KCWG+�+�)�'��о��=�S�u���s+��JE�1�%r���ƕ�����8�;��1Xh�|^D�H�v�/�m�e��3�,��<��FIl��Q}$�Y��zHgI���{}ma�_9�fY)��>ި�#���&����r�����������!���)I��5N�a�I����w�Ir�3C�
���4�t\bl.ϰ���ݝ"zb��qS�}�������^=�(��:��i]`<>.��C���V�RY�uB�O�?=��H�L�*�u��k���&̌j�U�*�������"o��
�o�O��&f��t��Pu��G��!�l��Ϥ��A��f3�319�a��4?�ʴ�#����l���B�-��\ł�-����*�\��=<U,�?�<�!\�l�4)P~���?����U���S�&��&Q���ZDs�P���������X�ޙ��VW�Ư~��]���ʪ&ۢ��S�,� +��fr��9���w�j'����f��X?��S���z��Z+�, �ڈ����� �ca&OE�l���d}��������R�v���ϻsï�s�e{%��������� ol�����p#7�Ì�jҝ̗��l�==�ɓ����~�/���8�}xu~�t~��JE�:DU�����x�"z|� ���&�=�C�LA��M���w�j�_���b��ɥk�������^&	 �{[���?���?�����{A)�qʮ�R?*8--� :��4L�.u_����'��>K?w�h�A=S�>6�7�m/d;u�y�����v����kǎ��m�p<�|���xs�I�lc��6�Ǚ|S��|Zd���J���*Pi��Ɋ9#����#vd���&l�@G   :��+ "�JFw[�цR�����*��{�KF%a3}O�(��a h1鹅��*{OF6�l�:L�6��ܭ$��-���[FP7���	�w�ʹ8��RL\a'|x��&��X���ʠvR���,[�q���c��j�q�Q��~����BYHe_C,p8�AVh\�y�xq( 0�ܝ�m8���N��6�goyޝ�&ag2��~ӹF%�b�[2>E([o��]w;ㇱ~����Y����չ�3�;+E���Ό�m�L�qw��cc��7�om�s"�˙W�i�/J���:�}�,�l��]Z�5�S6���ͳ
`Ȧ��d,Hv�������Ü&�Ӊ����9on�Z_!�O��t�5�c��'�V���s��\���5��%g�����u�lI�C&�LC�R��EwV�h���;r��y�k����|���<.���3��-�'�<8Ǒ��MF�\�C[1�IV�-^~��ŧ9
�,&-��4�p���������J��w�;V�.�(���Og۲������}(>���s^�~�.cW#��m=:�ݢ����5�/�bg����E� �9PH1�A�<1in��	N[�ҌS�>dU�Iнʓ�}z���K8�#Y�����:��\W��~��}�	�|g�]�,��p�
ϻ�7:��k�C�<�-�c
���1s0�P��8)h�2���i`�q�M�����i5۩���1ocM5��T�\(6w�n-s��#��j����y4���v�&�x���P�i��E�Pa����H΃��GO �	�ueg�:Z�F��"T�a	����|���,��;�1��{Cs;��x�o�{���mS�2~J���K�4��|!���2Իds�|[yޘ#�W +��TE�V1�N?�������0��Jc��!K�q5�
5�JJ�� Pl��(���Gr\&��Ab�9�.Yw�'YƄ����xg	Y��y\p�Q�w{��N�r){�7�<=@w��G��BypU;Ǥ��0�|޺�����;(@�@z���[�p��1X�?|�4��;�s2I��m���.z��fu	�u]o|��1��k<�g��^�,�`!ʜ����4�؁d�}2Y��q
���5x�w۵����������};H��6�UF�u�#ށ�^�/�R�̐x����Z���>u�5��Ơ��+�WT�>b^|-�Ӿpc^��`����n�2��M�Ĺ��YU��\.�82u�A5��
_�A���-�s���PiP/h������,nS�������b�F�9j�'4��.�oa3�M2+3�����1�؈S*U�3����xz�Y�\`���9l(K���n�[&�ی����^I��M�o���M��GUs�������ɫ�F2}#,�I�m���\��b�h^Q��骶w���XGrα�'7���v�s��� �3�{o�c�&W��&-	���5��nG�r�����Ֆ�:,U��~��k4�J���b$��H�>����JK���GsX�o$�=�eӅ"d�d@E�Y`c��3t�ې��N}3�b�%dxS��3���ٻ�wC��'r?���<jC7S�`�3���Gy��4�n��>���8�{�ڟ;$���yG�Q��t(�����{u�ٳ�T�G��ʘ��k{L��y��M�l8����X�"O�=�Oe�;�q\���u�_��W^�h@׭������ӓ�����������/�'u��K�Ө� `������$�E��<�2�AP~n���<Y�ا^f ����f�x+ 'N�$���6�D�� "7r8i�N3������@,䰝b|#���c\��@��l�0<�>�sTv�8 bK�v� ٪0��6���Y�)z��Б�����!%9ڟeRaD�e���Bơ�� �|���:�:����ᔃ�l>y���+�կ�FK$�؛g�N �����fν.4M(�@��;��SC:έ�u���ݽ*�  ��IDAT�;��%2�W�& 3Uc"�Dd��h:mW��ZǙGn|���F�&�΂M�D�fV���g2�'���^{��&ǣ�?���$���h8�4�!lh�og�����T6wsYG�1ï�s��t�|��<���UAbw&�J6옷}5�A`s��f' ���8���ĉ�|i9�p�w�i*�X���N�p�T�����@6����0 �)#�5��_6xՀ���cF[���j����6^wJ�|0��2��4�8�W�g�$v�S��Ժ35g�C�3����G4|_�p�^��x��$�>26�n��p�[7R8���GO�?�D����!����FX̯�Iv��}6����T�oq<��w,$�_�!��_$]����I�wa{�s/!o�y��P�E�-�SV��˙�r�H��x.K)�E?�P�e�<|GM<������X�\�Ad�ۋS����~8�םH�39M��H�1���UK`��~��1g�ĦeM�yi���G.�Y����.�$eH߉�N�w��~X�9��9����Y$�ªE��g̖5�rcj�x��\���lo9 xq-k��!;YF� �_m�^�r��C�a�8�T\^`�-dF�a����p�/�F����܄#{wl0��2U&�o�^�3�g���q3�<�؜��l�\&���վM���Y���R� �G�
�5�a|��Ǵ�>$�N~������6^�H�p�4�n�M�4�����Wm���0�}8l�G��}&GrE�i�S��k>D(��3���'b�t��`X[�·��H��i~g|rp�0�Kr�,���	�������>@V��G�D8����i����L3�k���7c�QzAs!ټ�c.� \A�/��W�Sީ���@l1隬y���|�pT��**!`L�x�Zw~Js%>���ez�<����1������4���9��*�#y5ڤ���'�0$���;y�7�V=�������Z[�V�w)@����~X��qS�� s!s�q"K��_�FN�&B��_��*5N�Z��/�v�x!l$H��֋9�������΀��Z�?��er�Bu�C��d�c���t����';`���X�^��"ЄO�'�QZs�3A�`��f�w"���[|ƿbm!�(v�B�o��1��֖]ܐ-����#X��P�g^8�}�ǈ��P��#�L/~����0D;�f������ix,��:J��'������$n)��ߩ����Zg���V�W�[A��晼Q����d�-�������|�8n�F�}�z���S�҅��X�pW+���z�Nػ��f|v q�O���m���V�5�z���L�$;��wΦX[6��Dr�\��I���M�_�_�=���[�:�����t�3��{7�A���/�/��ֵ���Ie ��cX��8f	�fX��Wqم�V_��:4��<>�oY�=
A1�ʣi�uJ���F �����j\z$ݝ���C�;�˔'�$N�{NUeh�
*Ln5�[C�k?���e�Ę�ROF�,z�aY>
hc��z�Oq�[�g�'�����ϯ�k��_��<|(�FD"����������MW �l;�o���������l/��w���,�`���iD��D(vZ��LU��	:�"se�RyA3���
4 ���.�L"M���\Tuج����Yc} S?�ئn��@f#k�l4z��`��7I)�������w4Z�ۥ�Q���ѰT:��������% �e��B� ~Ow��PV��N8�i<��='�0��}w�6|��+�ID��0�D�1�}Fn���?���	<�ߙ1d�MS����R(����MT*�D'0�i���|�.5`�1��@�n΄];�)�� |��M�Ԣ�:�X>�HA�A�Ssóh�$���&���Ham�85 l�
e�`���S�6��D߃v b�ػ����ݳ{��U?w�v��VK�L����]�M3��jLQZ��?�]=x<��s�X�LD��:зF�!=��KD���g���B�s�@[A|��~�3����0��t�Kµ������'d(a^"���������Y.�n�~�='���\ۄnT��g��y��I���������8t�e2�y�^�Q��:wD$_i��遾$6��N8&tW@��^-�Cf0�=��u�H/J8krT���ځ�yO��O��D�jԈ�X��}qp�9�xPˆ%c�
�ԥ��I�k&I�f36ټ��U������X#�R����> �*��9�ҧ�Lu�����3R���v�0@%�X?��Z��^L�q��/r\1kN Sր��G`X��i��=��wT��3XW�[$���0۷@�Q�0+���Z$ua�0�̲������;���|�
b	B��9�ugRA��u���1�A�k�i�����hj���J���D�[�º}���HWzT���X]�� �~��7Z��z%���6�=v��w�x��H��tC)eK�ܝg6�W�@���#�Gi�L��1hHJu�y\��\W�7�ǻ��j�8J���;�؉V&�5����s8�ն��g��uR��Â��a[��#�i�_����X�Y�>>p���L���|J-�;H���oF���D�(��bN&�vLP$ TG�U
�JV�P/GX�N�-�_`�eN�U�1�X�E���7�-H�A2�5����^տ��:�w�bt����	�w��o$�@���q�;�ey;�B���u�z;�I�th��S���~�K��'G_��K{�y<��X�,���Low �Υ>ݮ>}����Q#P�.=�|��E�xʹE�F"c�5�������G��[�;Q`>s�8��˵R��}��ڒ��}��d���Q��S�����I�B���tg;'�tI+`��k��,Q`ڛm����UV��2P�+����D��3���q����.SdM�	���B }�׆�z3�W��;��546��얅mL".��Ebh��#�B�^T����G1ZTп��s8��/���|O��>bKhQ/GB�lޛY�L2�k!L��>i��s��'M�aA�=��6�5��irD���m#��T']�V=g�ù���5;^�X��n��ɨ����l����Z֚�n#_?�NK�,�U�W�.����%|���`,�m�Ϥ;�����k�u8�Sr녌���D�1��>d~���E���)�0�o��+��{'�������d<Tf5�����d��ۛ?��ݩښjf��m7ٶوm=�G��U��xᓘ�b%d(�}\S!�Tl�#�R� ��GX˫�ꍿ�?����7��ӿ�/��w�<y��o�y:��ʵ�_���u�_�g� ��ß���7��'�k�ܾ��c9���]7VA�;����@��Pz��n���p�`g��A3xt��4��X�	S��n�n�{�Wu�k��Qr="�t���5����i�mu�hR�ߊU��ӥ��R�s�)���l̍@R���]��IJA��?�ryϮ��H K雕=N�?���R'J3��Н I
����Q�Y�pؘA4� �gF�O�4�OxwvZĽ
:���F��N�+3"�IБ� ʋ(�:��d���y:�6�6T)0�>5|�$��7�O�A=���jƧ�Ap�jz�%S��Ш�X��V��el�0͗�F3�d�/�m8����<�|�4±E7V�*��,)�^XMU7�%�ظ��ǥg�w�8`[�b��羦4C52������5�Z��v?L ���}�_��:�?5�D�N���5 ��?�;�IR|F�4vPm0:{w�0_u��n0���K��`%��r���EF��f#�������X��|����p�.�$�f�t2�cL��I�Y�����`옺�r�S{�J�4�r1��pde�u�&�������N_�r�T�x-����x׋�ؙN��.s�v��i��;�2���f89y��k��X����mV/�u[C.Ww�t��q8�X�aaB����gv��-�/�\�/��k�nmqY~\s�=�`W�"X���y�:d��ㅃ@�[����0e�H����`F���$�)Xl�t���b��C�t���S�� |Ȋkc�������*_���o����LӶܡ��Lܥ'�}�v�"C�B�����Z5iW�r���t3cK*��dQ�ˉ��ĶB`��jr'*p�|���sd��l�I��'$���1�O�>L�_����;ovS�`��Ε��S��� �;~��b<ں�3uVڄ �AI��z��	_6C�&}�Ռm�%�k\s�I�nV�Z�iir���Ԁ'��M0�bI;Ū$U�p���9��`/dо��8O�e-*�4G�f`�w×aJ�2�v4u�&�������j3�Aw�[Z�L�hˊ�<�.�����׹�W��Z��z�N�r:��psc��bn��_�?�K><��,T_c+�I��v�rJ�C�?��%»���Qͪ���w��;eE�tx�OZ�4!��qHNV�k�LN�]��E'�.����7a����u��5����BvE��&��﵏��AT|��/k������(�}��c�;���[��Ɏ$틀��݄�@����轛��e@��l��n�;a;]O
����vl��8.���aCaF0L���X�^]� XTE�R�d�ĸ]� ��V��� �]L��.�&G�\�����`,!���t_<��I|n��<_���}��Jƛ��Q��֭��z�_Bm9�s��8�T���%��:O'O�K��:X���=�}�	= �2F���^"0|s�u��H��!4>�~�>�d�A�C������)[��;n���)�!�����+!@�bV�kXi܊����Ks܁��N�b(��1qؔgzo�^�h�I��̔�`ך������|��d�z2<��6iw?5�["�W�_�7����~�D�c����y���k������AN�'n�p?�JCK�r���e�i?Jߺ�f����mW����<
�:z���c4ś	qy��ې�I_W�<��+����&��ιI_�2����.ؙ�w�xQ��Gؚ�o\�7����÷���z�^����2&�Bî�����T��n6��:��nH�u �ͬi�}$���( ��;F�y�3!��@�#C�ѷ�n��^m1�_a��k&�n\q��h�����c�n�V�)oԇ߼����w��{����;���k2�X�_���u}���' |��Û��ѣV�o޴�ͳؽ�;��,-��Π"���J±�� -���CM`@�4h!�U��0��X@�v7�z��r�wL~VF3s��桗�T!�#.���Z\io5�*;�;w�W���B�L	2�q1Ga���>81�MN����ݵ/r��=��5��(���3 �R .,��`D�:��8�w�qC�#����v�!k�% ]8���nR���@��!�1�ʽ�bAT�l�b���A����g7��Log`}��m�g��Xt�?���O���x@s�#,����nA��:2�Á�6�wvKd�Gy�ՙe��\�`]�D$��֫�;����Zm]�d���w� �J��E�x�	�G[O#�g�og��g��{�Qbkf:5m{]=�ł�؄a��+3�f;�����8ϡ��}�Sw.P��,�7��OFڍ�`j�*��V��HбH���g�߃�l�ʲ������X;�p?wm�B9ɑ#k�S{�J�sFh�ݜ
hs���6�J�=��fTt�GN����:Y�����%��fuvs۠e�)h��c;������i*Wh�}bGuP��'.K��3h?�*u�EPl�}�@E!���(aΕ�`����@��U^�v[���л`���-���9Ü�Y��$v�c��N��a���y�����}�YN�oA�濛��1u`�Lv�]���,ϰ�������߷��p�����zHv|��ݸ����qe7]gо���v�88�����jF�����I&����o�/0N��_}��x|2tu�d3$�fG=��������{[�Cƞ����r�5�鎲����0�")�� Д�~�_kg�U��pC�n�5���w������9�N&[�SG>8������N�I%q�vc;1Sғ��
��Ƙ�v�%�c|�Nɍ&^j_���nN�C�V��l�+�l�}J�)ț!�j�[g8�e���A�y:Z��3){��xy8�9�ŝ�}��X�`Υ��5CN�[���L;���3:T��G�Msv<�Wr�8��N�$��
�C6^q[%�+�\%Ɉ����Gz�����h{s�s���t���d�3�@:���4�+0R��T�{�lT|����<t���ݱ�5��k��Ȳ>dS�_���+ż�:[���5���0�F�7�sJ;�-���c���r�zo�c_c��c��5�b�*�ܻ���
Vg~��{Q�D�
Y�1���Ph����W.ƞ�eg;�I�-�c~�>6�������Y����[$�A����������g�,�x�W��zC��tlp��U�'�Ko��`�
��&���i��y����ErR�c��B��������	/���9�?딸 �@�.��b�Ϡ�P�Q\�U�`��ܩ��yq�}��Ǧ��a�>9��1�GB9|Y_]�U�>;�qi߇nm^n�>�g�r[n����������LZ<�S-��̧?eoz�Hm@��U:O���@��ѷ�u^���%���n��E�QoI�yIKѼF�[�G=�s/�Q�E��خ]��ȯ�?�^���CōF_ldC�� ?�A)����6��`SJY�@�1ۆ��)���xz�&A��[�wk���)�a:U�o����_�Ty��ٹ���U ��=:�d{�)9�ͻ�u�x�)�G$�y�1������x!�.��@�nn#ߡuê_T���j����!�ÿ�&t{a��!�Ú����K�.�*��r� Q�>Y�H��}س�U�&o�f>�����x`T�xӦ�!�"�u�����r��c��:+���7J�0�j�����Y�Ħ�&BsS/��d�&1������<���r�������k?��O�z��w_??��_���u}���' �����6���w��,�cw�^����5@ŁR���!|��0M��Y�P�Z�g��EAE'C�b�C��Cp���қ��gZ٥��G
C�j�d���nt�G�
��� 9 ��x5v\��v��R��b��(� ��5�:�4��M1ο-L�{��ǻVb��"����c��c?-l���ͨ�c����}0���F�E8x��;0`8��cp,:��9s{1�[�
��3�u�-�,_�Vy]�{�n��;�����oo��`�������ϝ� ��w��<���,0��S5�I��P�ǒ=�R�v܂e�v�/9�5����U�Q��Ù3��tG�g��r��( �s�@=Wҍ���F4�]��t��˧�_ru�(Ȍ�r ^Z��N�{���b
8q�m9?ۊe�?;mo#q�|�V���>w�je�A���N�V����t���˗�œ/��/U�߻_�!��\d&����Z���h�[��5�U��j�G��![+�a�p/��3{Q�{�Y��8��{�5�]�N�N�Hl�q_�
}o�!lLU���^��t������]i�B�ł�3��zR���.��N�5>�i��~�vv0�#���9�S���	����4�s��Q�EE_4�*>O:f����U�"N�p�Q/K��+L|ނF��Z��.�Џ� \&�y��2��:ذw�>��̃p��eTc4HZ�X�Ƨ=xW��{�ߘh�W���� ����~S�V�D�]�_�P����Vzʉ�4г��ٰ�	��w)-�˕)f5F&w�Ǚ��&(V|�GA�/�S|��_W�4#~�>C�O���[5�?Ɗ�T���%��y[B%��B�G��7�b� �[2*�G�N�O>���^x�g�,aX�tTab.
�H�4ͫ9�E<Ac�ܻV�P��`Ni�D�%١,tY�[��"�h�\0M��%�w����m?�;���O��w�������<�O���޻Pno�r��2�:����f�@Ͼ��Ng�qs{;�g�Nz�;�S�^�bǰ;^�8`�+��=��sЇ�Ü�]�g)�Dp���s3m'�(����X�n3Pt��x��oc�{b����5�PgR�%��+Vh��8�m�B;�F���Mw;OgA<DP�'�@��~���S�n��M��g�j�=�7�3Όo�21�؆�6qD��͎�:�r��<{��~��������~6�l�S�:�m7[b����
���˨��_�ǈj1HX;���-����B.��V�V�B;H�f1Y�[[����v�v��"���u�>������&�\�a�}����iNr]I����8`%=�^���ֶ�N)~��MB~���5�N'���E��a[��\#�t<�8�a� Ыͤ�Y��C�� c�������x-p/���ʟH��;ÛO��b�+dZ���<�xGpqqGY`����]�"�A��H�;�����5�� ͗�Kz�oׇ����um��`�c�i�		F;1?Ǝ��]R|��l~Ǉ�>x���N�e��~_�(����l�rYq�%�c��d�" �BѢ}�X������aլ��G�E�����������A'�s[�<Nح��1/z�?������IZ��Է�ԘkG~�RS/�Nc�Y�4��?c�L�����H~�����|�7���G�m�����>���3�o�X��?E�T�TNl�� ����W���ݶ>�����K�v�uh~㶛r����(c���iV��l���䌀��'w��3q��O&�
�Ȩ64z}xQeaaYU���s�¯4�U��M��,�y<3����w�i�V:�D�U�A�_6��r��r�1����6=�]wk�����g`0O�i�4���B�k?vF��x�ӳ�~|��|��G��y���t;���]�~�ͪ���|Dz��8��m�h!�j<7��$�Y�^�ӻ\Kt�g�ӓ�� O]���P�w�< ���=�HB����L�q0����H
:�k��BNy�d��5Ya��7�Y` ַ᷽��JB7;v$�*�DK�6! �U1���}��*�#H�n��;�F*��B��tK����2���'t�t�ި2ױ<t�on�����k9>U�a���h��8[�������+�o:��z���;?��W�o=����/^���?�c�d��*��+���ʥ��I���@0���������%Ja3̇���X�2��: � 5�_UlB�릝P�r�U���mm436�-����ϡ�l����;пqE)�T]�ci��qo��&��΍����wԢ;��'^�V�x��W�Ky�&Jڍ1mhĥ���kQ��̱���h��x�V��R�g���T	��u����k�f���6v&b%��+�d6�>�o�׿���_�W�_���?�nO����a�q�Ӓ�e��m0�K�ن��5}wM-�v�F�	:�?���׶d���\�|ݪz����W���m��d���[����!&�H�� K`�%{�$&�B��G�H�e�E��v�n����]��s�^+���\���6R!!�U�u��{�\������HG̘L0B�9������F��.$=�52$�3d@��<3Yi�����M( �D�	�B����9�Ssw�f����n(����m������ߍ�m���gј#��ޔ絼���.أ�@��n �Y/��>������������ʷܷ��o�IN�@���`/Q��JJ#�܍��`j�,.t6ɚȐN2&
�?���`��+��M� `�;)8���A�o��rC�-ك�KD�$�e�O�l8N�I�A��	�X��G:���j�r����-!����t�/�E��/�'�mvJ�~@yB2�ʬy�'��wH�4�yL�]���f����Y�?�Я�����Ei�3ݭ��B�BO�`w~��l�K�'�L�aw4n3m����\�IT���F-+���H���u���z/��Ei̠g�$�&�T�g:�$����;#�����z�=�5�%�X���/���;�Ȃ�A?��1]�WY��ďd.O�/�	$��09.��k�q�6kw��QX��6�e+#.��%�SK��\���~�|���_k8bMo"5';���r�ҐPm����@�1uҹ��h���i��7ʮ*�%�G�Ue[-L�R�!7su]���O�f����ʭͻ�z��oz�Vƚ2
W�V�-��w>���?�g���o��Gw�wk�'�]���r]ֱ-��<�*h`Q�˗�(�B�v�l��4�
��I0��e�����Tfς�b�����p�|Yu!�m�F��H�]G���m[b����U-�F��zְ%sT�B҅R[��5c@}$���-A��j���(�Pm����­�F����d�nZ�}�/�>�U���ߍ}sî]Pj�*��Q�D@�D��;&߇���������������Ͼ�{K�kY�U /'�A]�	1dkar���ɽpR���?$�S:�|��B+��gB�%}�nIETb��J�L�>?�{���U�cU�1~	��χ�:��ֿl-���/������T�}�����Q̙e���H����9>����������MG���<��,�����j�G���ާy��O�����;��qQ�H!X ������x�A޹�~��*��[�G�Ŕ�5T�ry�v3�F��A���=c,J�=�|���Uc�����TWk@5�i�h��QR�{Z�6���>��`.�9r�N<Y�\tT&1 ���^Mc����!h�~���c��z�7p;f���]�QM'���Hn~?ǎ�`Ʊ%R�Ъ��vA����}N䄜��� s��Y̵3҄���ح{麼�b�5���Fwg�����s���m���(�p,蔯f����#�?v��1fv?����F�{c�ۚ��7*����w�CqLW�7 �ڰ�~�G�éo.��?�����_�g���]�}�p����ӎ7֑����7�쭟�w�0�^S59�	Di}�e�Pg��0\$����8�D�x��0=�]��`�6���Nv�B����V�T3d�?��e6���`;��nVw@��æo@��ͻc0/��8A��tl�"�������r�Γ%L��l#�y��������w�Q���+L�lXG�M]5�纒����ҞF����]>���_�����}~���JM�1�3.!�x�sW������m�n���b����W�_�5���>�H��6�G��p��=�%�m�I��=� y��,����b�@�b.G���<T���"�~��9�-"0�'��M���-��Uf4]�H6SN�7"u����_�XrF'8�]>a-��w���ѫ�9�w-`���������v>��X�N4���DQ��Mry$�S;SY�z}|h��?��/�����Ԟ�����r�\/�t}�	 �����ږ������ʏ�������Oo駶�p��؃����g㎒`�rM�7 �U�vG��1��j�/�{��
1{�VEG���)�s�1�[��D��Z3���v��^UģrAK2{6flG��BK����� 6RE2tM�fԐ�:��8��ܑ$c��˺���#JT�7�5�1w��I��!Ŭ;V)���{
���\&�F8��,eu~H�;*$$�
c�����8t́@юn�;�7B�=b�f7�g:��vl���mG�]@�}]�{�]�'~�/޾����?��n-���v��L��h��^��,\*^��/�`R�KS톡��e�a�KKH�jݜB
;q�{`g�I@��	�$�KT�/�٧���:`���&ۨ Jfa痽R�W^�-j���m��Wf^�7�������|�"�bS�	Rl�qt���q�b8NF6����4�^��.��v����hzZ��|�ܽ�y|�������@���i����]; ���Vt�%�gP��!�k��ɢڜ`��]ʐ˘c�=�3_jk�C ;!�S�\�mJz2���{��ԩ�%9¬�X$oe�dW�;�s�m��pz�T�������Y�@����l��yp)�'���V��wg��vF��)H��:6�����3-�;���xw}��GiL�q�]��/ꨂ ��ĺ�`qv�e������<�)�˱[�[I|���|9���4t^�d���,����9#"T��#�Sm��^w����!���n72X�`�l%��N��
=Z\�Xrh�:"�����"�<�њ��xn�#F2��4O�Fu��r�!G�S�p,��!r-�MZ)��|^�v�8	�u�}�F�*H���t�e:!���Pg������-��d��	�H�+���cN߉�l����D"�2�%#�h{8��:@J4�:<d�B��F��(k�Cp�5�d����nr�OX���kЃ���
8UX����ݏ*㤟͎.�*�F���ݮ?s���߻�����ݥ��`���}����:��&�~Ƅ�L���C� #�D��?=��,E�Xl��k��K�t��V1�ړ���̈́zU��p���+�Y�Z8+V�X�����#�_K2� e������G�Č 97.�˭����ﾐ��n����\�|$Pd��қ�<�w��/8�}��'�fo��Wm��es5��B�VI�Y���uk�K+;�{�Q^������Թ�1�m�*�!gl�jqD�[F��� y��m��E�����\�Y�z战���K���堷ݑ ��eH�#���oM������zx���<c���Z:l%|�@���G�LAI�#G� ���g(�b��@��΄CSU�!��ݢ�̓�E�;���b���o��)XGц�0$t�L�7�2�N����uio� �ʜFH�����(��A`�x֜�'8�g���׀Ж9|&"	��7���f <���=Q��8������*���ǹA�V�`7_����dq[�v����f���&�;>r���1k�p�va�1D����a=`��<��� �m)�X�G��d!�Œ����}ѣ)ɗl,�ŭ�43v0<.����r��3j�p$f�dE��Q�RN\	��|v�C���a��!�����̎"�Ӽ��s�m���3��������c�>+��j%���9h���|�Q6��N�;��Ї|g�?������GK������[o�e �����vz�����k������<;�:��#��|���؆��ZoC��/0��y@bArQ,��[�}픳�B!6�-����ma ئ�U}j�&����i�la�q�ڏ#/fRӞ0�%��ʫ<��Fk ɦ�6���ٚ:��2��VW���e�;1$^��N��;�����GB�8TJ���M���CE�v7U����=�v7�\[������]=�Q���y�H�P6��`������z����0�j/'���0�#)&|8��BwA�ਤ8jI���b��V�~�Y�~r��&?��Q��X{�ol�G�����>�C��c���a�9�̄cx���>��^7Ǚ�)��c�1�=�z}���:�?�;ب|� ��Q��S���{�������h�v�b ͭ_ن׻�+�f�4�M�p6����G�;q�gz؋��m$�4z�����c���?���[�^��W�[
k��z�^�����kO ��m7���?���_������?���{<��[O;*���V�Æ��Z��,7�p6��_2y�E��,�E1�(;�MC����ǅLPo|�4�A%��ֆ@\��{����

�;R��P�ˋ�1!{}���2v�l�h�q��FK7%�;3�;F��ޟlLf�EI�r�Y���[��6,��y}\IR�pV�/�kɎ� �蓚�e�����X##Oi�9ኾ�3O[Ӡ�a�� `{}'-H`�%[I��IV�9����޶Z��>n������V���O�o���c����M��fT�盛Լ��p�c�X��!��6��YЛ�0~�X�H��h�(��C'�ͦ��'��c{6�r{t�=_��W�e�N�BI��n�����]�w�m����=Ms��o�} ��i�@7���.3�ٛ��o����?�۟��[:ib ���hs�M��N�"sB|�+��7�ޭ�^�g���	�&e�e
w�"�,�I*MA���H<�[��͍'7C6�\2��Q�q���s����G��弲�T^�Q#UvE5�y���脒�;�[bK�PǱ�ZA��|�u��\V��y"B\�o*�k�9[��[��&��Jj��T�������0���
粲G���g�;���7{�y�����)�%N_�ʆ�a5�w�#"�m�ww�ޜ,��t'�y��熤�;R[����W��uc�K�?�w+ikH"�o����<3�c��6��&��4AK�,=y�)�u;{�-;�/�XO���%=iN��Y#x��[f�H+�\������Ө!QBu�8@�n�p���\9�K����z�9�e�#�m,��j��ng�� ��zP���Ҷ��<�َ�1�g��+)����<A�4���}36���^Z�5KNP�����r��v||���N�����׃�@��q|���j?x��Dbº�>����%�j.��-xc| %�v���uY&t%s�٘�icխlγ�!�.6��~�4�Io[�FÎ�`ӂ�I����L�s��ī'7��`�Z�۝}�n�y��K������oSm�wm�q^��TVن!^P�����7ͺ2�8��(6[hi��;ۧ&ٔt�^���7]㸴>Xk컏�����~�NǛ�;�|?���V���,��������������Ne�%*t_F�u̛8�G2�-F;y+�J2�~߾�N�5yj�c��0�lw�������������6�u��xx��@�ڋ��o���G��UMH7���ٝ~�i"�W�Q��rg�]k6��z&�`�g�G�G�a���F ����<�"�˃�nkյ+�NŹ鎲�{����#�`�ʀmM���y����X{�eS�ǋ�^5+�Q �lP68����U�ĳ��rEu�8�^��G����K%�Dy�)�F"�@��Y�;o���,��锇�ք�j�0,�p����G��P1]ًᎌC�f�y�k2,�^G4w��D����^�/�cǆ�n��sж5��	uߘ�UW7K��1��/ ���ѓd��V�	]����Tji5s1��/�fZK�2�6��U�/������C�}^�^C�^oU,f^���g"!�m9ϵ�@����y�Wp�������%'����[I��� �1XA_.	/K�L9�D�jP}���uXJ"K6��YA j�1@($�=�/uǳ��7��R�l�o�4���l�ðo�	����dk�T{�9���M5�'%/S��V�$[_��'hMsr7h�e��E�a9��֗T��/&A+��W��R	e�h�y*��z��~��O�z���r�[�����R~T�]n�Õ��m�w��v��uoJ�Ʃ�����.~����>��^��>��ޝ�~���V�'Gf�J��QJ���>J�Θ눳p)uFPم�*����0,�dLQ�~���*��Y��8F�޿�ԆR%����b��~��Π�Z�����.dc�b��-��'n|��x�����~�a����a������:1��W�-��ێ���ݼ]�]�V.�~�<����������ީl���RB�I��������!5�����P�6��.��d��T����%���7�0|-#V�c�Jl:;����M�˚�}��M�^Ӥ��-���1A��*�4Aϓm4~DBzN�>�r2� �>�慃;��D�!]w������&�D:��lhv�%5:�i�]TZӣT�xd;j�B7�m�y��	u�I��y��B@��s���њ�dYRͨ_8���|i�5q��r#4�|mI�69�*�#��f��O��O��_�����N'�����K����;���z�^��ˮ�5����m9��,�懿����������^��G)���;���9�' �vW��,��\J�wdbG�|�(��>�MT�t��N��hw����`�6,/̄}��3���{�m8]���P�P.��$ʒ2���׶�t⤕����Ϟr�淜C��g����\���
͹��.fT؋P`] 8$�LJr�R�>~7��q��R"ALs���fP��%�y��y�8J��߅R�paN8��4��z]�[K�{�J����v���}<-�O�w}2|�����\̀��#;}�����n2;�EW���Xp*G`<����O��Yw�8��!�/M���F�ٟ%*h�ǻ�C������ �Ŀ�w��5v�o^�n��ګQS�gݍ�!;�s�����W�4ʿ�S���Fuq>��è���F��$<ҡ�Q4��q��Rk]n���v�H�0�t�餎�Bm���/䆁�Ql.Jl�9p��n8^e����W�X�%&���A�h���:" %�ʨ�ڎYw��Y�V���Zv1���B��N88t�ٛ��t��66 8�}�H�!�n��S�NP�7��r�t��G��C�Z����c��±�r�G����Fo�J=���Bi0/\���9��	DLIoq�p��d���Su�?8����L򖐤F�l������*��EIub��fd~�
?��<�v"gz��d�96#�X�Qu����s�SwV�6e�-�w�*U���z� ��Ɠ�X�>@�:v�1���ג���`}`Nĸ��K�k@鸥u�Џ�N>��8.a!0I�ϛ�Y�����H��x����T\C��eYk�5gOG�6ߐuٱ�� �`%N�%Js�a�wиcf|�_�Xh�@��F����6"�W��2u���d)��F>�8-?��:_���D�)�[M*+&���n��v����٦OL��9�V�]rP����{��!7/M������';�~w��j_��>�?��X��b���a���ё�E�{zKo�=��C
|���D�6v�ܒ~��A�#�G��Q������[NW�?�}~�w>�g朶������ts�O�3���v��{�;�)Ļ@���3��	cl*�ַu�r��a=է��wi6���fГ�:��$,�
~��w���V��l rO �8���"]��X�~�:(QA�$
�l��Np$Z���daG��.�5 m	s 	M�� ���C�2L����"���dB�"�S�����(��l}��hO�5�OIeھ����*be�j�K����.�*Y.S�H����wn[�X�{����P;Kez�뉘ר��>|�`�X�p��~+n��D�\<9Hw�;ΤX���n�����
��F����
���I�o�o��EpZ��'$�@� 69�=�dS��&J"YR�%��R(��\�e�u�9��G���ǖyu���gI����7���{��#��$O�#��icIɳ��-W���Ԅ3�B������_MR��D��ʣ���J�x7�2���'�9�#ǰYn��z���t����(�In_�"$���c3m�7��o�2��0[��h4���F�w��!����<��H���3������$_�`!���.��:���]��R��6U��۹\�H<�f�v��������T�Ǖ��������^Gp���.���.��+��W-����3�y���H x��.I 4�{?Kj�:|AV�yv��ޒ��}�<]}��`%�ku��e|v� �t/O�Ս�}j*���ʱ-I)Ys�r�QV���B߱��M�l�ϖ�G[8K��c�K������w8K��F�ٟ|g�W�wk�wul~0o�QH�&�QL�?����d�>�O��;��\�e$oK+��nm5=7��M*���U(-���dw�$�%�F-M�?��T�&	���Sw{�I>ٰe(��d���Wx	��1|�8E�E�|��)�,��+(�)Y���OÎAT�c����2�*dZbؚ nu��E��~�����aG �Z�;M��4�1�Ղ�G�ns� ~}{�b��1�ѫ��ű�^���)���&��
��6��}��b#b1ʐ�{ty%̌�s�_\q�ez�]��R|ٗۥ��g�7�ԏ[-_}������z�~���  ׶I
ݛ���/_ݿ:Wz�u�V�p+�(�r2g��(��GF�JqF%����:ڐ {��L��%�²��`�Ȧg�/�,({�$�nA���I�P쐴7�8�+ێ��i���̤%�Ls1��Rw��	��c��U�vM�1��]���Rr+�3�N$@���� I������3���t8��P�2��0=Ϊ����Qz��,N���)C�yknjmV�'9Ip^.�`l�.H����Hi�,h�
�ǹdc3���y��T�����i���^m��Z6�b��j�R 	 D,��3�@8��U؂u@� %��������͘QP68��y��W��q�!�������vx&?'�ڟQ��aC���5Gj����;{��3��w8��x� �,&<�G��|!�n���un��Ǻ��gK۶���'���Zm�xw��5gWB�q�X�p����v3�c�_�vt��Ț�b=A7(C(G	J�g]3pĐ�cdVG�}#��n/�q�6��� �ϲ����
[� ���ex����̆��M�����>��+}��Sv�Q�D�d��VV*9�Y�V�;��%�׺�<��TBr���lW���l���)�)���< &m�m����.��)v���'X-|�"LM2�22�S	P�t�\7�Tm�[�8X[�D:���s��F�yI�GE��wE�T�_�R���MR���A'��S�o�.1��ϋ{c���V�35cB�~�������~�GӢ/T|�[8����4����}}��{r��;I�#^Ε�z�'ٺG
5K��H���#�� ߵ�#��v :�
k/v��b}��:Hw��;�����p�N)$0��ul{txr�m1�ήva]�#�
��ͥ�k��'w�js�I�ٳƳ���\Z��<'��z���Bu���,��u��6^48��1��M��;ݗe��=݆�}�fB�y�P�V��!�V��J��V��f�ۺ��߾����N\GD��>�l�d'�U3�-�q�Ш�j�7��&����:���Y~�����m�3������m�s�����>��S9�v$��?�����#�\����㧧��1g��S:���֕����˥�����ߧ�˶�����{��}XZ}���]�l_YO��*{�6�]��G����n��.��d�MΥ�q�2֠�����Y��B�i��a�fP�d�j�R��(6}X"X	dS,�:����n�B��V�M����-�����ի2�>l�h"r]!����s��Z%��q���
G-Y��l:��I�"�5L�!�(SC��;��
�&��ǲ��b�-U���o�}�
������x��-tp��g�a��lN�#�t�M|f���lO��ױ��J�s#�܆}�د�D�D�cj�[����1�N��b}�b'`=��!�f��}:��c���P^����Փ%����lu��TM�����થ�&�n�z�F��Mӧ`v�<`e��0�k2��Vf�>���|�\"lHv��
{c����ϻ��d����AG�]+�|jI$�G��<�u�*S�O����q:M�T�Q{9�k`�im'���Vc3k��cP�>�<,0d�=�RT���@��d� 79^���8���>��wz�hW�?*}�1�u����ov��K��G�~�b$�'���-���T��]s˿S_�Ì����~�|���z�g/ΎX�XBW���������|�*��.v3_.:1!��(�}O��7���X0��?m��e�g��H4xj�&^��)��y��,�q|waM��%�w���X+e��DRB��e��>cOk��=��|qs~��26RK�*�T>��""G���1l����M��.z���	2̄���{�t���I���?�����T����#ߣ�B^	]n��Cr��F&�B�ߢ��b��W.8�k~N���裶&��6��զ=�9�W�S|/�9t�ebU�+��k�.��VN��������c� ���:�Cɏ�}09�O����s�/��X+��N�?�%���c�ƚ��T~��o�w#�ӝk>]����Qݽ\/���rM��	 \���~�������}����}�Y�W�E�Z,�܆F�U�q����p>�c�z�;� #5JPNE2n�)�0dr�Q�B	�!�%�Bx���҄��(�m�ڨ^� mF[n�!�<�y�,�j������s�s�r�d����*�����4O�w�s�U�5c� QU��zEn��1�<����
>�C'��q�}[�䖚�?���L�2 ��?�l4��1.qPXo����V�NB���#ey�ۛ�������f�s�ie;�K9�(�U�"y��3u��"ʳ{#`������� R_ ܙ-ύ�������A�m#�^���f�ePȦ`ToE��U�3�����8 $э�^m2��짝;+� �r"�m8�����F6l�*2�����5yF����2u[�l��Z.�3��u;����&��� �0j�ˉ��c� ��� Ƌ�0k���^|	:��9��c3�j�@ws��>�QAT�LkH։]��Ea<	�;�Op"ib�u��i�w�9ʂ5�Y�!� ��������U�2s_�yfBf�/�|]K!��8o�t~�X-�	$�G0Y��/��d� 5^�ɠ@�G�y�f��4n����P��H}��$8�sryvz���K�#���=�I}��:�;<��e���?�#�$�b�ܠ?��#�,�Ž�I�q8��7u�1}!�%󗁂�˶t�9�lD*��~M�#�����x�p48iS���9��B�C����i���eӵ�,��E��Ziqn J�Gg��b�qH7���b�?�'��3t��b4��&��6�G��>��H��D�X�֓_[8��3A9h�ʱ�:m!��t�s��3y� 瀔�=`�Ч��+e�x���!��<��po�O!��ݩ/m)6�ӆCp
1�,V}����������Rd�9����-�c�ɛ��<]v��t�T�ޯk�p�K����r�� ��4��r���`�V�]��O�l_�&l�q�W]L�ϕ��~�9��R��'^	�ɟ��~���f�Ɵ�,��xj���ڏ$ q6���K������G19�������H���?��|y�u=���B��ֹ����8�c��L`	|g0<k\��*ǖ��"�ʤ��.�h����Ǥ��Ě������2ź�&�#��{)���$O�{g���P�8�����&�a�e������>�Ԟ�	%��I�3�H�C'%7�6X��;��C�wS|���1���6�b�}FZ�CC�,�Pq/���8Ǩ��=2z[�ڮf�Fr{��o��[�'��С���TD�~�F��q* �(�o��9g��Tr}�g��0��S����n�B���"'�A�`������NG	s����vP!-��:�{�ʾJ��)���$3���0����9��9���'�z���7����N�-)Y���%��s<�vOw$�Tlj8V��٦`BZ��q��������hi�M����os��0u�/1CzJ��'��ʏ��z]'��A^��r%U�(h �cr��)�b=C�gI]�Ic�4�f�q��"�Y�p<K�� rt�3���:��9prT|�mׯ�&в���������n�[.Ou��M�|����vW�7�;n�,�����g����G:_�㿔m�m[��~��~�O�L��8�;��؏��q�e�{�k��3����1%@�6��]�Rn��Bp�)�/tfĈ[���0�H���h�V�W���������쨮������k����g|�w`@FI�xk�/� XՂ����M*_�r�v����͛����\�)��y@{�%s�.��1(�PX%�2O��l�Ǳ&�[@R�塏�f��!`�����=*u
�V��!C�����]��?Ҥ#���7��|��	����IԦw__6��
	T�e���I$a�ƥBQj;��z
w�ԏ��X��>�6��c��|;��~��l����(��a#�6������9N}s����{�������M,���=������zss�0�r�\/������& XЋonn~������������|^�#В�� �w"O �0�gV
!��w8���!�<�V�
��@
�����o����fƿ;oRP�BM�ąq�8r��呞�� Z6r�Ya+ �V+�߻;u�ad�ݬ�`ΰ���b�FP��d$�����w"�]��`��7k~�(V�����1���0����8�_('�w0�bT[5'�M�=�#�{0�D����swz�O��3�@���3�Qu;�yok�lt��w�\v������}��7��w��j헻��� ����.(�.z<����u?���������e��.���G�C>�>��I���l�4kS�?Gp_�&�@8.`$d�ۘ�yO����O���5���2�v����Ri��7��.N�:��x///���i�E^,��`���/uT 8����V�/ޖ�n�#K��Z*�݂��-�Ca�]�%��"��[��A/ݨg�Ơ��b�,�l��=c�7[�4Nc��(Q6>D]���^r4��S�e�s*�����qQ>����R�@�d1ڢ�4�p�{̓H��������hh�������ȸ���b�8Ι�@�|�A�=1.�E�Z��?G`:v�uC?��;�x�����7ϒ<ѫ��#����{(TB�,������]8���L��y���t�J�L�N�y�N�#�zz\q��1��y��۶�����:֖d%b�w�Z^uד',&�P٠_�x`�w��9�z�ǜ��hǩO�YJ>�p�%E�\-x⳰�/��zd��E�ep��/�6['8�(B/��Q�����񟭂^}�=��P���Uʕ�͇<��t;~d<3v6�Y���w������!��+�}��F���+�?ƚ�[�k>���>��:2����d�$�I[^e/���i((��CW�Zq��*��±��J�cu�tKL0��@7q����	����q�{{9g��?z~,���oQ�O���
�v�O�B?�zk�1u�mT�Gg#l��j�9/��v�R��#S�t�Me��̓étᐵK����8Fv��P�4MR>�+�Kv�(�p)����3g����+�v�P��[���D��3I�	g�m
����2��6^O��o\��e�>�?G �7g���u�e'�y�꼷����ַӎ������g����ڗ�þ���C�����SUʬ��!�������%�sX�k�@0��\�q��W���w��L�ԴB<�!��3�[Uy
S�;O��ɦ>�RଞdF����������!�9�� �+��ְ̔�.;Y�qR#���m@�Ov���3p|�3*֪��n%�U�d��>F�Y�M 1��Oo�y(��-H�Qn�N!�K��{�y�{�ɳb�Ih���'�K�.��s���{�S﹧�װ6z�b-H���;�.�]�$z����C/$��h���cN��������[יGem9v�-%�kM�G����[�ů�U(�qC��lW�c'�9ٌ�U�X�^A��h��ܲS���$��O���&3�&Mk?�1O�a|�~u���`�/��c|�����nKkZ�I����Cџ�̟�c��v��a7�7k�9'�?L���,�LN.�!"�4�	@[߂H��6*��U����MB^oBO��lgl�O�b`z�K̿��$WFO�o��'��y�{~��z����x3L����H+ P{�������u�����0�h�c[F+����7ݤ.y�}�.6������]�?>ρ{;5��&wA�,��ON H~6�Cǟ�7
�5l�O`5�*�)�5���A�����Y-SHa�oU�.��S����io���A��F��V1W�{U��3"B����E�l��|z�����?�����i=jz\�dY�T��	��%�yбӼ���y�w`�"�|<� MJ�Z��	���3��f��ӥ�:O�q%�������eD��ݰ�m-%�!R�9y��˥)% $mxE�w�xon��#��z�n֌c���b.��r���l�Š�v�&�.F�֧cN�?�^�h!���r��\���</���^=4�c������g��NT���>��錘���6/~�a>V�}����������~�g?�y���.�9��e_����z����+ ���^_��_���g~��������"��ze�Hk����C��B�2
@��ɍ+�S@�=@F.���lw\~�NR�Q�%$�ʓ�9�{6�`,�/��;{T=�VE��	X\5� �s��0�?yCۓAZs~b7���JRgo��}��
�q�0V"�[���nn���A����JR�I��ŀ��YD	m�e<+�gdIe�n�22�u���,
���4I�@If�s�@
l,R�6�W��q#�{  a b���y`�p�NZsTd�����R��o���Q����w�߹��W��e���\�u���,��K��z�t:y e�G�K��U(ݺ��{Ø�A{{����F����9EޞN�ڊ��fC��~�@,i��;��u�݊ٗ]���V}j}���83�I�����0xv�.L&�l����}<��h�0r�|ՊE�.�}�Y��^#�LMuYڲ#�z:ɱ��v�>�]~�߬������S�e�v���_�,ruh��f}���a��P�9!���٢���X^Fp�=[$r��:�y+Hka9�6�qZ�{|���#�s��^���AtH��S
�I����T�*���Y?���=�>�֒�a�đ#�+H��0�:C�"����m�n���ƕ������59~pM�T��u�u�h�w��5��6ۢ*�.+\	�O2D�q��*ϋ)����1�ig�J7,�;��ܶ��$���a���'��j�Z����t�o_U�����8��40�;���	�*�a�m������	W�]"�1�5�炓�ı��/�p=<~�E�\����	Yq�i�u�5��Xc'���w�w3�8ΞU�r�6>V[k�{��ΐ`@>w2���
��51��l9��q�J#�G&����M�E؍�l���\8�&vބ�1�qq��r㱥����D=��;7x����a�a�¸)�?A����7D-�+J�۽��������b�3s�Ck��TE�0���!Vx�l~�D#h1�bg?�A������n�R6zzM$wr�$��;��r���8�p�]�+�$J�qUy��Y���:�&�<���3^H�+Pm�y�� lع����g�ݺ��:[i��hY;�������?�Ͽuõ-��ݾ*~a���]N8���t�jAfٖnz_�����sZ�ն��tZDI�������������U0��)��ꂮu��#�m
�{s�;v��<�����kfg�ʒ9좲��,���}�K;��B���;v�S��x�s�`0Um�~�<���W�`�g8E{�R�UF1`�9�n��4B�!ހ;y�C��-�T�N�V���>�0�4F嫵,�c���式�2Nv���w�<~�S��ۿ���ö��Î�ތ,��8^*�!���F�ϐ+���)��Pg%�eD~@WM���&��7bcO��k�#�Eu�$�����k��7��1>ώ����8� =U�XA��@�Ű���c�2���?M��$EY�n�R�VW�@<@)a��X{����9��I���]�w��宇৐OV��1&��V���i�3��09m	[w>�d˜�n�.r����%�M�����V.S�ڣ����؏ �	|d}B�F8Ǎ�s�:���f;���Qڝ�&͝�K�O���H�)>͘5�U�g����ai���8�[*�Iڼ�����=��F�uZ�y��7z�'Ɋ3��)�r��o"�5I���Hh|���i��o0�i��b�����;lG���tL%t�����"�x�5�RBhK���z�� D��[M�́����b�a�����Dk�R��g�MT�ZX.�f`p�V�ϑ'?������%�hj�'P���f�Ye)p&��M٭�CI[����ҋ�W؛�;%�����a� N4j~&w�M/K?�?�_��_���y�����M�y���K�;mrl��.7dz���\�f��hc	ⷮ�iz�6���wx��O�dM"�m���K�]��p�gx���tڵ��p��&���u��⨡/;��J���{��{�L�o����n�G\:�(�)*�$Bh!�`�@:J��ٻj4'����o�_��Ǚ������5���Li2Nߗ�
�+��w��������x~[�ܼ�����ޖ�y�h��~ٻvQ�3��ht1���C4ۃ�x^l����u��,ÇV5`��7R����V���1��ڼ�r�7q�����N�����X� U-�6���B���f����,Qp����e��|V8���䣢��IV1 ���/��>�t�춾,�T�K7��C,�A�aSY�B<���?p��4�{��r?�u�{V��q�&�gc�~(S�c�K���p@A����`�������z���w���u���5�,�N������������?�+��~���A0����r�\/�W\_w��z�����~����7�����w����n�q�J�F ����(�!�5Hn��;w:X*��l��0��C�n������?38ZYd�oj�:%�2@�vmؚ��sS�0Sfy�](��^��>�W�J�㓞L�I�NM�'��s<g�crs���g�q|�-�x�N\TE,�r�#���n��f��n�	�W��;#�y�0�6DH�,E-S�&9� �d�v�g�<`��?v��9$߳ϱ�V���e�ѹA鳀�������J�_n?Z>��;�:�L���𕵝�Ro��|g�Ϗ�p���tC�#8�����!9 �@
fysIkJ4p��q�ih���1Lfd�:X�k��^����O�l5d{v,� 
��c����6b�k����PQ~���շ��L�3�$�#��GA�� �!�.Y#�8�����M+���T����ELۥi?�8�y6ۉE.��X�.ú913��D�7YZr����I�v2!�Z����>5wH�[�m]��<J�L3�����pǭtp%�%�)�*�i�hdt7|�S�#�a��	y�t2#.2}cw2ͭ}k�w�~K&���@��H��N�h��)�mXo��\U���������!�ͺ�M�Es����I+���Y���y���:�Rh'�}ig�������������8�=���1�j|gSLzG;��
O�Iz*�r�|�#ET'�fE��a��|�_��6=F;�k�o ne�O��S���c�ޭ���.��wo׾BV�4'�t�\F1h�k�Ne��[�l��A�p!e	�V|ƪ��5C�C�����s:��Q^l���1��rL��I^��A�R��k!'p�u�z�Gp΃�t1)��Dъ������]��-�cA�w���m�dMHrH��1�	ͪ�(�i�_�s���$��M=��|������ӧۛ��}w�IO�K��X'c���ui���RC!f��^
����?�Fxd�]������4H&��R�lpw���H$s��kL�.A�O�i�Ϸ�+��[$dJ���y_���̒�š�Q%��N�z�5��9�m��)��Y�XSH,ՀM|��n��X�2��ƫ�y]��n����n|�����&���äI���,Pi�d�%Òa!��u��,-�3��Q A�ߓu��k
��q��`����&Yf7���I�g�'�E����:���^.8�MҚ}��(*� [	�[X���Z�~dK�A�.�4C��\�qEc��lu=gT��imf�\;�� ���fJ$N4�C�g��Ѱ���g{�����p�u�\<1#Ӝs�;�.�TiǾ�U|����d'�Q$���g��<��n*��ʧ~1�7�}��	�'>u���zG��D��a����d���9� ���w���.t�n!d8�z�oΥx&F��"�\�1���D��w]g�9�j��y��46�a�Nr��z��2<2����-�|���E�&P���	�{7_3S?��ŪhS�%�0Q2�y�Nr�T}o�\��s`'�y�+ٓ6#�7��:�:�5��ؓMN*�+�$TW��Jrr�&mi�%{bj���F���A���X�+�������$�K{wۡ�J�`���,�O�������zXn�zS�wO\���{����uGʎD@��p}'�N�&�����4`�V5=$آ݈cO��*�Yc�[X���XB$���&�̉�������W���� o��0ցՌ56���N�J"����6�o��1w�E钀J��?�d�FXJU��ͨ��67�V' �q��w���V̬�%��X��3_��֕�{۩�_^q�{���b�]O�G����`u�����1�t��^x�����c-����c��s�kl�����$�7�c�9�K�H�F_U�R�;ᐨ��:�o�C^��0�A�����N}��p�;Pz��'yf!��>2A��e��۝���+�*�w����ݖ�X����D��[��FQ�`=u
�m�ìW9}����v��I�����w��(�2`ۧ6a	���X��8����R\l�2�� �mlhz����_���������;���W����=�|y����z�^��=�>�䓺U�y\����{�;�=��?ϐ��-��t�20Y^�%*o��UHk@;Γ6	��� #���9lc���:^�/3�FFߒ�:��4!����� �ΖgEuW�ͳ�k�~'+��S��>��)z��k]�_yc�v���der����r��,&�9�7��F��@g<�v��T��r�A�M�~a\s:O�P3�����R�U�,��mŻ-c��6pz��W�Hę�������W7����A't�/
���q� m�O�/�:@�Y���W������rw�#�E�%n�IA>�2q�@{�k�d���x^ñ�%AJ'j�Vj;�z�:�� Iiw�Ｈb�f'Lv��>����z�p��]�ݴK
-�0�k���t�i7$��;�u.2;��v�E=\�7���W6��41��*s�NT$P��O9�	���2�ɸE[S}<�&Gj�y=D�z�v=h�����+g���l�7l�oɗ���#�9�N0�=�ʣ��e�X����;�dz�]Z�ݮwB��v���p����)�5��o�K}�Q����e#�.!���S
���X2B�j�sRq��y�Z:�ڏ~I���g������gQ�5LNJϛ��
�z/�y�5�q�۴V�&YG�9�,E�;���^�<
YNh�����=[��S�]~v{�;oc�=���y/��yyT�	|v�������Kh�C�	A��%IQY�5�%��0ԂEO���:��� �%N�ˠ/�"����]��7�>�I��	<��Yr��/��1sq�f����o)t�j�k���$]XK�q�^.�M�9�v\�Xw�k&gR� ��gL#br���eT�<����^tsOmM��܏�N�x>'����Fk?�,�*��))5t��}�����6C��zU�@N��G���=���@�;Zj�Yݝ�����ZJ��5\�N�-���!>��I?2:ZR������Ӝ�:���S}U����8��Q�=ԓ�h��v�wfKܑ����_���'�9�'	X�*h�3cd��D3�9�7d�}[r�Շ�#�'ل��`���źL�f��4Be:�wzO�_;Ňc�{�5����ؐ �@���u��A�'8�;������F+�A��>I�>�Č��Y��M�j�+0M|	;������H!���9 ?" ���y�ŭ�WX�sڄg[�ׁ�c=�7:��L[N���t�f��M7v��Y�f(2a���q+Y;Ӛe����I�l�]��eO�˱�E;a�g�ֹB�F����AH7�Հ���U>u�u<"��n�e�u�B�<�6s���N�5��.4L��Jck.�A�N�?��dz_���g�Pײ��Z�M�c�S.r�A�m�g|�u/����0�, ���-,0ױ������x3�&.A�rb��Wr��b�q�qk���v�����-*ҫ>c�\��LVhP[{r��*X! �㕟��q�Ql�q�5U�P,�yہ鰆����|�Z��y�����6�VZp=�<:�$��NC&��9���<FS�{1�)m�+��R��+�e4�AwZmS����l��zH�d���Q�`�7�J0�a�2d���.�kX��mv�����5���	gYkm��%,�+�aW,�	g[пg�/N#�<3��Bg_/�q���$��~��Bg���6�ߎM)=k�6�1�Y�S��A��<������c_$ưv�.Rzu�D��a��v��*���$sR�|��x�%�<]�瀅��O�g��R�N��s�gbQ��ʧ�Ǯ���Q5d�۪���:N����������r�����5a^����z����' ���'ӫS��\�����\��wS�hF.���� �ƥ@'��k6�g��{,�f@4k���+��e����ߪG�;�∿]�ȜF{Y��<���:�!�۝��niy���l�Œ%Ck#��a� �؃YHK���걆�(;���]���(�]�V?P'��s@���״��hr�������U XJN;J`~�	�m���8����a�v?+}Y�O,��մ���۹�㰳�r���X�9�0ڎ{ϩܑ�I���Kv� V^��:�΁�w�仏���O�֙���u a�`���<�0�g�[�f�ꈱs�%��I���sxt2���c(�Ȗ]�X#0pr9K{Gv�mca��ri�uޕ"K��f&�8�ֱ�}��Ľj6�_AB���i%��M�?{�2�S֪͏�����	؝��2��¦�@���x����kv��l4������N�7�z��#���_q�;����i�g��ӯ��sqESMtp���]�R�[�����IKz.ў���0ݗ�?�to�IO|���M4E�Zs��Oc�LD�;�lC��O�����~X�:E�V�������!s�%t�7y�P��]��e�=��;v���?�?5��v|�w�B?|��Hs��.�3�p�u�(��z ����c	}���~���|�K��t��{v���2���y9��:i�G-�E�ԏ�#"H���f����I�������f��*�x~��{��8sܚ����$�/Os���JW��l��&�{|}h3�h��<Ƴ�1��\(ͰFݝ�t��R1C�S�@Ъ8�����2�8	n���|�v|�4A�|0�T�!C���#Ɛ��*�o�^��1g�������y}#X^�N��r$�!7��h������x�}�XO��6�iH�b���JK���L6�t�Jc��7��(�|~�imV@�����8D��p؏�j�~#uZq�(W�A0�[\g?I�YN~"O������wXezO�3�����+�|\;_*�P�g�@'an3+��9y�'�g�g���S�)�����%�˗���zfZP`��%������=f��W�I�W�1^ao��i�KXǳ�;�L�$�->@"K�ñ@1��>���``s��V����y�X
�k�	8���M3/2�>�����]'�<G��EE��3�e ��p�3�����q�p,���p����َN�f�/&��C=ǿr���������h[
O,�<K�Kȕ|����s֓��tv6�x�e:��0�� �?'�P�����J>��,�yc���W��&��N����5��B7����.pČ�rW���e��ɾ����:�T�^S$�;&ɨt���9�ϖQ"Hh6J��ꆗ�g;�7�Cי�9�a�u��H�&k��*�D�y�FJ����٦�N�6�E����$���4U��`NU��
��'Ǻ�E����'�;�_wՇOiZ��&�N$�OX�w��"�f�}�H�Oi"Bq�U�OG��BO�{}�F���;��Z�g���Y�0|�]����VFa�1��h�zP_��~&in{�}�1M��ˤ-�4���Ռ��5>H	W�P����:O�P�g}������$[���{��+���y���>�K�z�v��2�>cC�$�X����r�a��f����Z� {�}A�%��l'���?�e��ݏ58?��=���M��@��ms~d�X���eW�[;��x�o��������r�\/�W]_{��￿}����_���/>������Kw��+��;�z����?�U��9.�C.<G���7D�i54�jƠ*� ɐK�ђi�$�,�	E3ềƹCde�)�d�. k����/��,�`k&f=kv�z^�d�U���N�2Gb�lg�P����J��\�n���cϴ��gAXeU�q��	��<�)J��1d{f�d|�R�<� �R���(���a�����U�9�29�D
�𔋴�� ���&@BwY�1r�5��&�Өx�� �q��O8;x���κ +� �����V���O���#ce>�υ�����Α������s7�.��12qV��3(�����o�hΆ:[_Q�#;KC��[����MW���p��u K���;�[�ޝHE�Po�{8RipҊ#������¨�� �i=�UV�n�.F�8Ŕ������.��_���ǒ��9 ���N�����D;1b��z�l�s�֙�$�X����,#:�&�@�ۭ�EZ�6����V��GBN�lV��S-ɇٹ2G�"W7�`�%��N����+F8d&Jd���+���kdw�!���C����z��tD@��R������`�3/d�]fh��.�V�;�pV&�؛h�b���'��ϚP��;�|�L~�9�l��J�p�<�+x���tk'�u�]Y�'=���;�y��:� C+���2�b�ij��+;���h΁w�3�A�4�I�␳N3vm� ��x�j^YƄUn��}.��MkPD-ık/�����,.�2��m-%��Z���4%��ӽ�۝6�=�#+�|`A�|�0�I�t��H�Q�b�P;B��NOJ8�Z��[�h�ߕm�N4s�+y#S�:O�ɟr�/�A}��-���a��Y&�J*�S���2�e�S���C_�m��b��mJ�j��S�pk����45h�ք)"H��c϶Ư[n��ٲ�h�w��nɇ^�m"��g[�)�L��d��}Ʈ��ώ�m���Ki�����;���A�UK���޸V�R�>�?��"�eJ�Yi�(�v�W}�w����`Z$��,S�%Ly(�H�s��0'����`��]����WiZ��u:5�ɘ�ξ�k�������{OB!_�ǹ��)���ӱGӳ���(��� �T�e��&M���� �#���1�s������B�AliJ��4w#�>>գH4=Z7�fl�Al��1�����,�OP�RMfC�9h�rS�L�a�[r;����.P�[�忎�:-�k���y3^��&ǫk�7�Fsٮ��9��h��p�v�fX2�K]+�l��k2鷎y�1�P���a�+�d��K_�?՞1���k�2��5�ô,�p�OD���� ��]럝Ì�5q��aIZ̖C|����6��,�B?VUO��ہ�W~�2G9��y�5j8-�O2��<����d��N�9��Q�AA��A���t�ܑ���{q����0[���٣�8w��:��_6OF�I�^��8A���;�.w,vpu�-�Ԧ%I����y�·�����=�Jkk�:���T�	����\7ϐ�ҤOxb`����-�r<�{�4:`��}�?�|U��3���6Ƴn�c1?$�q��/�[�Ѧ�(?�xW.W�9$�S����U6�*	��̛t�w��u��i��_�!֪~�/�Sdz?���s:���^}��� ����H�1���&��W�i��%�@�c��x���¥�I��<��f����nc&�{? �æf�B㩢&d�clCW}9t�X�)��lXw>���nK���>'ȑ�v��l�ގ�~�Ҿg�Q���l��H�fJ�<�����x��؁��k_߇��]��Ye��Xl��z$,���՞�u��4ӻ]��._wCo��馝���/���?������tz"z�9Ny�^�������N B������O��_�����������o��~{�|�����Z��P�fEC���bM%�@�
�9�	�\&A9U��
��~�LA��<�����ՙ2i�[�D';����g�!a!�;#� J��3W�w���ov0v)b�j9�*F�h ��o0:�7�I	�&�ꎬ���x����o�����ާ]WƳA�������'��>����wl���<��k8R��|�`��9���9�u]�,��8�w�Co����B¼k�$x��
��1��٩��5g?�da��pF���k>X�9����i���S�|�-X8�=�n��# ��҉>�U@�$2�0��+�ݦ���"��p�7�O���!k�ڎ8��B�n�:l|m����B�X�)9�@��#N0�¸1`���K�Gu>��gv�c�[�w�	�W�<���悏s�0��-��D=ʘ)��#�����+��sj���L�g��Z�h�A45aN�6��.�
��e7Z]�s���L�J]������155��U��2�T�gz�n�b��uKp ���)���,���g	�W#}>�@��Y��G]��Ӂg��,O�.�u&��0�>��tvryE�C�}��Y8����'Y��MmL�;9q&>8�/aĹ<'���x8.�2$c"�Ypz$�'�2�>D�#I I$��a�'2��;N"������ϒ���K��e?c��c,l�J�����+�H���b��9�z�/��J���!�%�`8Ƕ6�8���0�^6��I�SZ?<���pn��rI��O�<;d�;�A[#�$�xZH�Ę=����%r�*/9�9a�;J}rE��	g���)��8㙙�����ZdSq�fJ<��s��*�}jt�_���z��,p`C�Ki�<��#�X%��4I[�	�����l��\���c�d��*�6����~M23LTG��&/�bVIr!�f��������b��X��@_+��#�>zb�ɑ����s�VB'Qg����l��M�~��(�S}@��A�p��iI&y�eQ1�E=9�L�mZGĜ��.��~��f��_�8ä7�&`2Ų�M�#�Je��5���tdM�"����u1W�d����s,��p-���2���tpEC��%s�iԧy�X\ov�BrE��Up��l�W������0������-���'��r�,�f�6a��F����i8ɬ�T�}V��::����C%��I���Q�,�J�'�͂�� ����r��'5�?M���lS	�z��Y��[!SM ��atJ���5��+���\Yg�a�����O��n!m�+vd�5NBIJDngR��{1oб�f��a���o� 5v�d
���?g�i��@���|�	�z�`j����lc�(�S��Yq���1q�Oi�F �Sr��w�3�]��;�ڶ��/p`�w�n����{��0�θL�V�+#�&��>R�X��=v����f�t�r:|A�����A_�^�4�d�u��z�l`�.pה��@�v
�s=@�>�/�5B�!�@�wԚd}���_����?�}�����A�Q>�}�Ml�u_��dSF���L�t۰[Rk�~I�+�d�&�!�g��`m^��b?��`w`]�GB��������%�?Kx�1����Ә�`����+�3B�f�;�.��t9��"o�>���������/���n�~|{{���v�2�^����z���O h��~���o���������������]ڟ�H�Χ*J��pw0BY�g(2�,���j����,��5�������$��As�&7Ƴ֛�yO��\LY���1'�:Ɠ}��K���F5���ߟ���7�K�Ϟ���U,�F~[7+}�9��X�2,�� OpJ���n̤�aD<�4�K��F��A?/��,�L	�3h%S�J�d� �0$����4i���מ��>$�������PPfs�0���qv��`�@�0�l��L��l>�g�ޫc~��g���Ƙ���w�}q����������;P ' ��2���]��0�r"A��(���.�빖�m��aa|���ˣ׻�Y68$���j��Fv{�gXE�fO���mۼ�f�˄��BsVM��TaCh�]�pN��G>�uَ���]��:m���ݖ�����l�%7��U5p8���#b*��r��w��r��|,������N����P����dB��������kX��E�M��'Ƚ��Ӿ�3�a������
"�H�dCB���N}�;��r|~/��cJf�.2"H�38�R�>����?�N-�5�#k;�I�
"KM���u�A@��c��;��g���Կ�����o��<��(٬��3� � iܛU�h�6�Y�o�4�B�Sd�-[?��4>�	�A!	�J��7��"����D��������ݡ��u,�P��'><�CH�6ə�S=�k8k��5�"�z>���DU�Κv��;4hÓOs�љ�nI�5�f�mW����a&;C��	6���أ��w�[�M�d�*�;�_{rX�3Oԧv�ε>�%�:��@�ʖ6�]74�إX� �(�9X�����d���:�c~��_�msߦ����y��+v�m~?�U��Tm��:�]�9��2�I�>���۱�y=f�e��˶y�"l<�%����$�zx3�֑D"o��|�Ac�	DH�b1�\�Fs��cB��Y�<��1����iW���p��a�U?�_�sRU�2:5�����zB'}o�8��~�{��k��E~k�}ι����U��U�[4�QcY<G,F�� $�Bb�Z��1`�? s`��d!�C0 a�,�	B�� �~�����Uu_�}�����������>պ5�WVݳ��V~������|i�],PE���f�H�FN:1���8�����ݏ7�;U�Ԏ3����XF|�n��+�ܭ�褌M�7�[K6[$%���Cw)���VNB�G�T�:�U�vi5'���*�����[�5�y��V�s�o芡/$Ɓ��ϭ\9��*�����7���^ q��ې}W謏abM�@�zg�*��ت\Z?㢻^4+�,�7�����s��}T?���-��X��'e��j*�_=T.���zRq�����[���J9��ۆOm-����!]Mj��AC'��4f���%�w�ě�M��;��[��������a���R�Jٵ1�-���u,��^N��I�_\L�46߮�y]0ٻ�`X��n"�p!f4��zC���0�-����(�]d�8�R�Ɍ��͍Ơ>�5����	\�g���}�;9�`\0"�V�j>��l{oI}h�G��������X�=bw駵-����Y�\O���ݖw?��p�/2������O����X�~u�鱋�od�aYф:�����,�X��r=���oW:^�r>Hub��2~��b�	*F�8I�&믶h�G<��L��P�x1���?W�����ۻ�U"�2��j����B�Ĝ�wJ�/�L����W��o����=�:�:����Q�����tI�tI-}� �
��o�ܾ}p�����я~�������gw��:��6CRF^A{hΧ�T��M���QJ�
U�3���f��"P%F�A&Nx�$��KS�:
��t��ɂ�^b��=V�@��b���rl����|��>�h{�ѻWo����W���e�h�w+���W�&q>��\�]"�����p%%�pJ�`	�#�#�Ω�Ǻ[��(/#mń]9(@Z'�zvᣬ�>���.�>e]m�������ה�d�U�P*��O��PN�F��շ�E#��q9*v7�OK3:�R':Qz��v��cy�L<NvmN��BV�V��#XT0�@XOH�	~n���XR��-�J/��@
B���ihw�B�
	ҝ�|L[��ǋ���zt�^��,6�a�H�8�2|�NW���4=�����.��ϝ[�1�9�g{�?�t6��w;�D�&`�Y�9,��Fs-����S/N�,�@�\h(A?��ɲR��C�@�a9�]N��â�\�C�Uy�ؽ�T�Ҥ}��D��Z�qtN1��D:�9NNb�"3�?)F��c��9��ZӔ�@c�Us����m[@���&�2ԝ8�hQy�?�,�[�tS��v%�6R��*ϓ�3� ��"勝��(k����rߨA���G>Ha'�k���x�C2t����L�4K`]���횶1��ln���c�'n��f�Ǫ�fT�9hZ�s;m�ٍ�Ĝ�	o�	%(��1^�	v� NC�#���a�*�����I��^AI�\�d{Ͻ�vB��T.J��������_h��I�B#�Gݮ�@��I�@s�%[���o����U�pQºj�"_Rg4a���K�1�}ݝ��D�E>��,}��Ŗvk;z�mL�p����z��JS��W-�Q��k�.Z-�0�
�L����YHmhlp�w�,�1�m|�]�ݮ�$�,�O��L�H�0NK���}r��,]��It�������GTtz��WDψ���6w��Yڔ�tİ���b_�>h��[�'�Q�}���>t�e+�y��6"�˓�zǳ�������
�_~�j�w���i��S}S��՘|����ON�}^��'���oc�/�Kp�v)Sƙ�XX%�c��L�q�.�2y�v�.�Gݒ��l���-�p�Yu?� ��*�N0� :C&�:�&��؏F hS,��Hq��3��󵍋*+�"3��uxO����N�v����ۺ4L�d1���2�D3�	I�DO�z��H��/̐���)��Ƕ.8����}��7X-���p���x(t��0��E8�&�1A�g����f؟ÿ,��ă~��8)�I\IO]ԅ�@��2-8���B��q5��pF{a��O��b�n���������� ��緛Ct��|��b"�B�b�����e�l���m�R�v�$�( ��Y�V��B����ݱ�Qm�k?Q)�zd$>5Oǭ�eޅ�zQS�^�氿����62.�H$�q,}=�H+��
HO{��7�u��ґ���Az(�?��a�}���8M�@x�P��u�w,tW�ATpC��|D��9��ӈ�Iu��1�/�4�?p�R���&�:��,��R�V����&X�D=w{n������uW�}�0��8��T0���Ҟ*��9�����*�uy��o���ۗWWW��Fx~I�tI���7}@M��'3����z\�~;�]��I��Q���*���[C`A��� ���A�s~�O���N�	8( ���oԉO�nyG������۩-fx��;��h1Ve���dx�N���)��w�x}@������g�����9�� g�c{ԡ�zp"|����H��<��.e�`���c��},�?��X�Ӛ�qo�@0}�:m�+X3�H�8���m��Lx��)��I�?�CĿ�
B����2�:- �N˲���Й
��1n\�N�aD���՘�\�!����g+C\�:��I�����8�}�����$VGQ����-o�Ed�B	�����벀�� �$��-��������C�;'9�a��qE�\@�օcG����?���<ТoR�eX�N��$؁�܅��3	/���w"g��qM�h���?�_�_l�1*z���`��%p���10`��N�¤�W	=�����ft�D��L0���Fi��Af��)a�v��%�JQ�,b�H�e�f$u;����~���7o/|�d2G﫳vS��7�6c�pb�M�����£��_;����Lro9�6��8Ts�׎���U&�P7��������|��Fr;/d�V_ēd1��e�52C ڧu��K�ݼ�ؔ4�H�L�W2)&�ד�V[�!���S�|�:�Z�B����#�h~�	���H��ӌz��^_]�O�5{�8ER�qt���'�����Y&&a|��b~l0��+�JP���>�k	���Glo��t%����P�d���z�O�H%�/��-WmI2�L�ma���^����&�c��7mS^K�,�Ӛ�q.Dg�`C�([���oE�+�0���w}mt���1�
��-�7Xc�cq,�S3��7�C�d�oz�Ջ�� (SV8���fԅ(7Y%8�ߥ��ˑI\�����?qci۲��m�2�C��G�}��:<�:ʩV��đ�q��8��jk�����JV�W������.*���m���)<슰6-.�@8^m��s�e��a;�H'_�w]��q�Or-����Sg��Ə~FI+��^`���7��?V�R�k+r��1�p��x��}� �gWL��!���X�ߞW��l���q�Ot|cl�q�m����U[Z�7�=��w;=��ؼg���)C~n�l��l�[� �N���2�$<����Q�-�ܨ9��tW?��ڞ�m����mc��5�?����.\Xz}(6F��h�ly��z�g"#�^f�{\L����b"A���S�i�~�+�2�ca}&�<˿��zcQ��,3{��x�F�p���\�J^���, �J�q��7�1?�x��v�U�m��4
>S��X"Gƌ�GKM���Յ�o���B�Mb��,������JO�#zEw�����f9�a�c����u�'�[��xC܈>��G�Y*ގ����iQRZ�"�`�IJ��Oi߶���B��� �%mi�D2�^�u�>x����݉���|�����%]�%]R��� ��BJO鋗Ͼ�?����+���?��'���mQ�ѻq�"-�����.V��l0i �c��e�"gà���6ؠ�(h\]�u�I��T?���+�V�������F���Go���G:~��>Xo��O�����`�%-�c����v>��)��~R�9GƂ,e�y<�^�(�ƿm�l�l� ۣ���$�n@����30�Z�i�i�֏��q�PF�+�׸�lxGǍ WY͏2��.�o��dx@�˦�#��2ʝU\V��mq���H;�6�%@Ab�������oϴ��~W&���I[s��0�+~V}bA#�6��ߎ흣�:T2_��ra!�z�H4��͔��1�q%�5{��i�2�i��(�K��{�oq��E?� ���h�ǱleN����S��Ӵf��9H-_�6LW�#�Q��+�Hݲ����e�t캢C�|D���i���ԁ�
��w�⤚t˂�V�T���du(�qj��R���@�Oގ�s�g�f�q�6�ؐl���x`Ny�U#t��fSO�g�M]Yp�e���ү����P���)��|yg#���-�m��-���wh�]��Uv��)��U�v>�6�S��s��n�����&a�����}7� $�.��*�-[Ȥȸ�fP����0Gfk�;�"�~� �w�Qo��2,��6��<j�mHB~ӭ��/�ͨkF�'c#�-���i��9��D�t��Ń�9��_�F��Լ�ྐྵF!�=��]U1lٗ�Ό5��'=i@�&-�7D�awX#@�m.40t����h+o~�ڶ��^�[�	���e��p
�ٶA"��D�\�.l.h�w��H~�(�:�fȪ+;`3��SYt+�x��}�R���xk��U�<��J��`�yQ���x=�)2�;X<ż_�7Ns�u�:d�����h�GZB�^$�t��\�4��e)?Pn��6�O"j�G~2]-�Z�כ�GL�
����8jZR���N������	 )�m<���q1��\ʮ��AH��MD�'7��0z��UW��)r���v�������/;vBN�!��,�D���M��]�`�2Y��r«nh�'�X��Eڀ�ml.��	���?����Ǭ��.�Pk�ge#��i�3���b[�Ő��Y��A���>�̻�׶H[ډKb;��TU�V�`s]�	 �h�z����A�O\(ƒ|O
�}V���.�EB�+M>.f;EG2N���~ǿ\��[��P-��-�Cw飞LP&��nB�{ۥN�P�j'm��y�����!^���A�f�i?�<��u�F�`?�Κ���������:�k�Y���Y���.��:ǌ���a��z�h��Y/�=ҟ���ᗞҷ>~B_>���+J7�zj�ڮ6H���krH$�E`;�Ά���N�El�ǧ^Nk-�Dt],�KU����W�}b�	�R�Z:��Y\���F��++�>�����_=����y�����y�b��GqI�tI��/���������/�������Ͻ{�?<^�C��R��>\]W�,w�-p4*m=>�|� H���;����B8�)�O]����`��R�
�~�0�u�;(j����Y�L��NƳYv�_����▎_����C�ΓO��O�ӫ/�������J�o�hJm�A�[�0��l�a�Z�2 R�42�H��Ge%^��=��1�����}��61� �mU^vG�8Y���y.9l�0�A�@���~^6eH�!</H�ws%�}-��;��~���$�ʳL9�/�q)CPW!�p���$��k�!rĿon��D�S�Z�S_��	1+�:ҏ��q�At��s7EAB����߁��7�aƹ��98*�n�y��:��=��$�Ȟ���Q(�R;.�=�e�ں9��k'���u힓�Ι:�vU��a�ViP�*���j'�j�YF���N�W��g/��?:���yx_�q�S��n�Av禔�(�<�<��^�=�Z�K�w��L_{����F:B��^�>��+8/w9��Iݾ��<+i�lo\R؏cҦ���w��xWۗ{ cJ�1H8n�X��9=��PR��[��<?1�m �u�$Т��j�k���'#��"/���R{;�?C�J���8m1�a^)������ݷ�Χ4����n�hx���a �S��>x����3��Rw~G��27�=�Q��T�2�m��`�����1,�m�^=��o=߲�	�Q>���s<�Gq����Q��+>Aen7�w�(�O-#~/���i�6���1����'A�u��h��= },4�	�*0:5g#K�;�aY��<ΰ�B��� �%��Ǔ�אf}i4�����{!��}�w@C��b����GB+��N�g8l'�[
h�>%x��=�0\H���qH����k_j$[�����3TG�_[l!������G�ۻ~!���.uy�&����-�OUNJ�s�Q��986t�׶%����]@���h�:��`��BO�{c�	�VO���u����O���iX��*oӝ���~2�2�zΛ�����ƅ��0>��T���L����HW�-!SnC��Xt�A�ƉM��ݞ%o�$���c��
9���n�^�Ȳ�[߷������D�]�b�zɨw�,fZ�������#�0by�&·:���@�ou�(�3��Q���&f3b.�O 5��QJ�i~9NN.-WU��_o�^�ї����r������úɱ�|�e��g�E���q�sG�&-�T��?�Q�8�m=6r�}�N	���}�6O�G$qw�Q{�����8�f��|��u*Xtg9�q;��v������������w?���ן�x���ӧOo�.�.i'}� ������������_����ۧ�mMW��iY�nÓR\My�j;�z A�w5P
�rW�xd�&�l^�7���jҕ~���1��YW�W��U)ReQ�-��*?�f�o��7���׷t��}�<��R'�_|�u]���1�zA�f7�,�|�y?X ;�9r����,u|�_���'��͎qRzfu�9+-�Ti�"����C��#��w!۪�zL�??BR�|
h����'�|y�Y�TW{笠O�	@f�R��ߴ����N��:�#�0�SƸkY� ;��^zo� F���%�Y�����վ�iJj�\�����������kұ;q��C��8�����sf��Ǚ椈m��=���S�Xg(��c0�m6�(Q�K�\�=���of����	e4 _�ǋ�{6����o�G2y�;���x�ʘ�q����4L���6�\жGc���}_E}4������+�W�b��1�ϗ"~	~'|�w�m0�e���4^K���b?��(�!�pt-C�޷:Hpv�b0m�'��e��/
g"rb��[����d�SGvƖ�80�����.��à��\d�gc�\���?
�IbzF�[z#�U>>}���b���6�y��{]���A�q�9�2��cюӺ��VU��6����T�w��t��1�}ϦHf�M�M݋�)N󾨍�����q���O�;w21�˗��~�w��ڳ�q۔�g���Qδ��C�<���)���?�Y�mW���GX���>����O�k����L�|)�h��r��ڟHo�?��9}{ډ���s6��,Z��3�R���[�/kc-}�;��:@������F�a���4�/G�^�������%b̝iO�#�iE?�/��v��Gd(;����m�r@����з^�b�x�����/��/��G\���>�ŋ���g���f9mw�k�.`�WV��L�J�\��-�^�Ԗڞ��&��5�G즴�Y�<��6�I�3�/��\�>�}���i%�Uťor[�5�k ʉ:��B_��O�[�����L_={G�O��Z��+��¹��UvE�:��������V7߻�ȘU}S��E�x\�e�TZ�'��L�+�0-���^��ܮYc�������|������o�'������o��?�OOo�9�K~�%]�%]RK��	 ?���_>{����ן���[��=�tH��zr�x�;��ʪ0T�lp����B�`��a�@�jZ��d�2ޓ�A(�д�q��,�V��'W�5>B��z\   `�ƴO����(����ڝ|q]�;f:>{K��w�����'��g���/��e[���e�@=�8��m��kF'����as<-X���@���*�5W_�U��pvg�9�#�_F`n�����x��`u^v�Ú�΂{���Q](�6x����g{�5�F��!rn[�50���1�r|�2)3:R�I�L�'zǂ�1�4*P�y�9V%��0���h��P4%S9b�u�l���K�PR1�����׽�@���'�&ߎ��.�z�.lwD�q`=q ��p}J8����?�~��>��0ߗ^����}��H���@�8�:n���.���_<]v��\������a[�<F4E�Eυf��������8**�-[���V/G�G����q/Xj���h������;�1//ߘ�v껺+x�LV�S�����e�Wp{�A���x%F�%_��ڰ�86��$�����ԫO�c/�{���(G{2�ͱ���j��1f��� �(�w�^�vl���x� }��U�.�\��|�z^{=���/˯� 0���iۗZ��8��O�C��F�XD~?�?q�>M�L�ɸ��1����}�a���9:�<���!F��i�߰��W�b?FN���'z/��a��>�vB���_�ۋ����_O_�Q�g�{��S����7�ձ��c�������}|�g��p�L�����F�G1�b�����{8&�e/Ec�.�dsVfLc-]m����G����I�(����H$X��1ҩ�\p�j��ߙL��$RloH�����Y˩��� �9ޖ��̆E4 ���>.�����4��v������i䙭w66�~��c�/��Y�Ř���c/?ڏ��2��1q]��	�T�Q�UDmN�WY8L�x�}�'���,u��/��p����K��ԁ��_�O'h�H�]�ؾ���ɞj彷����n]˲�g�Pе��d ���S�N�g�]��?��>�ߪs�/�����7�]�~`1�jk.���2'�t�T.�%����c���u��z5�8����I��L�@Ȇͪ��B]H@!?q�Jӌl�A�������R�ws<,�n?ؖWO���Ǉ�M� ��K���_�oz@Ui�8�w�zu\��꺮�.��++���$F��WR�H�3j��#�8��� @q��B]�_�i����oݪ��n<Ԁ��)�w �q�p}������E|uA�rb	�5#SHC���z@���8����\���;���G������O���_=����Xj86���*E��v��-x�ٴ�#�}�4/��E�r�;$����ߥu�`�s������ʢ���=�Xp�;��A�сM�?\U�z���/� �9Z����mZ��V��i=r�8��9v 2��A� ��N���
|�r�q�H����Q��0X�5Hd�d���v������o��a���qfƄ6�c����,�2�-h&�(F��>�~�E[��l\�ꈂ���\�/
�� ��Y����I$u����YwIx��=z|�Y�Li���4剝��ӱ�~��f˰����I>��E�Ae��ݒJ��{���*�8����`�� �MҶu�K)�.R�wc�ɗ(��xO�^`������0���	JK��1��9�MbD:!j{���t�SL����q�L���q��ǟN��nC�]�3c��5�*L(���S��"0�'��׻��Ѥ��ߕ�}P���Wo��I_���*�$XA��.�^�B�XJ�X[�+Cq~�;�.�+>�b���gŊ��\���e�I~��X��}}�uj�D��3�+��U��i�؍��`%?v����]�h�e1��x1[L�Ǆ���Ի?���`p_�4��ta�;�x�1^�f���I���-��W��]�c�n�� ��Z���4� ���D��w�\l��j�v&����.����r5�3{�v����N��/cf}�����h�v�����a-_���k��{?�_�؊h��<ئ��G���1�(�sF��/�]�G~T,��nF<�m���x���7.4�x�H��]��yթi�cy���"����s���g�!�q������e�!麴�[�`T�ȡ�Zi:H1�bK�q�;S݊2jۛ�v)��&v�q3
�]��b?#bs�?.��#�\�.���*�`^�u.��j�/�ҭ�K���ȗ�Xg��u�ݸ����F����c^�^�":ݏ;/�6&'x�&U��c�F��Y0�sD#{�9r�IO�Xv�K����u��3��q�t
L��g����oK���F.��W&�w$�ND��6({�c��X���3��>����t��t��c�}aM��̝�uP�6-�g]`@m��}�4�&3ϓ,�`��r�c����9�.>R�\kWIpf]	P|���r���*MK�����[��yU���,�0X����8 ]�P[q�0��v��ay�ѷ���x ї�l��%]�%]�,}� �g�}��������w��W�u[��/:�'-�ճ^80W����)���A� O�.�5[��o c��}^����=߲�e�,�[�7��W, �$��X5�b0�6QR�!�b ^-{�����U���S�����}��������9�x���q76FuaA�E03ߝ'�#r�{���2yW����Q�Ԩg�t���"gNh�J�me�����NNt<ƄN�Xoh����>:���
�v�]�[��7�&t��.a۽��N
�]0��u�{�s+H���9	��`�}w~��p�m�Ą�����m��5OQ���(b��w)[+Y�&
x�l���dwĎΌoK�ܗ�����A��>���ɎY��Jc`"Mޱe��������~*�gt����V�0�U$^�G.��e�G��P���r���16��OHx>F��.��q�ù�<?��?��VG�zL�,H��Ʋ<��>�~�q?.�B�@}Bi�v�y��?91�;���l֗^fg�D|��a~�KD���A��#�˗��ni�63�@Zf�閾�Ӝ�=�
��ѿ� ��ݬ���mϖ�0���G��.�8a���l�����'�'r�-��;���,�[y�I#3�z-���V��y��/<�(ȶ���7~f�2��˶4+ְ�4���8��"�AM/ٝ���쌯�0�?:^e�.�8�ЧeE�� 1Yd�}^g��H�p̞�Դ�w+}y8��g��gy(��*�'u`�#�F6�>n���s�#z/�K������Ggvx��Q��M�W���]�/7~�H�=la���B��|��"��/�6$�b���Ot����o����Et݇��2�"����/�D=�y��[��#zf��x��Kc�i�/}9���v�'/�V���e[���B����ہH/����:mQ]^�{���{� �QHB�0ӅZ��7[��b��,}c;"��>=a͍0��C
�Z�㉙����^k�m�Ɗ7�/R���}ߗ�]��?���C�cD������g�GzʏO+��j��m*��}h/s���iT��������9���1��>�r��푾�������җ���c>��S[nʤ��2���b��o��e�ܦ`�" iO�q��Z?�w���z���O�pb������B��E	Dmi�϶p��q=��ex���St��R���Q}g�������@o^�[��Ys=N�����.��L�o|�����������'^���ً�����C>,9�eW��cW߽@oD����$�v*C`�3��b�Mvt����0�
䲮�*Jyi����5Wmť:uޱ��f��?W��%�Ud5���OϾ��姯黏�>{�	����޾|]~=՟��\v0�d�\�wH���ή, ��<CٵT� �-�Oq@�]��l�j��FZ0���@����3G˃E\����F�ʊJ�Q��y�|��l�-i�O�
�:��\��f��|ȓs���2�	�o��s.a�\�¿��H�|���8I������7��<�g�%X5<q�f�جLy>K�Ϩ�Y�C>��=���!*�-���}�6DA�s���E2#�����&u#g�Dܱ�t{:}�Q��ڧ/b��,�ۑ>��,��u�oK�Vߞsr�i�މ�.�L�hP�Vs����y_��6)қ������S�ᩧ�O�l�/Gb�͊�y��t\�{�?�F~�i�� aT�}Ҟ�lVDCDg�i����~�[<�K��>��z=nR�'�Ͽۣk�� ,Ĭ#vO�-�ϴ.�{�����l� �����bz��f��=�*�O�؅_���݌�Y�=�숌aM���v����=��8_��h6�"ڴ�s��x��]�m�}�Q���Q9��s'��G�{~G��\�������d��C�B��|Q�F8X~�ۋQ�h��#�@�z�9㵔}����-���^�ʋ�=.sl�^�g�>��׃�"ٙ�ȟ����9�6k?��Y�Y{���÷�b�Cq=��sl;�����L��^_J}SRIxe���u��c�6�4��Ɣ>ϛ�c����b�NQ�'��������M`����$�^����x�����ئ2'�7,�,ދƿ�SOc�n��'σ<D�D�źUNm��/��"�����o�3��ԗ-�>QZ���g�c*�k���i���A;2b�y�Z�3�[������kE�w_��_��g��_����>zDۃ��r�q�2�d_���I���	J�!��c�9#��yP���,�r_м�1i�{ ���SyR�״5:�~R��	�{%2��^�\��n8KZ������pX�
˚���$��i�K��?{������Wۻ�As��%]�%]�M�� ���ۿ��?����O^���?��і�dy�v2)�`@^��L�)G��1�6ȦI��#7�`�r7��� �J���s�pGM�-� jk���z��RƣMu�"A{��ۘ`�cC�ޥj��SI_���#���_���>���ѻ�oO�z ��;�&��/VD{+�t�=����t .��� h�Pm���- u/83:������{t�c@;���7�/�{��z�6���dC��4Dc��/b�+
���ݟ6x���k�����AqT|��6�p�김�^�(r��s�m�M�W�~���:�H7M���G$�3����'����X�/g�=z�|�s<�����<�m������(h��?��(�Tۘ؞����>�vG�9���v����}9��(Em��������ȸ=h��G�f�|ڢgQ?��è�(`r��������%��lh�N�Q{%�Ĉ�Ģ�~l���<7�-�Pl7���O�o�w��Q�ky�eD�����lO��6��Jm~�K�l�ۙ1>���w�Nv>��W�x���t����	AW���\��Z������..��6F�Z�����[lu��P�E��^/�黟�W��O2�Q�E,�+L�4J�,�c@��������|I���6':¿$�[o��svw��`䉧��q��گ����Œ�n�Y>l��s� �7��=�CT�wE�z�1�#_יִ�۱���sm�h���Y�s��t�����<>]�<�>����`>֥ퟟ0�G�d1�/�G�;�9{��w�ͰO�sfm�����_<m�a��H�St���B�UVՏG�%����t?ӎng�y�5H��WCҽ��};��t�����13O~�YNzU�`mP����,̬�������c���F���F���\�:�#PF:{J�B�ң4�u�;"�����}}c�L��C6�	Q���S�[=�(i�B[��o�.��H�|���C�+'>������iF�H����2s/i�����]헶Do�~M�'�������Dw�;���J7e�����q��F�$s��ʷ�y��;�ſ��§6��W�w�v��ʌ����Փ5����"��y����=2d� _�y��+o*-�b��U[V���6�Sʽ�'�Gǿ����o���������7T�K��K�I��������W����_�������~<�e��J��;4c�X�e�O���E6HŊ��ϟ��~_M�jL������-�R&�]wuh�L�L���^�j�l��R���)��O��LO��/`�]���w�<_闞~�l7���#z��-5��0���k�O�{fzKЍ �w��������x8��旺�	����	ƾ�U��.���кBOA�_�;w���'�y�Y�3xS��`�:o���cFzI"��2�}� �X6GH����=�����=RZ�<������'�{�ev]��:J>8�=}�k�(�,��-���Ć%/;=M�G{�>w]0i.8���8�� ���sG��Hg�w��xe����i�Y�c���M��w�j����������Ϲ@�w����n� ���so��hC�������E}?{��}F��!�e���:��O�^�f}�w�Fz��si&={v`6Q�<O��2�'��f�t$j���W��q�X����qL��F����n�/�me����6��_K���V�.�W�"?ٞۂ �0[v�ԗ�u��A��ݽq1痵����1�ъ@d�g�q�~F�`�(���ƫ$�CF�G�(�+���m�}Ww����r�����KMd��$�����س%���<����~��x�4�#�t:��+a9Q�����w���g��v[���<�OԖȦާ��~����}ʞ��ǒ����ʌ|��5�/���fO�X���`}����E')�Ï��0�σ9�����G��$�p׹�0�σ���F$K�g���6�E�.K����'�xژ��}%�����G���򸇻�.���E���;J���+-KmmJ��I>�̱�[�R6�0���/璕���4�&��ŉ�iii�~Wr���x��"���H���"�����|(��F�O���1�k����i���5�`��86<���O���!<�No�#���=��1�ǰ�Vx��w����e��-�g#��PI�Dƾ�؞���`\\+���΋$z��Z����M?~�9�K�h�䆖�T7��,����?�S�j��>N��Uc��-���e�f�|`H�<��d�����\/M��X�8^[y��r5�{y\���k���R��{^�P��͉���p�Ǜۿ���կN�?�N��G|�. .�.�L�F ��Io�T��mtx��ӧ��o��\�]9�H��E]F�8�ՓD�bP���v��vދ�݀r�
�0@��nQة�f�;�j���\��VV{mǕW���v�M�����D1~oOF��t�*�w�n�W���~N���n��21H�v�L��[`n��"���+-�<�{G�M��~�G��K����~�����I�>��$�uB����u�+�e#_6�W{����{pR��3���.&���3�$�~/����`�[�P���F���N�w�nvi�,�ث���y�K�#�wi�'i�3:�V�!PE ��!4Z�}#��ٛ�{x��u[>�\�]*�0�b�X����GW��n��$+��*�1��۪����H�m�`�}_��؏h���,�'	}�ǿ��i��fܑ��v�|��Gv�Eu��%*��;��l��(�����t���>����"���qq�,x��#>���^?���	��Kd����$_w$?Q�D�F�k�6�7 oH�{�c��=}�y,��@׌_��_Dc�O��z�6�Gw�����{���l�|?`���i�9�O�Y�}��NA�d�K������F���v�z�$x֋uҠ#8�b}�ZB���y$S�mj��kM�	����1�g�a�1ʤ`���`�g3���2\���x��~B��5��3�o��1��Sd���:�w��Yfm�k�Lg���o���h�����+�#������}�l�F<����1�����j�D4�~̅��f��n��|�(��O{ܵ.,�6;d����:gxl��<1�E
�1�}\�n�Id�↙��0�o�>�_p�WG��o�&?nS��Tˌ��}|%K��#�t��]̌��mʨ��b�饨=3�3�a��+i�/S4.Q�H\b�����K}o��-c~���[m��1`�ym�xSZ�J������_���ӉN�}�ql��m&�ui���9��?n&���(�-P?�'��R��T�9F�!�����ǓP"�D�#�ÿ!9��@��q��-2���zs>�lj;D���A��o-��V���O���n�g�|J_�>�7Ϗ�<==����p๑T�E�ƥl�˲{?����E���c����R�y�e2�Q����`icB���O��g�k2�����xm���G�Z����l.-3W���-�����ӏ�>?�~~�Sv��A��tI�tIa�E� PR��v����}�]��n�K�Ц�rCP�Vou��z��L6S���y�	v�Fa�:`����ˊ�"�!Z:�bx�X,�4�����/���l
�Ũml�|*���z����-=xsE�{�-�z���_�����t��Ik-��]IM��h� �qU�����pD'�@y���
WF`��(�
- 0�e�7s�U���#'~�����Z��+=y��Ԓ,�Cۈ�փ��^�N6��ԥ�:J�]ۄud�48��=�Y���4:]����5KZ��r�8��+v�Ə�c�#��Ȓ	�9�<:y�Yt�,��P��A��i]�m�C���o<Р������{�I�c^��U�Cg>iE�2���6�ɳmcL�~��i��L���Z��a�Gz<��n<ߦ��Ic�9�v�O�f�"���._�1q�ͳ1bo��^���Ɓl_�>b%K;��/�8�<��܈����ZKD����r�0���ʚ뽱�������1�K��s�(��?�g֟ѻ��|�~�d��xt%��'�����3VF���.���8FM����0VHDƾN��S.�>��3����$,���n�F�*��*�'N(O3��q� �'HKf�y�+�c{F��~j���i�(0�L��d���8&��*�:���ý�M�Du�<Q�ܷAqSޥ�]��3��{����6�<�<�>Q�Mf�h�9�5�u4&���>_�؈�Jd�|�{X0�7�|�3y��g�"�JQ�>�o���>�8�ǜOc�~���w{��b}���1�˳��1�v�z��<��B��E�3]6���8�7k���o�,_��6��٘�^�d7<���(W&�l}hO�t¸��]3?j6VQwҮ��~��DmW|_j�S�2��}�2k�B�E�a�[ZG̵��2cޱM�����k��񀱅�*��.?�*�,�p���J�=����ݤfqaɢW1��3��LlO��޶عy�M��a��������/������߂s����S�� ��>�g��~M7��>���^����;Z�^����~�^�Rv���M�3�9�����b2�M�4�Rjy�;��&W~w�k�7���9%<���]��������o��e3գ�O�������7Y����K��K�M����h���z����O����?|�|�}���R:\��ZU��1�'�'�Do�=x�*�c�F'�d�c�=/e��k��9=����`�Ro*������������a]�����l裫'���������7�wtR�J�����#1�{��>UYЁ���/��Y`��	��om���Ohj���.R����j4��K{ԓ�]��jL�e��L%;.¶&%�Ev��h�p۽?.�_e�K��}�/8�4K#��A��36s�����h)��X���đ��`��8 ��&�e��X��x�rƝ4�Z�ޭw���LOi e?X;��Bi��3�Y�2�a�:�cG�}�}�zܙ�c5��>�W�(oU��'LY����4f��P�����Bod��I�� �X�����T��1�zc>P�ǧ�D��$�,`}�ъ�a�3��;���d?����E��8��DxF����}d.j�}�bѨ'=��n�Y_���у����������=��<�q$�X�w�?��W�����@���=��m[������Y?u���ido]:���lˉ�5�.�gc߯:NƤ+�'�7�"��7^gi���A�Q��oֶ���گ����2Y�7$��bz2e��À�͸�6j�}h������Y����}Q�я�������4�h�Ft����k�vI��^�Q�,��l�Q3�1ӡX'O>�\����N��i��]�ya�^����+k�w�t댇3"9�k����<���h��;�[�._T./��M1�w���`�/y�cO�����c�c�d�+ſ��Q/J��>�����{�_@�*)�X&��δ�vJ���lo��+��1�1W����O)_N��#��2QوE�/>�i\�4�?+����Fi�N��@^NrF9�8'���x}�ʘ?Q��4ڴX��;���q�1+�nR��D�t�������Q�}bSƐ�s<�b���l��J-�J/�T�X���w���x��^ߌn�t�c �;�k�x����L8�;E�U�h�:V�>ٰ��x����e��,%O�6��s9e��{����n�|I���o@:�۷wt����:�W�rR��Bw�H����X�&���e1 %-(0FZi�}����v���`��
x�Q�t%�U�_<v��R��c��g]]6p69>˕1�ί�����w��_�g<I77��zwtI�tI����� �V;�zu|�_����~�������r"���蚚��;���F�S����C}9��DY����5[�-j�R6u�Zq�d�����'�ٍ��sk�H��-�p�P.߯)7ZOF���J��_�ջ=�7��ѓ�]�&z���}�O
hǕf�ش����7�t�;���i��8La�آ�9� �p᩿���#m��/΂��x�b��2r�
2����\$六���7��V4�2wG j�ؔ��}��Gc ��ra�|yl��ޤ1�4.�`��zm�U�3�-mB���dM�'�M-@xk��{��:i2�409�;�./�+]qQ��Yy�>��8u]��āX�SCO��ٝhۓ.�;����N]ė�i��m�K�����:�4.�Q]���;{I
�!���5�'�1L��f�E_ҏ2vEm��U��N���E����]uV;��;j�{A�Y`K����9"Z�} ��|�4�/�>{/:�>�HWyڣ;�-]5�}�8h����Ó J���� �s�-X���(p��̭���H�vy"���
D���Q�E��36���<C�7ګ�N�K2��'���
�����du�,INm��^��<Ҽ�2U�h`$�q1�gu��[���1�XO���J#�b��L��NR���L���]2�/�z���JGU3uhw@��'>��t�v*R�|�L�[�v_�z:���c��V��QZl��	������r(zQ&�P��qa����`�&G��f�rI�5E=��yL����k���H&��t�<��\y#����v��]�"�X��>wT��i�� �M�-�s�
��{z>I���v��ܱ[��Q��M �t'�_�z1�,��$��5���:�يa���=hЗl�F�'c�����^����bm�b�|W��tAl��W�ÿ��#³�O�ݿ�ydb�]1�d7�t�eu{e�nF���.�ya���4���������#�����w�dy"�	������S�7�h��J��=�F�^���Zq�[E����;��N�>�#�a����#�[m���L�Ȥ�c�#j�X����w������_���]��N��P��.�/�a��큄�̽܄��rm[6ڠ'��پ�w�GC?,�UְeW$|[�vC�ҷ%��r���E��;�1�Cp>�����F�U����/�VЍe!��Y�m���\��)=�+�A�CaP�1.������	}]|'�Y(��e[Ǉ�i�o��*s�U��W�u���=x|M���m��w��N��z��Ghyp�����	7�����X��?�8*�7����46 �"��y��95�ׅ.u����zq��97�(�A�3ʰ��ķE�W��Jw�ۇ���>�������_��?޶���<yr{�q�K��K��I��, ��?�{?��o��p��x<><)����5ez�/,e���[Z�*p����DC`�9��
9�P*��p3�� s��r��:Q7\.��ʒUg�'��s���3��ٿp�]��}E���[3=:<��n>��(���>ټb�^�xEo��<��ڂ��;���;�fI�C����:߹Ԍ��x�W���l;%�U#����=3'����"����&�P���s�Q���k�&@���;o䝡ѱ�T�[�;;�ԏGg��i�j	9��z{��bޕ��{l����3�f�m�.��,�o�+������q0��:$����F�D.쐷��2�����I��ԶE���it�D>���D�Up�o��V� t�+�twZ���pa� {��>�N�\�"=j����%���Hi�Y�I��%7�����TX�\l:��7���u-�y�ϧFl����:K�>:s�q^U�)P%h��s�*K:��0�K�lc_Z w����$�F�h ��1'C�c�S���Ă��ġr��}�0)�6y@On�]f�Q�Q*�'�[�y?����;2��YU���v�����m0���EqW�d[��ү��A�j���ȞQ�C�I�/S>#q�w����'�Ѷo�o�"Ɛrf-c�����}�����@�V���;�B��<5~I0D��c����h�@��{D����6=m��'~y�6������ő��l�Zel�$�͖��|�ӌ��<Γ���_��o�U��6�J�SN+hy����3��Y}��gڠ��[I%��u�"qk��;,��/�Ks/� dc�}��C _H��)o�9�x蟕��b"��x�.�1�Ԝ������]�a�k/3���������z�C��mӱ�:	�}�6oq�Hع�;o�o=���@�5M��i�Oi2��Zj|��,�&��y��n����֬�Lc�:L�n��&x�2�6�7�X���-��IQo�m���/g��b+�s_��?�7�k���;	.J�r�!��nA�<Kr �BB�;\5�~��Ꮵ���>�d�ʳ`{o8_�9ʁO�.���V?&��*~\	�qd��θ�v��8��e�b6��H��b\��1�c�W�����5MZRÝY��������+5�	=��g#��Z٩<��J;�Q#~X`�;�v��Ef���bJ�B�mf�$:_��R�8@m��FgE5���F��Ӂy��Կ�Ld~��25�4�'�SS����EPNo1Ț�a����d]o�W>�����+�fW���k���E�����-��������I�u"�rx�els�"������5�0b .����O�k�m��e����5J˻DO�#��n���kzs�����P^3O8�p������Տ���'�\$�ԕ�˔,OH�_��҅���;U�7��C��C��`q@)�����������^������FW�^9}w�����͛�?�����|����/��G�_�%]�%]�N�� �������뷏n���ՖxTj;��e�t�!;l�3����48*� 4�0NzT�)@��4vv��KG� ��J)˂��s�l'��(*+oO��pwR�W�����}���r��W'��������՛SSZ;k�%��w\��Fg)rN�w���
v�{Z����^�g�#�|
r��}��I߷�l,K��t�n�#�����Q>��4��89~MV0*P�ݡ��'\^W�#Ͷ���}.`I�6��{�Х��!|� �8�:��c���t܁�8���vrkl�u�b>ā��t�5Pd8斀��$���}��σ8�f��a��\�$��ݩO�^N�y��A��.��w� �,����Z���P�G�����A�r�k���Lz����Y�s�U�^�k���]bu,�=���=/�1䇖o�0{���2�Q�J?X�e��.MSϛ��%_��$�6�	��Ni$^FQ)�?���~�;�FA!mH7� ���K�DJ��V�1D&�0�E6a.�ʮ��R�]��#�g�B��ei�3mbt�2��������2�o����tqi�TI���~?�	��p�6
v��Iy]ǐ˸������Q��ٝ�oM2��*ʢ�q���t���£�c hn#���B�G��+Y$���b{ZYd�_���LN��#��۪1�=`8Y�~K�{�:9m�b��!(K����}ƅ�Po��g)>��n
�r�����)�C���i��3<IE���:�Tמ�){&G�OTG�8#=$:J��g<Y3ʵ�m��"���g���c�镜��Ģ+�I�)���~��m<Bm3�z�@�f��n?��~y.�0�#�o<���Nr����?&���~�2���+\D���Λ��/W��M&1��yBK��}=(�t9��ͳ�2��٤����N�a�c)����[�����6�k�����ψ����]3R�K'�=,���g�C
���1;y�:%�}E9�Qƫ��_��`}�0n'K�i!zm�Ŕv��@���x��ܷ��oGy���6�F�����;���WJ_,��1��N�e&�#�G��=�Kukn��u�����B���}�0o��|�]���4�ޅ|�Vۢt�z�xT�M:Ш��6mb���kʝ�[�1�H[�ᐄV�3�4^�����������z�{���Z���g�GΧ��b�-�S�F�Kh���XD\�j��U�.�cv�I�N;�O�L|�b�$y��_��s��[���Ձ�n˕��˼Ɂ���O|]pݡ΃,ikcN1��v�,���ί�����i����9-���,�>,�-�-�֫+Թx��x�lr�c���%�c1����C�'~����<�7�ן���=<��)��s�^�%]ҟ���/ ��O�W՝,˲�&eW�FwX�-��0�W�1����S8,����f|R�ȈE&rj9�,���� R`T�@��{�7�'X���&o˩n�x�Ѓ�=ܮ��d���S����ћ�|�5Ֆ��vs��N���qTP�:F@+��`u#e�?�A��3�	x����l�z�������_{�):�c�����ލ��� Q��}&w�w�l��E��]�6��ʄ�߱cˋS��2>�讫fxNCc�c?q#�����(�X4���G�m{�C"e�j�?�.��|Za���W��UAB���Q�1�MFH8u�rE��%���O\����Q���XI�N��A{�74��0?�q�LFۊv�o�}V�fE��=K��e�=���Y>�.>�&�vY�� ��A,#�@��| Ԗm۶�<�N�TH��!�8����Ʃb

�
��,}�{���Z"����s�1p�zpO�|n�l��"@j: �����Ik�]��x-�$˂P�i�5'��I�B��6J���4Ч�,�ˠ��]��=D���Ⱘ�; �{�ܮ �A�o���|w�|k��P>�)�i��t؀6�k��~��7�"Զ�|b/�j���gQ���x�;�l�y�}�/����:W�i���cC�h����uք'L5o�Y��S��%�R�؇z�gV�Tٕ _���j! �����[�/�����8���48�/�c�oǲ
}h�����d�+�K�}�c���\ur;�	0�]���E�VάN���n�M���E���ۢ�}��$G�OIt��u��n�;��s�o���yh�������v�C��,]�7Q���U[	�&�n�.k�}�8�m�(;Q�c��v�d�.�'W�S���&��l��V&�EdjR�d��c}�xzi�ɵ��?ɂ�L|��h�e����W�9�cǦb�h1S{�pQ��n�u��7�9Nȃsc���.*�	�B>b���L ��6v,�(t���M~W�l�<�$"<�O�\@�ƙ��L�-q�cL�UQN\�v������KwULR����_� ����f0ɯ�a-�1����Ko7���1�w#�c�x������Q�ڲ,$�r��ʻ#��/]��j�A�ɀ����5�f��Fc�3�������]�W���Y$MG��gt�PC�1�ױ����1�񆧭-��8Nƶy���?�7䯭����@���+c���/'"�0���}���tsw�'���S�c��9�	 ��XZ< �)A�Ji��:��O��m���}ѿے����\�qM��S�Ա,٘��N��������`����qV>�#�kzw��~���w~��s���.�.	�7� ह��~���ݷo�����o^�㚏ԃ>E������� U�Z~��8��,�a�Ftd�4�ow��J�T5;��C#��h�ؠ-v���KA�
�`Xꒂ�\rp}���.�u���<�u-TO�k s�����1��:vz��G�x,�5h�5��[G�1P1,$q��_��"��'ϒ��V��u�[A��&Vq7K����5/Т����`�r�u�ؖj�QA��c(�V'TwzD���k� ��U��ϟ�ыНt2.�?�oʋ}^�Kv��n?�Q=��y|��η���S���������ո�q��d���F�ʊ~��1���ڱi��i������
'�2��I)~��~?m�/�]x;�٘��; �{��2�����*�(����tt�)I�pfW|`�j�ˌj�=&����Q~h;�@ڢ����Wy�X����){g�w�-Z��-*�㘱���&���n/kk�@5�i��ׇ�]mQ�,U��1���z�}O�`��A�]8�t��!T�8�ʆ��������Ϫ��ʒ�X=������wd�h�\?�M��(mC�;�Wl+�.8�vAh���켁�!��'R~���;,��vL>h�L��B;�Ǡ����=V�':���r85������D���$�U�0�	�<ް�O��^ϖw�^ɤW�lَ�(�~�q������y��$��q��[���s}x^��4��[i[o��\��p4�d20�Y;3�=b�=�� ۣ�}p�Y��_]}�$2�O^�4j6�I(�Dc��g� ��S���Gx"�,}L��ҟ+�mqGoK��\�<؞�_���βW�t�c=Ʒ#����Ca_��V�ӟ%�'~-	��C"����[��d?{�F���:+9������N���m},d1�Kw���>O�ߥ������I�����w�v�\����x.����h8^Y{j�!
tX����3N�,����ز���ľ��|&��G-o�ʾ=UǢ�.X�#3��im����wm�H�r\�7N-f:D�.��هlt�UF�-�Ʉ��[����scH�6 �S-_zQ�VĠ�c�jC`�r2�~���5�D�K&Ն)
����m��o:y�6��"���uex�m���}���x��G��by���?��n/��Ȼa���xP�
��p������-��vYH&��X���vBi=oq���Q�Eގt��>^��<���J[�:�R�/��S�cO��T���֖T�e���j�*r�G�z�	�n�'j���i����,��"�znGDU���n�dIW���q�փ_^��Ƿ�o>y}}}���kM����tI����� N:��G���~���?��Ϗ/pxR�fK�;"��d�bIj�}�X�P�`[�0���Y�DyK�-'X=�����K)��K=	&$��VP6直*nq~jF�ݥˀ|��C����')�Ou�e�[�g�[4A�YC~� I@T���g�	�KrW<��x42�PŨΎkN� �����&/)�n$���ۉ�j'	��jsy�쮮�}�NǠ^�3�|�AΞc�KkN��GD�@L<�^/�;��w"xlw�g�t��?3ַ.SB���r �]�<��\����s�{I4�3�I�����Wl����sm5��P�Rд� 2�� _�]��w)��u�t�2�Q�Ǐ=�]V��t5{G�C\�.�����5#}юzMv��ȍ��HG
�~b��������՚a9�o���;OA�|�Yk)���A�p"�m�'�A�2�q��P��b,�������#o��P�2mP )��@ �]���yڜ�h�"A��-<�<D�$:���:_���x��/䕽���z�OdJ�l�����5P<	�4r�؜n��&�񻞬�-K����8�#f�j�N1V�v�b0"rz��S^2]�>X=�2��Z����{�0�3���s� kKr�6�W����L+��g֦[Y���S�K����4}��7jǃ�E�ۯ��T'��&��ocQ`7u��
O�q+�o������_ұ����t�X]�K�v�@6}��@�t��h�0܋���ZDgw�����p4�����KPǭ�	яr� �xr�ʙ�y	�Ei�m�>�rel��i�Z}�|�%9]�\~�.��-f281����_b^�g
`Rz{���x�?Z�
�&-�ӎ:Em'����k�''�/���<hݩamrz	��zW����Q�B�>b_.o�@ڶ�mB=��=�>h��o8^um�:��{=&��ض���/W�kM��hs����`�x��w�K��l���8���l��W�<�!Ť1&�v�1�g��hY�g˙���s�yx�\�cB]���Ɔ��',���l���?���p��,6���DO,GD>���8����E��;���3�|h����������N���� "���f]4B��S�d6"�ϖ�����?t9��� L��*���c�<�>�2i1��ɍ��N��+G1�^n��� +߳�6��ͱ4�7�K�H���U���V���8���*XC��y�|_!)��h�����Wx��~�S�׍y|~�['�E�1.�߉�ݯ'=��R�G�	K�5<��@ZOSҍ����1��'a���&eAJc�螒s�S���e���F��M��欌^W�C)�X�ʹ�G�ⷔw��1�Z�:��Z��޼|�o�ο���?|u<����wxI�tI&�/� Z��ǯ�_��?��?����?�;�Ft��TwL����%��$0��j46:�3A��V%�^�ņ/4��.�����d��W�.�=�sSD�;��ySvZ_���m����Nvs���l�$p�����΂v�|�g�X`���'�NN ��,�3[������s�G�6�eAiP�|H�)� @ۦ��3�3�zg�F�A��y�{|.w��>U:}?������()�������?�ͱ�L��Y�  ��IDAT�-ڇ0|���$U'j�h�<�?���5��cd�'ti������F���\����~��U$��Z�f���3�J�|�"ғl_������L�h0̷c�!�Z�I%rr& }��d̂m�$���;��7��{�ymJ^J����z�-;� �.t��Ǒu�a����ef�W!�����9�.~G���-�N��Լ�J��eI6��:��'�ډ]�g�v��)O��'J9NH�P���eb����d����D���~� Ү��j҅_zݓ��N(X\��Ca{���Y[��;�vշ�Τf�K���+ L;ƿ��U;+�Y}��[$�N�!f�o[����v��˿��9?��m��n^�Lfmk+�׉m�	U��,�('��΃���}Ӻ�A�Z17�ǲ"ܒ�sk�c{�~)��6b}VW��(���|�t�@l��{�Ե�D���=�|e;T|GY��yϵx;0�_�7�d=�M�|P��H4���x3��/~��')���	�h1"��OT���h���]L��Q� �R+-Ig��eoxd�����q������\O�p���jI�L��b��Q���H���x�,�~	��m#�����S�g�4��Ѿ��dr�۰Bm���BL�k<��	�Ƨz�����0K�~f���6Ȼ6�F��s'���������>��#���}]���A��z�ǲo�f\,�����G|����2Wm��3�%Q���ws�
�fV?��C�.�+��N������x��i�|9�`�P�g�#��b������kk���yp7���4��z��bF�����c�a� �?���,;,F���?ǶlYq��kE�y�׏q-�KV��Ғ�{ٵ��_��&B��k�>SG���d��⣒W�ױ���B��Ff+S���2r�������w���?�񨾉�M2~�m����l��8m�d�� ���,W/el;-����I<��^ʋ�m�ɽ\a��A�㼼��W��X_����LFq�߬v�|_nh���#�����W}����>{��iY 0�SyI�tI��q@�Y׷�W�����W����������p<�ՊĊ�*�� �b�9�,	t`�W�lrƇ'pZ9.@�k��f �y� bC�N���'�TJ�]�G+�-�z�&�,�-h�
u�go��6�3<���K|w~�,UGN@k�-����(��["X1\~sAYm���t��L����;T�w���NZۙ�'�z]Q���#8�vXp���ѣ!��ɘh� �~H�k�9"i��	�X����A�ؼ)���:Ǡ��{x��7�_�?�j�䨫� 9���^G�y�:v#9��P�х�9:-�o�}��:�*	���.K��Zʄ��;�Q��M����w���[�w:�3��~��=<)��$}�G8j�[^�z�����<��FyÁ���Qw�:��_̣���PG���S�,�:�N��c���m1'�=k/��q9F@;�D�`��%�=ʤ�����ޣ݈����z2��_Ԃ���_��[Y���đ�'��`�Ԉ�?�$�~�^�0�h;0�#@��*��P��`y�WLY]����u�`F���}��6���RZl���l���Y��0�ώ�ռ*�s�8.
��)���;ʺ�;#V�2��]d����؎J ]0��K]V��w�X���w��8f��-��^�k;����]���}�y
Ǝ�q��`�&��=����[��D�0��D��(�Ҟ��>;���泋|��Z~��Ņ��X�צH7�>$i�<�������e䔷���b�gw�[+�y�]� ���]�g�FJ?Em�tE����	�c���hL�1��nh>#\�'�m0�4�g��m�]�Ivr;�n)w���4đ`O���E<�W<�Q�Ђ���E���cl;�?�W�>�;&!>����wU`�GT]����)N9���V���<�4�vm������S�="��z�ܖʮ������46qRN�D���&���I}�4.��{����ڱ3����D��HW�;�x�wv!���Iq+�9�=�ˏ�+e-���q�����c��D�qF��ד\k��q���u���|��{ܠ��X�g��ʅoF��o#o�Y �8@x��<��3*r�Pe��<�~��T���m����;���쉔�a���EN��3Z�tq�'�������8e���ۋ�(���;z�u�����O���	���ˏ%>�ٞ�a�eM�q<�#�P[���<���,�{�:,�=5��l;WcwP�J�[�`�x7�5��VM^=��������w���pux�m��S�;�� pI�tIg�7� ��N:.�u]�'����G�>z��ݗ���ӱ�:����d#�9�N��/�c#ࡾЌ{+�@������we�,���Nb�6��4ڪ+�kac���t8=;��vB�䈰�)S]�K��,��A��0���Ϥ��:r�":J��Xc��c� $��$� ⁝dA`GA^t� ��bu�F��+�-��bH�6k��B�=���;��K�m�\�KXE���:�%����~E�{T� x�r1��.�x�>��}$r0�(o|�:���Ȼ�!G!z�1�or�X=���˝��8l@���O���7�7
\�op�I;������^��籨��.�:e�M0�L�m�$B�������# }�[�����4ئ�K@Kc����m�`�/�����޵��tsn:�D����>J=޶�q6��:���Ƀ�WY��5粐4>�h�\�vDv;��/�Z0���7~��%�Ń��^5cy����@\@��>���7jG�ݓ�X��w@�m���0F�V�x�X�$@�;$�fu�F2��t������3�8����8�l?�u+~���c�]zm[����1�>�[�^׋r���d� aD�Dς�	Y�!7p?��A�$#�mh@�n@�e$�K��r�l�-��[��9g���H�Ȉ/�/2s�s�ҭN�q��k�9��Gdd��̬r�Ҵ�ss�\�B��c7�6<�{]�J������3�wׇ���]z$zb晕��}-g�U�޵�z�:-Q|I:?r��.�r�w�b��9�Ԯ��5��ش�\[i��������3�]�Ү[-���Z�}��J�Y?����m������4?P�Q�v��X�� �q�T_�O!�x|�6����������3ȁ]��ꀨ5V�;T�7�Uus)����-k��p�&_N���,�Bw!(>˦�a��L����ǣ��Ӽ\��9�Y�Q;7o[���](vs��ܭXb�}�f�w]�\�ʨ�fW���U�Ϋ�����j<��Ah�;���ڜ�lMz�����;{YYiP}9�Pǿ�H�R�<�>�]���$=v�F��V�L$�v��k_��6�a��\�d-�\����B��n��dw�U�/��s=�g{O�	�.�.P5�!�^ګ�|VCշ���f��?&��Xiw]�����AM߅�ESgmڹ�ͯ���M��}�>{�hd������g��ϳޛe��ON!>x4G4ie�K�V��U�/%�}��Yw�:�Gp�]֥xb�s������m�:͌+�U�=.���̼<��Ok��~l�d��ɒ#(�z����D��Q��߶�AZ��PLl ̥�����c�ټ������r���sL�J|��)W����߇�m�i#.�� ��z�U��r2�<�;I/W=$Ik�;Ę\��r\v0�G{��2˿�6���2� $8�l������Y;~��ݻ{��]o���-�k@��*�~??��_�g���o_}�u38��"P ��\&�mP�8���[im����k�:�:�S�p�δp�^�T���/
�DS g�iJ��R������jZ�H�N�
�� ��FU��+(��g���T���Q	�D5f�X������e��Ƕ
�bқ�l�M=;��{���j�D��'P#�_����'V�g}b���:y��H�7��Eڞ�#�Ҷh2��j����Ғ��mHN�ϗ���A5�wB�1��7q񡖽w�pW�5۷��B���,q�w�Kk�t>z��I�-�e�#~���S��$���5�Y������l׏!�W>��fVh���~�O�p,Qe�.�t����4;hu���:�=�$��4���l����>41�86�K&�M�����zL�nm,�eUF���"o`���+�k�v��#���^�ԛ��?D����Q��l���Z7ue�7E�\�<{�3HZĻ�td�6\��rՑ����=�U�U�����iܺ���Ga�7tEE�����4�+�֝���:V��8a���ȳ���쬞e��2���|��U��N�!Ko7�7M
�+�+�c(�z���Y�����{�9��������y-��<
����e,���e�J^e�^����Y�2�%|��ݙ���ٿ�[`f6r���Gל������k��q�Z3�>�_�Q��e���̳�HQ��/;G5��#kݫ�V���ⰵ��>���ߊa�s����:��|vmKb�-.�V>���]��^\թ5�䨢mx�A�~���-t�ӑG3�V=����I�k���8ˤ��X�*���e��l�����KL�`��W��ܓ�/�K��X��9�Rx�,�r��n.΁�]0�~W�[�f�sT��.���,Ѝ��43~x�?0�5�D�O\�lK�3�huF���[���U62`r�����+������v;A��j#ؗ�/�kN��vE;�D'��1�P2%��[C�_�+yFV�^�N^/2�U�$�N�U���.d���W��(P6c�jy�f�?��V�S{n��+���gس�xQ�Y����4R>��7i����(����	b/v����Ҳ���W,��鶎k/ײַg�ee%�"W^O͞�Nmh�Kx��pƗ�/�/{��t�e"���~^��U�f�q�qٺh���.���+�v���}r�Ҥ~���?a3�rW3}�>ߥ=��w}�sf��.�>쟉��EC��O�+��W����~�f�j?�Xb��E}#�n�1E/��v\WU!�>Ǵ����{�_Η�����˯[���x~m�G:s��z�ޮ�+�ߏ# ����'_?�������~�7����w���y�p[�5�B
IUZ�d�BX�T"h��$�G=�6��m�P�QT��=�lQ��D �-�8��}��ml{+��Z!�:(`�� �
7�n!�vSѪ!� �I?U!��#��lHT���]��
�5x��@~W0�}����<��\���
��h���զ{6�c���N��Z��ޮ���2=t�"��Q�lR�л����b
0�2�8�.�dXN�@�x�,�]Y�j10���x�H��&09�_����?ղq��40Z���=]�RhǾ������ֳ��0�+^ض��աS�=���k0��$cd.L��¶t��%�9���Bû=�xv�}���p�:f�а�2���ų��FW��h[��V$�U�9��i�y;�Z_WY��?�u�֪�( ��iu�2�ܭ4��U˧Az��)j!���R��?݂}�9𯫼ئǫ�|���+
�0�툹��~;G d7p��g'�ٜ���̔7��4|1�g�B�2�	pL1�e��}8%��JD�F�8'���w4qrH�c��1����9�2��V�;�ks=�ج-����sk�/��`N���-Ю����)��� e�:�f��AB/��}�s}{�G[Q'��c�3%'��uv|[>�o����(�G9�j�	t�������D�U��?Z�i;�a�W��^�;7��I�6�"c��ʠ��i�@�/VQ�c��X��Y���䱚�V�[8��8��+�X�M+��y�˜�z6��zA�u��,i1�g6t�[�\G�4�rB)��O;��T��ϔ3�{�]�4��2��`1�;���m=�x`=Ae�N�+M�\�9h�j��Y^�&;���_;��1y�R�,�.�PE�sV�Ŋ3�.s�{�ij-[��F;+��ҟz0ɧ�J8Ƨ�ع��)�]��l�"kH ݭ��t,C�8?����m���sG�jT��27�N���xW繎!�,��F@Ni>�v_e������;VcNh�ARf��xhǿ���}�yؘf�+s�t��:?Z�k��hU�IY��
+e)t,�zY�>��oV�y�/;���i_�CE-����d'?����[u��}MHf��������ƹ�xW�6'aT~�ޏoS}�M�g���%fmmy6�9�0iP�g%5��"	�lN*	0��{(�%x*O��un̻�=PA����'�c�Q�#�{_hY�:,`?�Z��Mm��fr�'�op?7�o�@3K�7y��1���)�^����U��X �)a�Q�z ��� ��!��4�\���V%Ɏ�^&*Y�\�[�f�i����'>s5��IeJ�~���n�w/��������_�����?1��=���v�]o��w�%���}~���/���ޯ��?�����y�糽�3�G
�3��$\��a���30��&�r��z�}u@#֭\7�.`w�����^�|�X�ߢ?cw��$��d9�5��hTQ��:�g'J���D����j,�G������R��O�~�۬Y��>��7��ع������F
r��3�A��E�,R�ҵi�+u�*����ѥ�/������e
Z��m�����L-+���Gl2�W��G���0�ۇ��D�	\�M�}W�<�u�i�h9�����	cş�9tT����;�^,���~��-1�Z�90�9�=����W�:���Z �i�խi�b��. ���.�W�}SG�RL��"���=��dۣ�����m/u�_V�����7��]��m ���~���~v���:�7��U�ަ��0�^��(d�U�t>�Y��>�+�91��Q_���$Yׂ���'}y9*��)�z�욓)��vƪD���A�#���C(���6�!���S%��m7�*�}>�����[�X�8���:��B���˺�KW(곍�"�R�����<m�=�Z���K��*w4h�ET����=�h���1~f��Uy~�_������>�^��l�9Z�����������,��Q��0FY��>���c�U��t{\�c�<_��Z�yB�,��)�Á��b���2_�]�G3͆��"a����{X��^�q!W�u]#]2����kyspɷ�=Jٴ�kN۷���6V�m]-��
����심@V��T��m�,�\B� �⬚`�����^�C��-��9g1t���QnP�s��-�37���z����OCo�}][�Rl��?*�)m�W��)�2�#��{����'�,��vsI��1,�BZ⬞�oA�u�	ʹ�B�?�����[���ғ�Q~�˚q/���6�%oF�S.i�%1g�öhB�*�f=�.;nc~TA:��>#�i�>�A�"�`��)q��ؽ͹B��<?��Z��/c�����ݺ����q�M�������=�V]���,e���<Y���k�>�ɩM�y]���>�f����S˩I�5�X+X�V����M8S�I�8*���:�ٶ�(�ӽ+ٵ�E���#�^��>��o�y�hm���{<R��K�L��,��_�)��Ƥ�Y�>�~Ӥ+u=�Y�.cVe��3�O�����K�؋�9��lm����_� ��]���<�t�q;�K4��]�V}�~1�`.C���mLb.s�1��o����G��G��[����C�ɟ��y~~��{����v��v�]o������H x�g���g�����{����ΗO�~o�̒��Tn�^������u�u��$��\�Y���n({|����t�!S����-2	��*n����F�D�\�o��*�]�.��l4OO*��-g.w�}�I+(X��=�U���wi;�����l�{�n�{^����o	/&��>�7W�j�&�l��s0}c#��ᬻ�mj���ђ�w�����CQ@)V�����.�܇�A�� �9�1�л��ן��̓B����X�j�k@Z��PM)!��M#^��)�QV��G���*G��Av\�	��sg})k"��f���gǗ:Z'"�6���Fv5&wr�۟g�-����j���N�SϚ�o�>�o���VW�ɘ��B���e�<p5����Q�V�4u���;�G��U�#��E�������N�W״�Y?T�������Ag�,���(sȇÊ>mX����㏹�������-�K�L�y�YE�Yf��� T�iZO�͆}���+���cV2�9�]���I̃ ^��s���	g�{���9!"��zk�i�m��EG�WV�ØV�T]iС{��%��2�;^1K�{q�t��PA�G&��o���ǊX��mJ��֐Ҧ�{���)�~��a�	�Ď�j�)uw��r� @�g$;��	l�֛�OA�g�US�|=s�/�V�o��˕:�[!��Xw��ڔ�]�TƢټ{Y-{��@����Wd(�ԅ5x�����R��}i�]<�xB���k�,�gbS�Y�m�&��&�d�K`1kr�`�㻝s����	���_� ��9��&	X#Q׮;���Hm�+G��4s��q?Ϗn�W,;��A�-m�u�8�o���i��m��M"�骁�I���JuY�y|�=�V��X��t�|�[/|���W�I����#2"�E�t�I�\q��x[0�����G�s�.�͕��*fK������gJL1��q����>NY+eȭ�s�R�����B��Kx9|��񤓊-���@`�Hj���I����Q�̟|���Aa�հ�g����`��~���]�iC��/�*�n��A�m=�"m��~��֚��Ue��C۪�2�.|�N�)�sN�-��ha���Ծ�*��H�� x�lymw��ܙ��)A�5�h��2>�w-eΡ���@l�w�تN����L�b�o����Nܼ�J�}��	�i_��2��&����i1�����}����5�ku�]�ݣ����G���2c=
Y�]|o��V;`�P�b|�T8ut��&	V�裏����uO�7=Nv��5jE���o����_����������/�����������/_�{-��8��z�ޮ?H׏���������O__}����;��˻KT~uDv��s﯋[��ip]7�CATKcBtky�_��h�!+�+l��^��uZ�����9����Հ3�'�{��{�@#)n����pb۞�8|� A�@%H��S���1���J�ڷR�s٪��6>�hu�@+ ����{����#����m2� nV�.�>�3�k��̰M�j��ꦶ��-W#�����~LmMeL��դ�D�E���vȖ�+# ���z�;����x�P�p�Ӡ��g�g�.>&^������q�����h���:���$�lS}�o�J}�n/��.�A�o�tj�!����ܽ��:����C�΃L���8d��S[Ӂ��������r��hS�Ŝ��;�;s۔ge΄n�gUV����;��y5�8�P�u#������i�N���\�B�z�9�K�Ao��_�� �\�q;�lO��l��܊B�Vڷ���`[�0vT�����z�W�@}��_;R���Ր�t+q�<��P���o:e�j:�������Z?1 �綶�4?�۴B�	�8.��j)��3�I�6������ ϋ����y��K��>�L2���� m&�>���wrQrm��� ��)(�Uo�Yu^��Q�蠫rA�-h��;�K�"&��c�K4|r�:���>nR}n^��Sdk�옕�y��� i������D;(�{�_���O��*�s���`n��9&z�@�H����<��K?�'�����؎I�����yi��s�=l*ɩ�[]���__�k��ò|Q�D�9�o��خ}��<ţ���‒h�k:�ٶ^����q��D�c{F�+e��zq�,+�$fp��}���EnC���G=Z�s��Z��^�>w�����IMy�z�a�6�gh��펠�������nݴ�5�;HY�6�����!�Ԭ�0_TF&~l��<�3i30)ӗ8��!�Ab�#e���v�I:tХW^���%9Ϻ�A��vy�U�� si���z�;��q�꿩�2n7�y��C�+�e�8����6���=Ϲ�s��y0���+ܡ�,0A����cL�[��<�T>��УQ.�-���Y�������ejPjO�:�����+sʔ�jpT�5��~�Q��9o�YjD����X�D�J��Z�S�b�`���k�b?��A�rl��+���Vh`��E=����W\��^#o�|`K�9���)7�����W�:�s�H��d��b��-�y�>J<��:(��ՎN:L|=�ƶ� ����͠/g��§��-����c&`�7̓ �'>z����c9�Wۡ�Cwl�g�9f�񂾙}����+�'�a6;�i2o���������6�}_ v^�e�=��M����f�պk�ԫZ��5�8m��
�u� ���{BƦ,��W)NK���]��@f��˻ðX4���"�˝�GGIV�hˎW��� f{1�L��h,�|�Kڋ��q�}�>n�>�O���޿*�O?��߮������ ~�U.��'�����;���o�-����>��0;s�g�C�� e��b�U |�a�+�V�8�)8�/��.� �pbV�J��M�[�EM��\ڳP�����@ �B�Cu���]W}��F�N�W�n���s�����p�߽~�*���e�M 0���"��\A`8�`�y�ON�� uPڄ�3�t��;�^+�@[��XT����	EV�:��6I+m#ݴ�<w\�~��#K�Z���@�:���>�;�S��h5���-�5#���Ӽ�@!��劎�X,������>�:N4���"���5xrly�LM��Q�����3���3����<O�%���
�ʫ���';p��q�h?݁�� �Պ�-e�@����<i8(9ߔ7�{#߃����}u��*�^�U.y.cݞ��ev,��f?y��S<τ�H|�uL�y��C��(��F����;�|gu�������6}��8�j)�����6�݊����� ߏ���3m�[p��L���㐕2P����N�Ҏ5@��Q�-���v<��~UVŻ�1�a��+u�]�__c�z��dv^��`��'�`��צ�V��vCFI��ߍ�-��:�*�K�E�|�rk(o��
�L| |	�x�l/dx� �{-r^p����!�����G��Oq����!!���^���_�$����B���4]�Ѷ3����d@e�����1�h/x�8ǧkBV�h2ӂ�;?���zU����p�m�2o=Z�񜎣=v��W�U�."8VZ�*��ɴi#��l�rk���!�z@���JF)�f����a�:z	�Yۙs]��>�g$���+0�.2���'�C]{,�`�T|��?%�1ޫ�b�7l5�ΰ�?w3����X=o����뚱��� >s����z�������`mu����0���梆���3!k��,�|���5e�X��hǾ��>u���~\���@�c��C��i�������A�]՛�Pe��|��0:|�y���'uێ� �n�:�9K�m���~���"�Eu�����a@z|?� �D�me|�?!��_��2g:�u4�3^,�$�ď���7U��_-{�T٢�o�Z�w\8�����<��9�.�N�^���ńf�����ت�(����y0숾`^���^W�5�g|Y��^.u�#m�6K���Ͽ�#΋c��J���'�6`�����]CΓ6E^	��"�[+u�넌��cJ��Mq��35����3l�n�Kg��x��}G�g���������Ѷ��U��Q����Xy5}�F����Kw�\�s}�iHG"�e,���~�������͊��W�G���`y��h~��:ە�lߌo� ��������ZbD��:�@R* C�z��<�X>��&�1�����]����q#�Օ����^^�|n���t{��;�������v�]oׇ�w��Z�����?��O}�����_�|�����L� x��)�RY2�܅�n�J�:�)�{�W����M

&�D�2�- �1��]�}�ƙ D����h�:P[�R�x�����9��l&]%��l���� �l��f5��~�G Ý,�^p6�X��:C��w^M��e��\Q����A�m�.=���_/��Ȁx�Z�n+>:�{g~��C���Օ��d=�8���8�{j���\��`Pj��q+.��ma�y�~��������I&���:���\���#�;���ZA4�:�>�vg���q�j<U�Ϲ��t�Բ��l�?��SZ�'X���*]�<���˻@��;׵�u���m����e����.�!n4`������N�>M�X�i�Uz�q��#��z�``�y�z�ԇ����o�Miæ�(/4h��#e��A����y�]ydo8�9������T�����9�k w�-g���ʴ�^��)����l	\���7$���sD���w+������*35��y��-ty�f�,��dҀ
�9�V�VJW���ShK���M�.��k�Br����H��ޫ<~�Jb��zz�J8w^�����]��g����n�w<�t6�q
=IC�Iy�:Du��Ӟj�oL�uV��e������΁Zy�c�xU�t�k�i��:O�}�<⇝<�?W]@\��؏di4�e��5�7c�5�tb}��Z�|An����[}f�5������۲�51�v��G㮘G���/k��M�z�)�������Y��n�#8�ʾ��ww�ew����B��L|gk�w���=����%���4�O��#?�];죿��X�K�x׆�8>��h�b��M��[1�e����SOO�mݵi�1�N��i�J�uQ���q���XǑY�7�0�6�w�*�c=�:���JW�\*�����P�J� 3_u���Q刎�1�.��3=��6<�6U�!���f��*��_�>�Mn7��92tj��E���Ď�m"ݮ�t�K�+��ڟU�<�)3���[�:��yw<4_5����y�f�����:�����s;������G;��5�G�q�o;�zc~~��*m���}]�����y�*{mCg��L��4���;mK�v��Z���w�{�#��ٍ���#��qL�N��Y������_��_dL�DK�;�]�����N��u}��lk-swq>�s��u�1G;��XO��A��e��c�u����D��97X�E�n���uW�x"�7����1�n�=zd��_l;��Z"d��+���}|~|����?���������?����g���9ޮ�����~�~$ ��ӟ��?������_����[_��{�������)����]�ճ�"t�s�~���`���p���M�'�NFU����PhHF`���.��Dk�k%�#=�SA�*��Y8E5�bLc|y_]-rU�{_������=�w��]��O���D�m���&�P�c3x�`N�|H{+��f����Z7��C����ou@ʂ���A/��۞	2�O���F�Ȃ�.�5�:GW����!��b4��H���4C��<����L[P�Z�Nf�b~w��*�Fݤ_(�BX��f��hdxݷ�;c�7s��U5gV�����d�a���3����g�:�_	�t5��逮�������Љt����܊4	�ďs3�;Ͱ�1H�E��H�jz���G!��;&uYp֤��>2;x�Gn�^d{5"ɭJ��o���ֆ����i�R.+�kNF��3�?�@�/4mS�(��y�����(�"�sWP׻�� ���r&����舔��r����86a8��?U
��v��]��+y����D{��'j����ٱ�Wk�\Z��� ����h`��uΏ��Z���Y�m���.=�Uu�Ι���ͳ�~˺R��������,?�V<�΋}�><�+����C�g�u�k�������諜����\���5�<�:�o�P��(+Rj;X���ʼ�L�����#;��B�#Q鷣鮎VA]f�i?uv��i��U��<�Xq���ͷG��,z����&�����.6I�l[d3�RN�ڛF��ԁz��տy�"g�����2p�������ˏ��xT��1'*�%�k�;�[��un$-�̪'�β�w<����,�R	_�r��<'� �U��K�2O�a#p�[X�����3yݴ�;�~����־̗�e�g�KQ����Zc׌	b<�'��e`�D���q܄�ز�Q���1���]'�G�z<a��o��\��I��M��v���{{ ���F/� |F�����\��ڻ��d
\n���V���E�����vⴒ ^ky| ���~�v�q�3�a�.���;���hS�b�}�����ۑ�&�&��sd��C8æ��!���ɹ�ڎ��K{g\��.^:��2�@�Imu��m�SH*�z(���^Э�#O��H8~bd��}�����/?<|���+<�,wtY�I��������3��w��2T�����sSd��O��}U�/���(�e�57!?����Ij�qP�GA�b^���ëM��`�Ȝ'�m�0��{�/v�؜ S���<�k;݉ŏ//w�������ׯ�_2I���Q�%�$�P_+u�2��Ա�g�As�l�?J����د0�{׋����ݵ}�U�NÍ�=ƣu�Ω���E�	�l/�/��cV��t0v�������=c�t{:>����?�����������>��'O���g�}��Ƚ�+:߮���z�����z�OOO_��?����������/��_͍��q�`b�A�p܇�e�����\h���d�� ����n�걛IɣM�B	uQQG�wfu��2x�d�8����\g�O��ň�������g�q�����4�iܐ������y�������w����>��c���h�U�:8W(� ���c@�{;#��j-�>w*�`&�q9��N��+pMäI]g� �+)�`(��׭��Q
в�:u�Q�ϼ���W܊ASqApuc���e�`]/8�hUp��rC\ޒNt��O�0J��0^!k���7���~�r��ԙ?�QI�G�K8�v����٩�˥�mO]���9Ҭ���v��kF�ҀF�-����[ywv�X�[yN�gRI��Gl�4($E�x6.��L�d����Ύ���^��T�5f����
��J�Ғ���<��'�ͺ5�6��\b���g�IgXO�/�C�ޒ�=4�$N���(tg�x�*N^8/��� ���;p�ţy�\����{:Q�8��F���R5a��}8@�{H�oHz28x�Sx5)�#�ȥf6����b&�>QB��M,}��t�=�k!�)t1��˪,��]�i�ܳ/[�3M�����o�\�9����y,A��:ZGVLU����Tb���}��u�!4�x�rX��qD�o�d"�)���W㈃+!lNȪ�
�:b�椎� �w
��v��g���;����ާ6����Y�Xu�����Zi��#���w�($'\�5ۉHY���� 0�Y{�z����	�m;������Z�B��"�#��4�7	p��;���݈W�����ؤE�Y)�Kg]�X�Lݙ�sr�{�y��ʘo��\� �O�4}Nh��g=��y_�(��:��z>�Ok�),#(�������c�����i�	f�"m$Ȗ�G؛]d�u����߉�.�r��k�q��`e���w��pl��UڤN�>ǡ��Ryw?S�?�|��˽���s�e_"y��L�,}�6//�Oy���ۯ+�ι�{&T�u�<�����V�
~k��+��z���ـ�[ІM�*轞c��Ʌ���"���X��:c�����e��/&�Q��w��N^b����cQ��s@��ie&�	�~?��Q��r�gK�yD`;N�<է�,l[��������^C�d�Oά~Vvk��� F�z��z�XH������:��j�.G����3��2����׶w[h�tN���}��@��{-����6A�."-e�J��&�]���&���,
G��rsp��PGP�^�1"�sԯUXLF#(��d�P��]w��rN��NE�ɫ�W���G��F����H:�nR�U�r�8u�y�	?f?����2��t��{�Es��6l�j3�}b;���������N�w΅���~�5���"�k����خM�9���/CBOsg�i�B�F�[72���}�d�>_�u�����2W��c�1ٮ��+C<��w���?���o}���o���w_o��� ޮ������ǚ �*��%����믎�?����W����������_�q���+II�4�&A��pR��� _*L��/nk�N�@�>]�s����dc�������U9I`����1��?%��/�~W�z��Ra��Ρ�&�������loE��e���=�=s��+�l\�]����_�$��O?�̾�ݟI �kE	^�9}�&��.A.X jQFo^�	/�����W�V�ZN�]���O1�P` +��8J��|~2J�G�m�̓hF�d;!�#\����<�a
x,]�l��=t;-�鰺�M@}���7�q�k�3 �A�@��4�a�|
 \o����Ɖ�2���" i����amI�y��1Kbbe��	�-�GI��Ҩ����ػ���0j�d���C�6��3c���̑L��#7�K�F9׹Z�n'�љ��"�a��I�U:n�<��AZ�1���½���6�����H }Dώ񟏾S����ڵCI������s��[:
E�G�5;�I+[��A�c�<���U{�8ݢ�V�>���=僳T]�x�X��M���r���1Ʒ,+���Eב�0�)�����b���0ӹ8x�)����߿���1W@��6��w%!�>�C���B�%�9O���v��U$��2�Rl�-� W@D߁g -��B�E��!�ʊQ��db�����Ig�7�ָ�D�c]`�t��U.���.L!e.#���O:�c���O��s�e���7*8bU�O-wdc��1��ㆱ�����夻T�U�F:���2H�q�q�~���Q��@gP�����L�%>�vQ?�^@��=�	��G9F:�W�p��P a󒥷��u�-1aCN8�y6��ͩT�J�V��!	*�[h]��#0�dt�7�9�c�IZ��9�)��G�Z	u�V�ݍ�8»ˢ��X�s��<��{ͻLz��D�ى�ۆ{p'Ƣ��bn���ҋ��ԧ���n�r[i�|��k���#px+������2����O9��{'n�B����P���Bg]f�� �
��<Y�(%E`D���t�3p���}�*�I�~�cN��k�ML���1�]��N�r�$���G�j�7ƶA'A�`��|�7uC��Cp�	�93��ڸcX�ޱR�h���m�c�?��vlU�QN��9�3�nǣ���S����TK�#��h��ZĠ��Svz�3��<F[}ת۫M�|6v�������7������d`�ۻ8�'pȮ2-��=8 r�6;���>����/��Ř9�Y�口Yc}������v&���x���zB�c.`gG(�䊜8Y���gB�3�}��v00n��nء���Aޘx�	�;��n2:wqھ��8��8�N���ﺺ_uk ��������n�P��I�8�h$�[��la��<9���������E���䋹a9$�����ۏ;��!FZ����	e����!sM��ؘ��zE�י�T��?�g�Cv�^睅r�v
�1�鲒�z����|���1Go���Rp��Ė�K`Dc?�'Ƴۥ�9�C��s7���.����i����[ӣQ����#\0X|v�����Mo�%ya��'��3I7�d��L���>7&?8�9;�B�17Ї�c�����Ē�1dʂ��:�� �����h�>�����ulԉ�#ү�����_����1��u�9��Gc�v,|A����1V�א�]��̊�$i�ﲨ����tT?�U�����g�~l_���>��{y-���n��=�{�B����?�_�T�{2��j�[��t�4��J=�,ߝ��AT�AR�=���buu>�/�S�����	�ȣ�L�B���q���Ys�#�g7bk(���������r��l�ۦ�?I6!h����/�O��_}�	������;/����v�]oW�~?v ��]����o��?�������ٜ�䯲��mU>UQa' ������ǩ\U��D������n��[i�G�3�\)����u�ЀbHu�,�P(s͠�Qşm	�]ٯm"�j=,�`fǡ@���e������]���}+��܏>��~�~�>����	�4����� wdVk��82���W���3�0m�i�j���x�u7�L�u>���u����|8�,~'m��Xv?A=�w�r��A1z��Ռ�0x�5%���C@����8�3ԝ;��\�r����"�$4Mfl�-%q����.�e9��"�O�r���ޒ�&�0d��~�j����u�+t����c+�rή�_�5:@����0������qY�+��A��4�"���15���pj�.9�ru���6떠:�����cz�#82ᓻ�?c.������,������ڦ�-�<{]����#1@�q.쁤����>/�ގ��=��|��A�(2Ji���m^��Qՠ�m-I��?�kr��A��'��Q�3�<;��>�^�p���m��f����#�z������td_X>�LCV��=�.XwAS�|:s�"%�a��%:>C��@<KG�lחE�9W�-Ap�F��ّ�g�8ct�
L�L�G�}@VF��$O�h7u��T��x.s�|�r�Y$��ĄH:j2�c�2�{#���V���B�k�YKG%ݔ��ئ��3H��������r�*.W�1���y؝B���Dײa�[O�B�Y���C<xi�F݉T�9����w�����C ����L�r��c�X=�/���8��4S�¡8��˽``�&u{�s��oxO��]B��b�.�)������^�g�TE%���Y�p��^�̃�������[-;�h�|GykO�ڮ��`��7��9:�/�\1�j�L�\.@���4k��5��c��h��h��VU�ei?sG��g8����3�k�U�g�	�J&t�^�m�;��ۙS�\�%2ɔ2���!d�-�́���^�����?�\���M��<�G�Q���h�_Y��d5�&�@b��=��>G9E���M����1� �6�eu�x���������>����αG"X�#��	۸��7# �}��4�-k�H�1�-���W���n�T3��v���,Ϥ�ă��qD ��{��jGݖڱ��PI.�C0Jg�M�I�q���+�5`�1P˹�xv��:΢�C$6F��P��-�G��Y�`+�l��a?(�e��\�yu��>h��2� ���j���D�;x1@�;�uA�S�` ñ=����[�ǉq�Ltl���7�%X�c����_�Qi@�����`�(_��x �G�en7`���GT����ӿ���Gȓ�9��'�G�T-�a�O��NK!�Fǰ��.p�����1 ��,;t��i;?h`6����x4J:'N
^? �c�s����f��\H�=���Y��jW0���G,�#���[�Ȗ���j�7�c2�$~��:� ��^�N8C�h_���ÛJ���Xo�.n�.�Z|����2ӏ:r̗(��^����u'����0 i��;}��|�����7{~��}��������GÏDl�e�uN|aZ��<��a7��t��Ք�T�/0;uk�\�2��1�,Hp-r!ڪ���S�j��t�ģХ)[sr{����M�)�����E��&�s>�|5P@����}{>���_��ﾾ�lT�o���v�]�ߗ�w�׏޿�ɿ�w���>?�}���|!�FG^[�̐^�D�TP��t��O'������!���!e�\�,���^�r�u��h���L���: ��v}�M��,y��*��L:k��P�*K:w@ �1���믳��>��>~5	�7��/c����sb�
��Gf���~����������ЌΣ�&�h�q`���:���>-1�����Ծ��������C+ʰ���78��V�sun���	��S�{Ov2S�M{��ӡg�����}[	�RV�w��8h�g���ot�ac_Х�ƠGןv���vb,l�n��v�U�%�Oh�9zt.�~&�oI��&
��F�7f�:-��t,'������J�'��g �̣���,�4Z����Fӻ����h�=�isG�=�,p ���]T��`�p�p�_0N��sׂܑ��zu��l�Q�>V��w�|,�F�0{�D�AG8�A�YG���s{��t���`��eiP�0�j��<t�Y��L]�@'��:�r:1T�R+��6Yv����NI�{�ʧ��uڌ��%{abW0i�Н^𡿕�z:�{���UO�gN�c�q���f8���Un��p���sy 'v���(�CVڤ'�-�)��]���T)�r4Ύ��y��h��I��#\5;
�Q&/���D�ݪ�G�O8�EΆ������S��<�֕o�RK�T;C�j  �6�w�������l8��������=���N�cƝ󂥣=Gʼ�[�
駹��ku�be�h2�c��Q�A���;�J�`9���Vޝ�C:"I���c�����,Se}��̖����!m��X|�չ�N*�M��ϮӜ���=7_�l���[-uF���XW�>��Ә�)µ/�$���)i�1YF�A�:U/�J�M\�r�qBV�uƪ�.����4�\6��U>�<��h�o��!!�o��N�{<��/����lOm���r%w�B�+ڙ�qڅ�1P�S~$?D�c>�Ni��ؖ܁�1%�����>P��ޥ|Ů���[�,X����I�Ĺ���n�x�ד�K��?"f�|&~����4Ұa(��K�P�""2�8�%΅=�ҧC���[��"7���c��v�l5���y`��4x���p��w=�	<{M�	w�psS����\��<�o�/c�1�i�'V��h�&�u蔐O�e,t%�,�5(*�F�-�^c�A5c�z$y!�%�^OR 3�����'RVѲ�H�~0�Y2O3`t���~&���|G�X�x}�6b���=�F�C.�I���;']#�J�#�as{U�����'��v6C���Ȟ�����p?O�t�-��La�\�ĉ,�8����
>)���$ �-�ĥ�)�B�#@k(�����a�?�p���cڑm��!��M	��@G�S��w���0��G��ȹ�֦�`g忔�z��a����,�T��C���F9�8F�^m��N�������Z��1((�n��g=u��o!_Zyn��L�Jz�}+�ҞEO�[�~�==����=��/~4��_��W_��r>�h��b:[�(�Vx����J���߫�I�^�S�.y߂�v��H�'���б''[�{)�b��ÿ'�r������ѹ��l����`zM�8�$Y�g��Sbξ�¯_?~�����{{��Dܽ]o���v}���& t�(�Oϟ���������?��_��w��u�fȬ��0�ec^)֪�����3x[*�p� �61=�S���\fJ�,]Ix]i�
�i�@��a����t��+��/u������N�X��&H�����" S�����3�)�w���'�~�F4pv�ցF6�y � �융��8HpFj:�'z�~W���6�}oY�Y�]�I0@H37�����A}un��1�W�"�H f���(��>UC�b[?�B[p����te`+d�q�}u���y>^���f����G�_:�q��Dj;�3��-L�G�D,�Yʌt����1Fs[q�#5�k� ��z�a�mBe��s0��vz*����a�+��<���{ү����^$��R�kS��N���?j��Fw��-�%y. �5�ruU�X����x�K�>�Rx����ᘐs���5ﱚ!WR�^ϴ,�tMgxn�}<��L���#;�r�^����Y�`'d{�w?
 ��@��Ϥ%V�^m��jXe/V�]�^U�P��^��쾟u�.�x���˸wȎBt�kB��ѣ�|�p��}�.
΁��nC9�xk9��HK�A��@&@��smɯ��lG@X������x>V�l�|� +X�G;���=�'�)7�=s;��{���)�t�������ٕX�
�d9��8�����R� �5�xe�ې�Ĥ�����|)|pĎ�s�\�ZV����:�r������s5�d�ǘ��W��߉ ;�ı��?�
M\���l)��^��9����)�+���P'�ٱ],�Q�׽�&r)�����;���LT��It�c�A�gz���w���q���g��cԊ��ܜ点��١���U��xTA�L\�6�O:έ�t��!Ws��/�/�`��d�V�~��h�I'k�jI�_0S���d}fyL4�q������睽S�N:��b��Z�B�/s~���l�V���
�\�J^i�56�H���N�rUǮy �[���������j=˩��9w��R��64�䉖�z/{�2tL���Q������X>��u&zUgʹ�+���r�6Y$Ή�(<gjǈA�K�)����;y�t��s�U���0m��G�q�����Q�
	�1�p��K���"���Y(�~"���K�k�1����)���.�"�L9t��-�����l�h#K]:^x�� a���A@�7�S����'VG;����X�<%�oф{�ǣ���6�Iowl�zQ�H��<���{���3�ˏi�ܨzm�ep3��||}�=�]Я�0pJ��
�cǍ����Mw��Bs'���?��@��n�;U��YY�3���3���܎��ch'x�� �<�1�����
���~�� �p]/���NY�Z��$b] ٤5�]�O��������Γ��9�iN`<n$I�)Ӟv7���$�^�c�8ڠ�y�C��݂6���EN�|��m��u?��@Y�J�w����M� �uj�	ݐ���,d9�P��W��%��ǧr?E�B?�R��~6"I~Sz4��w�*H`��	7g?�f<�2��,�����9�&6c��!�B�;�9cw|�K��y�h�.lH��kp+�^�W=���¨�>:9
Mw��-���'ٻ���˗w��=?cG]/�eb�M�O�^~��c˵�w�e��ղ�i"�Zn�o.Co32��=��Oxn%�&�p!��)�4�;ZE�-�l�\���X�쯞��P_�b�t#�tɣ�W9�5������w����������|���_q�����]o���v=�~�; \�����������������=�n�<B�i���ɻ���lBu��
���� �;�w�{<�mϱ�ŷ���:[U�P��q���Q����8H����t�$:�3#��{�ړ�|x��{W���@C�+~H��;= �3+
�{8��ÐT�����SlC��1���E��mU`Q�A�	�(����J�ٱ�V2HP�B�������3����e� ��K�K�>�>�f/�?��./�)���qF����q?�3�.���:}a�z�u�G�%�u,e��h?�����)��8�x1��Z���I]n�<T~C��yZ�}_8h��*��3w `�)��x���ك9�|FP;�+��[%���c;t�2�}++N�y\�!�
M��ΨN'�^���h�mN��3�Z��gl%=�#���;(����1/ ��0�Vq.�,?��Gs֕� �%�q��5��3A�c�O�+,�:���)%P1~���M�8Vq���,���p�"�ix¡+F��� ��4V*�,�R�IO��T�[I�8[�"�
���NXܾ:�����6�0
l�;h����J���yr�h3�{�%�q�A��:��E��)�jfy�7t�6X�'�-�.�I؞Ջ���8��*�Ҁ0�4��$�a��L����J��疁��U�}��9�*�P��u�ct5�#?D��.!#��<{n���ӠG��R�?��3�<Oa���=G���C�����1�_ub%��"�O+���z����dz�m�Ù2�5$�P?C�d�D��:�1Vn�|����L��aHy\Y�������z��O5��}Nyuj�Q��sY�9��M�e�����ย�2t-�e��:>s�I�Z�ò��gfKz��5�u�o�����l�M�����������B�Oo�`��7���1@�#�G������$|���<��M��@ۑ����dF�Pgiv�j�C��p�ic%j�F�J�F|�g��/�y:n:���+zv2��q�^H��|�_n�.rz��ߴLY��v���z�2�A���%��K[S��L���)�E��U�H�QN%a�`��O���Z�{�t��ðE�����-��Au��6j@��ֺU�(/�U�a�}�<���?�(�HX]�)y�!3BV����̓]
�O�����zK0r �������Մ1�~V��.�<���;\���h�q�D�Z�W��Pv	9s58��M�
�ɓ��+�N���:c>J��H��8
:������>�ف��#�}Wy-D;�i�H��XI/EZ�#�Ɋ�`�쫘�ؾ5]uެ�g�θ캀�f�cߙ�Ԓﳍ��%th�W����r>�C�ݕS���9�ۓ�Y�Ղ���RS9�w8c�'Sve��M�Q$� `�<^=�ǚP���M����~���}Db/�o���}��]����I�~�̤�>�r�]g�>挷�\;�����9��>F�JLU��?�
����!=,c��x�΍��.s�V���~$�WQ1l�}P|�ԯ��@6��櫌U(��lZ_���5Sm�����?|;�-�E��=��G�]�OH��D�ǂ��x��X�1��K	�x6�]��I#�Kbb[�n��l����_��_�ſ��������_��W��������@|K x�ޮ����cO ����������ӯ~�g����_:_�?�D�˻s��_@��(gu��Y�u�q�Jav�A^Bŧ��j��ޟ}��7�M �lggnO��{y?t��z�����_g�m��Ԁ@u(*(^��P���߬�OZ�A��׃vb�� *;�����+hM��. {S��^U�
��u��-۽w&���ǋ�'h�Թ�9����:�ځ3���~n{��)��3i����|�߫Q�[lw�8�,�M<�}�ga���^̦�A ,��f�Y��;^�
� -Z��օ�����Np��������@�M�� i	N�V��A��m��Wf��:�������иR����΃GF>=k�80FyL��6���WG=��
��m[<~�-�X�_�i'���س��VK�_]x��_����C�,���� ���<��s,p�]Ig�3�N��?OYؒ.����40i��]&��-�n�eAį�/�F���6�<��LGX���9���uvν�ȃ�6�E�_�2�/��`h������N�:�>��O��D�ˮ�آX��o�^_+p�78�<��Al�I��@D��s����Mq6����~�֪�>�2�zb��<��������\��?y�K��jk.Rs�s�*V��9�@��`FD9�E���#�N{��Y�����l�<� 1��ۘ�6������RO� m�����I��ә@Iq(��Sݔ��CQ�������p����d�1h�[�i�}tͲ|�}���g��6�I�l�����ig����:���{��:��3��Nϕ�����%�'g?�*��>���}jV�!.�]׉�C�Y�c��M�X�a�|��y�{��޹��̐��\�QO+6�1�;�Ց��;G�7�c b���Ё!� ~�j���s�n�t��'�TB����n#�7���hÍ>���{����I����OY�g�w�HV���$����+�cU�>��b��.V�x^��NK=1�u͒�pp���!"�2��õ*��գ]L��R���̛֫�,�,�[*ce�g2(Ԑ�$�5[������oÏ�;J���䟬_�h��Y�XZ���X�D�2l��&&��z�v���u��qܐ0�4����������$3df0ǔ?�<��9��AW�����Dʔ���=q�'��ߩ����J��r���c@���/6�b9ǽ���n$ӂ��Mb�A&��d�3wN�o����cv��2�fĠqP&"�	v���@��<�iW>�1N����4\SЌ��~��FU�Nxl�����mfk�i�b�?�:��y.s�Cj���n�>N�>�n�>��U���^��6+m����8�v�i�����K�gJ���J�ܘ\����D�?	�*F�}cJs|�c�6��?����<���x~�g�G��nǃ��곙�6|ٜ���qKK=M.nr�떅���o� �hLw���S]:���. ��3���$�������/py��_Y?tmX���q^ʋqj귍�:���8^-�?��*��z�A���V�D�#}s��x*��~].8_��n��x��<�~��t��w/���7~�W�������?��w�ܿ��>~}�������z�ޮ����cO x��n��壗��'�
��W1v;z�-��+ϔ5#8��J��
�`G�E�2��������+�v�0�m<���-qHC��4�h�E*z*�4�����Y�F�����}��=8�J��5�i����.5��Ykt(@#�𶽼�j�4hzҝ����F9��|@��M0+^8E(�g��ۤQ�6�lq��Ju�+O������!-�4�����E��y�
8{�g�H���t@�1���K_�hn�ow^�����h`?u�_-K˞�ߢA�v�U�����;��TC	�9�
���}g�$+ހ\�Z�j�j�v�TyS�]��f�x�gV�=}4�9��-��xf��ϲ�F�e�nk�̫Np}¨��m����ڝ���7��P&��gc'l�;����p8s�Ӗ�|��|q��2��-���d�K�A���rtƉ�Ew �S[����4���@�VM���ې{��*B�%��nm�ӍP��F�'qf��R'A��]`ҝ�M�Ξ>q�_��;I����Lz�6�p�sd����Ve��=���H1�����Yna�@_�h�:��>0y�+_M��^1c_�|�r�^֑狣��N綒�`�HǶ��c\S7Ǽ��GqƳ�φ2L�k�M�RL�T�0�r|�e2�������=p�����ӽ\�x�-���C��UR��W�J��	��H�ǔ�3��^����!Z�s]��gzē��3�h�ϫ��3�ڊ��Ѩ��>=��־+��6 (��A���lY11���Jg:��K�ɽ�P���J�����L/`JŢܽ�����|=z�,lCl��!_��M��N}~����ݳ�\�)��c"�8L�;�����ϕ�����?��־�����f"�ZX1��N�j����!�������f�F}L\����=��I�h�x��Y�j3�.RĖ����;4���=���A�����?��Gیi �.��8v��lV�\�@|ø�z�m�wo��)mx��ĤM��IC���ۢ|�Z~
�sK}5g���-��55�V��3����zF�d�A�8chl�8 ��_%���-V�;v�`��, <t9���oY�/1�O���'�9@#�GI����dNȱk%e�Ñ�L�;1���yf��W�H��D�؍�	I���G�J�Uvw;袉��&cM���К�΂s������u7Y�9Z�H�v!�L0����d��%%�|��ژW���;V}:x�h��N�N�����T�ϸNWU���� i��1b�Q&�f�+\W��	�:^�]�@@��6�r���,��DP6�S��������������������'�Ж��muG�Y��6]X���k�	��쟧��CW�V�����|W�ǚ�B�a'����c�#}t;�a]��������q+�U��ܪ�i�	Wg�{a+����t�1-V�K����
1��t~��t#mu>L%���=��7KGi�	���5t�����Y��/ p�V��Ӝ�3��,c�&>(v�U>�K�Ԉ��k�����~{��ݾ������u._Y ��3������v�]��w��>���>���7�q��Kt�����^n� h��_'�x,�Պ�<�#j�qW��q[�ޫ��wC�3����M27Eg�9�]��=���YC@r�x�Qc�Nfk� ���g�M� �Z����df�7�Rϱ�	~���K��O��>��
�vߡi�N���	޲tV��5 ����a9;2	�7������tFA���uN�f0
"+��lC�
۴�,��l��M��F�O*�aYz��:�z	&2u) KVB˵�.^˪�e��������q���f=5�N~� Dm���Q�fwq�S�4�XU��r6�1J5���3<�6�3����^�c}�tF$��s�ݲ�,�G�W��E .���Akp�0�%��A��Χ�p����G]��;y.�e� �eI�_xR+��&oTYkaZ��n�]���gx81�'�T0�$K:�sf�ј6�=����� /~�U���XyΓ t+I�Y�q(�r�J<:��a�����ww���=�P�Ƃc�>���K��A�3wJ����~��c�b:�s�(��	[�'��?R����K�y?����ѵ̍l�������S�����3'��g�j�>�3�`ٺhS8Ҩ��+��A�	����1�BPE���$Z��:&ρ�m���d�n/[k���E�/z�1�}��W�GeSϬ�u�Qv}��W|g�-�����ª�vL��>�^�κ�d`va�?#���'�=&��:W��s�B���?>���}��y�fy��گJ�ozv�u�3p��m)�i�$�^��~�-���8m궸��{L��P/���YGt0�#�:0]f��d�K^F<{
?�T��6ȴ4[�+u�#��\����u���sw`������[΅��r�.�Q�</c{��>7Şh��zb����Zy���A�>��k��n�3�2^ĮA.ΫI�C^���9��U�s�:��+蝅A8�:Ǭ��Ş��NٍF =y�`�$α{VxOUtz0	�9�u�0�î�O�OMl���Vq��
�X���@`\b���ց}�l�D~��M��N^J]o�2WSŸ���A�+��e�PN�3�;~�~�Rf+V``�I��E����G+�N�F�mî�}�L
ٮ���+Uޥ/
�'	���L�H��m��m����9��潮|�禂�����xH�E@K�溰ۣoG^1t!|�Ǌ�HC�KYg2'S��V�wZ���*f�B��M��R�qF,�C~%���{M�DY��QO"��yk}u׿&�sƮ�=�/n��I��R��$7�ե�U<X� u�����v�+Ʊ�,��т/t�/��h?�fݫO\�ǆ4Ÿ�3H<LL �;�o��͏��B����9M>��؏��b$l锲�o�[qd�	|(IcF[�Xz�!s��;x�m��L����������}hqӼ�>�6��q�N�L�m�lkzdSM���B�
ht�(����0y���g�v�v��kk����/�?����Ң���z�ޮG׏;�������?�'��W���?��?����o?���Kx=��e��4�k
@w��l�8 $��Ƌ?� �/�
�y�=~�p�ړ[�}t��*@Aܿ���}������ H�G���/r�a~��������5x��4(�vh�ׯ��/��w�ލdI�XS�OV/}f�Ӂ��ؾx�[����-�i� �� :�PR ?>@��m��QG�6�#�`�V/4��/4� �i�pl��RurW��ت���s���:��@G���/G�Jd���t�j$خ�� 3��y_�痁�j��eqvi��F���Q� 9o*XW�֫8��H�#t���=Vv����B�mC4i	։�����V}��p}g�,g��æ�op��|��D7u^��o8Yr{v�qA��|L�|�*�G��n�s�z�8���������c:��<:$di3�=ӷ��9��}Z	�1�5�a�1W��+d�g��s�X�豞��B��A����e�X�%ч>�x�~���kS��D"�qx�Ձ9��)I���8�\�C����S咭7���W#���V��{ώ�<W��&/6�Q�:��q�bU�I����*�W��� .脕�����Uq�U-���B�S/��f�3��#gy����!�h. ,N) M��n)���ܵQx4�\l�;��Ŗ���x�����ե�%@���4QGѣ�����G����WY�������uĘ-Ѿu�X��GW�쥞~+�W�������[��,:�K��h9G�lH��VG>�uO|�XQ�םǮ�.��衞XP1en��$X�D]��3���Z��T{����vǮi�'.�>���J�����on���p��=e�!��8�O|Qۍ2�k�JFm;�$:��YyO����\=�hp���,�#�x����Y��$�#m�x B�i#q,i7��{�BR��.����{���s�������Ml0#��d�!���U��Ye`,�,p����O�����.'`�s��/�..=�h�K��^NO|ȭ߃��|G�'�������D�{�@���W�=:}i���hs���������c'!]-���,��\U�{�:��9��������bx�4�v*���lCن�J��s�%���%+W����ݏU������O�߯w9V"��!��Μ �'�?��'grB7�-�$�`�q�~s�	�d�E�	젷��Dٱ�(�z~��y+��}Mu�z�=����� U�I~u���#U&T]_?c�3��(���=�νY?��;��g��tS^�X���(�9��A*��xЦ��4ޞ���D�����M��;��:j�<��; `���B.���S���a������t�`��#�
�?'�h�c��Rw��\o��{��ƀ?x'1v��������㘘�h�����˜���9fu~W��M֫�,��B�X��tW���<��#_@S���@ŋ�����k���e�R`b����K�ь�8�Na���AA�bI�yj�̵��yy;��㧧�3?����_����==}�����u�����ޮ��׏;�@�����������~���~�7�~�/}Կ����Y����rtW=ǓN*�t�A���-�<�[ͳWa(��i(0�F�#�k>^�!�g ���ψf�l�G\eܣ��ܑ��!�[G�Q3��x.JJ�fE:i�u��-0H�m��>��������IWuF\��/��O>��>��cà�qv_u���$܋3ǽ�T�s��J� 3�i}��$��^���pZԳ�QO�0�d<����]_,�~�J�삟���yb����'$% d�qa �[7Wg/�7o?����<5:,��U�
�53[g��N�C��Ը��rE�Yyc��@`����b/�r���Q����|f��|r@��B��<�?�����+E�@�����%�+o��מ1|��y��]��o���c����.���Ѵ�'�̷!�O80N���c����d��t2��=s�t��+�8g���=qV��/v/sMT�>:FR����s%�ѣcw:	#)��+C�6�$��,\� �s���p Z8NG�c�P$@����Ϯ'�<�����;�EEv�<������U#�l��N&j���W�gw������͇J�
}y���6�w>�ĚclE���z�-㏬s��vͱ;��:���I/ۺ��ת�wO�����)}��{��>g]�����y޲n�v+��X-�/w8��8Sp�{4��x��v�6x��37\1�l��:��@.�m�U�����Um�!������$�G��w=�+焏�9㙯pf&&��Ľ3���0�8:YU�yL�i��b���&���@�5��d�\�mH�`��A�|y�>xF �~�t/s��6l�<�Eux��Ԁ@ȩb8��t�V��8��^e��;ٽ_g�3��G�G���^��Ћ�'Y!���� ���Sǉ�V�gX�L9���2]Z�{/؃vC��!3]܊��}���IYh�Kb�uu{�����U�:Yw@-I	�
�@1�3 S�/Xpu(��F5@6l��a�S��+�Z����N�+��]��L��x���[C��`�D!�b�f�n��X}��v��WN��?~�g�5!|l�	+�wIӐX���il)��`����F�	M���45��W�d�+���t������%V�%I�\k�soս��]�vu�n����� 	d,K@3j,�,1�%<�bƀ9#$0��`�d1C�<��@�n#@���X�1�p?��֭�����d���"�����s�ܚxg�=��ן+��_DFf�.�5ץ����-Rm���p-_p��0T���Cu��X��BQ�m��և��}�S\�����D,�T�����X�5��;ƻ�U~�{#D�#c�޾�<sD����p�-~�y�7ʋ��fs�dŝ���8�'� ~��QP��`��k�n�|��y��!\?BlyH��_����C���az�t�M�����Z��᪄����n�$2}�-�쾃N�s�$��)�N�=��A�&��xs7��ۡ��If�s���xw��a-N�c���w=����a�_ O��kr�����;�&8��w,�+&�w� ��\�î���.�숰�|a�
��O��#�-����϶Q6
��q��;�t,�Q}:�	bW�m�إ�X��$,��}�tb����g��I��C�����L\���W�5R���b"s��S��z����́�6É�A�����Qy�XL��u��=��Ny�����q{�V&�ݻњ�3̅�}q�v0���=bܬ�ߜg�":d���g[m�7gس�g���r��+2쪈��._n����zc!�w3��y>$���k��g�r
�b��9�����U�1H��n��_�e��e����`��q+�3�S|��&(gS]t��y��&y������qI�q�8�7�v`ĳ�a��O����=��S�y�=k�q]4����̛B �e��*�v���Z�l��߿{/���w���;�?L�SP*�p ��}x�dҜ��c��s�ȧu�ʚ�\�O�4�BJ�w�%"���P9}��4��9�u\[C���"�J����,�	�~�����z�D��H^�ك��M�toj��@W�e[�����7�,�k����w�֯����W~��o���~���;��^�kzM�Gq���}������/�K���?��~�/��n��w�1d(�'v���ւ�Њ�E�N�H�$a�I�9�\���	$qL�����Y��_��X?���UB�H/��z�% �7���zqWy�;�~20V�@JS�`D���Z�	��=���* {͝h$��~��]Q9�z�����*�.�p^f>�aS��p�JF�K�q[���@½\<����V�'�RG~p�����i|�cJa�T:�]%|���[�Ս�`�q��#/R�4G��0L����hȴNN����G�m�3����$z|�lԇu��+NDP'�{��A
c������Z��47w�� ��~�nhhU��(�`����?3��#�%U:����OO��ew9��E��1v��1�h���S'���
��c������v1�7�#���g���w;������(G��N�n�O�}�c|u�o����d�h_�G�����8��������N����x�3��x���S<	�V-�����E`5�Og�prۨ���c�d�otX��-X/~?�%_$nXz�J;�|�:t�x���J=ok!���&z�CϜ��0�;6N�J��]��w*�p/���˳�c�g����͝yj��:u4o��;|E��t�l>݄�UhآC8� 󰸬czx@d��!+���a��2���?S�
��W`����Q�i?����=nPw��#�� j̟��<:޽��`2t���c3֣`���כ�/�Pt�#�|F���b�oA/8�pW2�K ԃ��!���OG���ݏ�ԉ�Ln���㈀瑣�8w	^N�޽���8%�m��g�s��~<^7�����2"����Q�肣P�s|�;tR�"�p�(��*�	�+\T�U���x�a]�����s���+�[�-�m]�,Ӧ�N�}V�_m�cj�f���G:��yU_&d�3�۹[���Ÿ�����X��}!���v�u��b�,pP�x!v��_��!K�a��mȔ���ǻ"#p����	[�Bu��~Sv.���G׀���	���D�%�p6��#��l:ۅ�[��Rۚ��Lp�8\]C#8��8�<�������?���UYx;B_]�L�[�S;, qs~�x�[���D�g���<G��m��� ��/�=ް� ���b�6X�>��<<P�A&2����E��x%�)�ư��|�^6N�;y��==>�"&�!7��m\ʶ�S�{�܌�0���#ׂ���8�,��j[�=a�;y��N#�k���w��/������]��gYv���IFw[ n�/���U�f��&��t�Iw�xe0D~j��!#����Q�F����d9kqO�>�Zӹ��<�]����2k�a���A�h�����Â�^c�H�!��~}�����m�{� �d8TO��4�e;��^qQ��ҽ+�y�@r���`��c"�f+��Ҧ�Iq�f�<`?�܏��fc�� ��u�sp�⊓����C��LG��4�Ͱ��6�F;j�/-x{�1�`(>`��{�o���[��I�c4�\�S92�P�s�g+�<��A�@�.��S����{{:����=/�g�U������u�i��R=��#�	�|h�c�����cQ����g����E������y���`��n�v�gҀ��<��!��l�Զ�>�E�e!`��;�ُ�Ή~Q`�nR$YJ�Q
���ƛxg��t��1-�lR�_��'�����I>�����oKߥ�+=���W���]6L>��6�\�\�S�B�lo���U��HT��^Z�t���Q��jD����7	X	tr�8Y��F�){DpP��5-��a�$mV��A�D-�tl=etz|z��_���}��O����?��5 �5����b�J ��޳�ǳ"����ַ�w�Ə�[_���7��顧��ڻ�� ,���1^(Й`]�m��prF;7� �w�5	�հ�l� �P��F	E��-���"�Z"�'���ω�yu�h�"���2%���?��y�� 6M��^�!�#��S
ٔ��k'0䠿,�m�}�94���6,^����$���Y@4uCBࠪA,v��ר���gC	��  �c������r�0��#�i���a(�\�s�iA�i��P&/^��v��+q�|�#�N���3������1Z�b�����Qy�|�;&����&9�Ji�m'����$�qP9�՜u��p�.8���%y%�C{s�i�O�����%$~O��K0祻�C:A�1>�.�۠w#g\jIa��}A)<�3��Ԛ�鬇�dDgV��{���S^<c��8�>4X�kT_�:�=���I���������	����u�a4����Sc|`@5G��s�H2��Xe<�q���!�99x ~��~����G��2�.kb��~Or�d}����e,�Q�Mn���x@t��O*ٱs��a�`㠘H����Q�x䌠߇��h�qۀ2Zw�lz�žAW|b���s�w�?�079�5�����RZ|�)���i�l���y�f�/B�M0O7P�0��ֽ�BCM�l}��q�HN'A��z��T~2g �%~R�h&���ȸ��&��4o��b9pj�R���]m�/�q>�L �jM��`���q�U�iܣ���_�����⹖ʈW�4~�,�ׄ�l�D��XE��N�c4/�gd墝���ވv�n�Q'��j�S�����C�mQg�X��$�%�e�E�Y�C��D���Tr�6���^?{ǩN��ݬ_���0�}C��a��e�k'm&��ޘ*�ǟO��9�f[I��n&�m�+���8��_Ho)�l�Oe5Lr��# �~�G�|�߁�M��d��Xl�]��E������u���X,�n��lTz �C���j��F���g4�������qb/��sA�R�`���& "�wSs�(ۼ�Pn÷�|����w">掗�i=� �mXp��v��h��z~�>X�4��>�t���M*o�0�G
v�q�9d2R�<��A�*��fӻg�vR��?`&ˇy7h��']��z���9�:�u]-u,ꇍ��k��B-����)G��.6�'�v/�EN�Xpd�Oآ��oZ��6�x ���Q��ĤQB�]������S�	�[�;���4;l���Ղi1��o�H��D=a�t�t���;P�7�!�W�8i�՝�)]T׍B:�\�
���N:�N�9�)�$1ق��c"�>�����'o&Rl�9�4�0F��_NI9�Ya:	��D�:؇%���?��f�O�~� �N:C��Nr�׌D��sF����ط@�G�|6�o��N;Ɂ�i����
 m��N�3����:��\���n��%�3Ɩ�L}0c���H��8�R��ۀ |>�6x�iVA���33F�6���݅5ƴg�P���<��<'�%������^�����}��.O$6hXt�Ҍ�ש�9%)ttz�/���l�dل�/�^���I6uC|�	t{��7��q:��ʐ����N1�.���B�z�O�1�]�Vt���{���8�i`�.o���g��w��'���{���g�rB����5�����<�(N �[�ǟ���_��Ѿ�Vo8��'#��K|�$����  �hYq#��㵞  �%;��+��*w۲񅀅P�=�%P.b�\IAl�@�X;��1�Z�;�P�5�;��+��C�-y�я���L��5~��?�^�.��\boP��ן��#� ρ��ݝ$b��ˢE R�����	��` ��_�xq�ꋢv'��(�;va���z�o�nr�z���xD����}�,GY�9QM��]���&χ."t�D[;-\$Ҁ�|_�k8"7�H<��-�Y��4э�$�I�R�ôI!;!c����
(3J�Kp���|T����n+��]�28 ��]^�r���Ａ��^��:_��sՃ�z�%�G�lo1$��X��
㟏�'�H�K�U��6��w��iN7�h�#&^�/�y��:šK9�!9Z�=2��"��4�3��y�}�o/g�xˏ��K8�����DwAv���B�AP��bK�@ea8R�H3Iv���C���6�uK.a��F;H�lAr��tǂ����K���1�A}Q��*G���;��U$?�n�&�vb'/��ug�����WBD%��y0+�|k,��"C[s_R��i+D������fHr{4����#��o��Ew9ɻYnv�.��D�=n˼�m����7�9 ��%ƃ ��s��.�(;Q��0p�"��߃�p|�hv�F���63.���\�����X�e�����Z:p���ι�c�s�o�A�B㯌U���F�,� ������x����f~�6���u�%С�#��R�l��3��=��u[�O�U�$���t��x��]�����m1���7��8hr��{��E�BGU=\Z+:�����v)�|7�s����$�I�mAM��2��1V�3A�38�7��*�:����i��B%%ˠ�<5y��b���Bևs:��e���2C���b=��h���߰���h�C7Afh@p`^/��&���L���渚�LԱ��:
��?DC\ѣ}����N8��Г�N^K�&��}:��-:��M`ڰ���#)F�w�EC�/��xn����?L&�|�y�O�t�-�;�׵�Y6�\݃7m4�.�k�[	���D�z�;/���Y�[�u�'Pe���:��U�a�S�,�K�C�|C �-�\T���~�E�P=������ߛս�3��)o2�����}��=�\����$t���ڐ�"^��	 ���>y���Ы,��u���b~�7q[�ulw�	:�L�:�AWl��Ӭ���ICm*�1x��a�*��w�_���ٮk����}n�`y�E���s�s`�~�}���B�(�,�s�_"($�{�P,;���=�N���f󆰙&�����Qn-�� tR���hz�{�Q7�ra]c��%N�4��dv�Ut_��;�)��3�u�+b�^��^��}K= �o�B^�{3�g��%�k|��<=��?��i{������~�7C����^�k��W ���������/������g��}�kv�fۏ��E�͎��_�N.�>��B@6v�;�
NC?�-v�d�$�HG���q�8rU��}yd<�wD�F[����NƟ/ ��4_�C�����*�Uq��rb��ΉUOM A+� F�Y=e��1/qj�e�En`T�cU���ߙ�Ч���~��<�*+p�;��Ǹ漥���:S`{�z+b�ˤ�����D�z���|����g&e��~�@L�滔���� ��m�.I$Z�Tv~>�hr�/R���2Q�;a�]�4��(����u,�˶�����e]˴�.>9��N�A��b�^.��L���ߙ�p�y;�흖M�n���]n�ep�ŉ9�p߰^���UG�����,�T&�y��ޭ�m�4���z2?�En�Ü����(?�;ʨ�x��K��Nڨ[�}�z�˙b��;���Y�c8�<��^�۫vG�}�V��(�Lt��|}ұ^8��,ud�q��v�{L�L�h_�%y��{�ײb�^3}�ӔhJ��w��c��g���<�ŕ�^�Y��&8��:�����Z�>�=�S5���g�ӱ|��}�ؚ�B�m�X�
;�dǊ�Wtn�KX}�ag%ϋ�WW80��s�W�Sy��Wi�;��Z�����vk�g1��2����qٯ�b~�6��θ�y9�y��p��_i�xf��R~�߸�A��O�X���m���!��m��7d��<�g]��C����y~G�hK�+����}�V1&�m��h�<��{�NŘG�O���;����#1���H����9�u���S"9_���s{]��800sng��
Odlȋ/Z�&|�bեY^�v������Q�5�R=5p݆,���1d���]����>�K����4]a!����Jǚ�l�j�_ۻ�#�����Ιm�%�`��O߿M����Kz?x0�X&cq��*3N О>��M��y+�B������Ϟ��r�y,4�J�D��w�`��oN��]� U�2�S�������>���c�F�s�gܝi��9�O��s�>�[yxN�1Щ3e����|�}�6���
��R�E��3U}5G6�-�1�8v�>��yL��
>����O��U[\�J@���:������j��0CʝA�^h���1�elc�g�2���۽^i��YO�|�'b�>C+U`h�gC�o�+��>y�Q�n���ۻ�w������o�Α ��5���Tҏ���������O��?�g��������?v��8�iK�F0�<�v������^~1�7"DMП���R��nG�ջ��G�4��ڷ��{w�#�仮�p�b�����z��۱q�r8�Q0���?�]�e��;㗆#�S>���u����ŕ{����t0b  <B��tf��VNT�'�K�����;�@]�yo�iA��Q���C{&p� (7F��*������d�����q�`|h��#�ʞ��y]*�ak��\Ji�`L|e2DnԍUY.u�[U��S�{�8ɣĂ��1A�-J{���a`��,���0�%�_4;�n�7��z�$���H�M"���ۈ�e�^�w��aY�Y�7F<CP����{�ўc�cȏ��y�NȞ�Z6z�O��������dˆ���sDu���ĄI�v�>�}G���~13t��mv�0�0"No���hpSG^��s����D�C����9�n�*g���(2.t��(=vDs����oZ�ع��F���>�y��u�5�W��p�nm
��㇖h�9��Ϛ\������<l}���.�o7ҏ��QY�&��l~xH�m'!��oֵ.��!ޅ�˄�ְ�A���T�R̲����ϸ�	=�H���)�ƤZ���+p��t �
>ay�j�ǻ�K���w�E�Ϸ���X,�N�Î����jM8�V�]�֝�WMrg˔�R��*sg�I��>=���9耓|�1���竅���v�W4=��y���ǖJ�;�]PA�DW.��ͭ8u�"���+^Y���R�@�yb��.�)�&�!ˠf2���"����%�m���S�G�'.����}A�a̳,Xڡ�8��;���@�}6�8
W�p�2;>0F��M�7�r:����=�����1乒�{�S�V��iW���^��[�E�4����`��»R�Oo�-��59f�����idߢ'��6S�'h�F� �<����+~��g8a)����
�7���-��#���k!b�7uG
���<�<^��A;�]��p�iJ����T� ӘD���۩�v�s�Qr�� N7G�cA���Qꩍ[����N��ze�C\�ac8��.t���vC&q�9  �u�)���>�a�3niK�Gf��:�籰���1�H�|fE#�#r�d�3s���׭�Q�tֿ�'ƪ�u�oD�����]�/xvazM��t�-�X���ۨ�:`��ͪC�'_f@g�'�i�����<������V��G�v��Q[El��'�	��WR�T�Y��_��>^�t�i�>�9ۉ�
MϿ9 7�;���iv����Mn������y|���si�b�-����#�#ȍSx�b�&��umt_�Q��}k��;+� �]F�cz׈F�?��+.�� ���C�+AG�&�E[���~��Ե����w�[�ο�;��?�o��O~��?y��FN��og7�kzM����U ���q|�O��?���~��O!_|��Y�=�8m�c�e��J
(�,h�SRx(�����sVDP��R����Iy׊fF#�)��;{�'���Yh�{[v���q*�*�5���V�be�%�ˋfGR��W~�Eh}+x0����� ���g �K�<��V1#Fz�#� Yw,��3x'��Q��p*���z�r�B���6����_�79ʻ����Nd������F% P�6>���x��tO1љAz**�O����ot<��k�V���Ǵ;�悳Hʣ���ӽ�J��F���P:ir��#�Xﾰl�������x��p(蛳���|,�����X���Y�,ީLn��M�#��
�9�oH��y�����q�����!��R�/݈���d���#�q/,[�<� ���'��q�E���	�_�C>ņ^�NçF��Ya�M�����.u���k���{}��⣇�k<���p��g����ҊC��b�9����me^D�a(-^h�3�$(ArLK�])�
3�1���hx��LI{~���Ŗԣ<֕��&�(�cU��Wp۴I�Y7���}1/�(����h�i��K�����,]��1�3����~̸t`0�s�K:��� �~7�c�c��X6tA0c����i�㴻9�}�4��Đ'I&�"iA#�'�����j(�U�6����r���'��Hc���a �����EZr�q��K�F�6�k!o\(��;�V�8.����Y�1����.��ː��p��s`��N�z����$����e�$=I�<Z�/S�$�)0�����}./��4�L�I��� �"�i�܍��L_����q	VS�F��Y�a���%�_8zwԹ�;�uM#c}����c���>Uf��VRz�A�2[͛���C�������amIs�lr�ϥ:O�t��#c���pJ�ҤS}a���mu��W����#�����G	��7���ve�4
p~'n�<���;�ʌ��uRB���,~uL����#�q�_Q�:��̕�Q�cWL�T'U�r����n��Z�-��e��]�f��3W���ښ���K�����$�L�z�Ss�=]c�AmW�`iam�<�u��p/V�2:��V�z^k�8~�Z�d��A�]z� �na�̶�8shi0<�T�>m�1��:�#��@����Oe�Jr����~�ѩ�*7~c����A�|4�@�?�56�x�hK�g���>jq�fS��4�bg��@�5�B�j���t
nNc�Ґ�ʍr�
��1��.o�/?%��'��"|��� �i���D 2p������?ͧ��x��</=�y^F���r�ߛ7F�C,kэf�������`���6�r9�D�w��|���V��t�PSF�
n�k`���ذ��F����_�63E�B����`x����/�O����t.�
�M�7�!��x?��Υ�Ono޽��7����?������O�O�����7��kzM��5�I_y ����>����������ǇۏO�7�ӓ�ʪ�w��}�`;^5���^*𤨠L �S3�2�zw4׹�o<J��� ي�q$�߳C> ޛ��d���ij������k3Xo�y����tU.=���RG�cW���a܁EC��^���(V�g�����@����Az����I�0:Lw�Z��/x�:��<I)�y��� xe��4z���1?��ǲ�ښ�ceH6n�����~߷lLa>�&N���f��X��`�z��g��^�W)(m)�	�]j�/�W���X ��jlr�Sy㱗4OP �૎��2��:��Ng'>��,���h���b/m�����<E��v1��=�c^4�6�/A�Xf�St|<��1��\��������N��K�˗��m|*��-��n{�ͭ]�a��j,���M�1�a�GO�WY�Sw����$v�;�{�ӵ�+�� ��z���!��:fK�=��-2���� 0W�O��d1�0~�"�g-�����e":�,�o7>Z��I̞��z��p{��U#M��|>xa�/���?�zV���7�y� V�h��is]��+fY�<�{rF�$?ߥݦ<E��/-��n��;�P���?$�M�qܷf��D�ub�������E��	�fs���k�*�8����đ���u,x��#��RCOb�*��b!>*m�:iC�+ �~�g��뺣6���/���ި�^�f���y^��W�jٗ��������}{-���k>�ק��~��W�[���$dS�ԯUe&��ޯ�͸�9�Eݲ�CZ��^r���8�0�x���C�͜��z���S��M�E��9tُ5�`�g�mA�y��9|�X��r�i����gx?pL����z�}ƺ1vܟ�p��>�%���e61_5�����2U��a�GJ��"V�4�_�I��������kЍ�DȪ�����~	�X����a��K�E�DE�W�O�$��4�R���>�&ٞdG<�;�`_$ez��=��7K�xئ/qI?�IsT��H�nʛ���x'+���\�Iһ��B��Q�j�Z8yI�e)TQN�v��{̏-��El��}�Mv���_iѥ_��왟���,� ��׹Zp��\栀��tmK�����"���kl������5�qj�;�n���漓�3���K2�d�����Ǻ����$ls]�����)�5���X�� Z_��}�K������؄�t��f,��{��i�s��[���o�sk_��㷾��~����#?��s���kzM��5�I_� ����_���۶�y�\�����tG��l��	M��5y(Z�E45@�͆(�!�q �h�sAz|�p7�)���ppl�|�Vt�سap@љf8?��B`��C�}�������������~���9�(R��Ӫ�5`;������x7��n������ �������nއ��f@�Yaـ�<��J�\�Fa�[!����5��~f^����l 2���6���/�vi)_M�řڇ0��[*'����\N�s@��6�_/t��Ҙ��y�m�ct�� 
1&�}no��c�N"ʞˈ1��mc�P�}�s���ݿ�4E��}����Nl�;�����1^���z����i�@C,���r/����٨����9��g�t��k]���������g�c��a����i9��� 	��|}5�Qg�Qȭچm�{c��wr��7]Č�>䄳��P�eI���������`��j	��a]d�U�_��H;*�̹�񙯓�޷�y�C㶭�?�E6��y���W}� mE�d۽9�ڒ�Yw�zu��:v�q0S`�����x�d��I��{yWS�{��^����>2� ���-�������Uy�PW�z��J���g٪}���2��~@�~�Ty!�Oȸ�ʶ����7��q�y�c犵���[��M�gгے��{��#�I��U��]���"�|�w���,��rvՎ1b��5�]��	݂gk��K1�n0}��,C%ZhT��r��X~+��O��s�x5_X�s'�(���Y�B�w�G]m��u�~���yp��g�gv�s�KL=�&�"5�,��<��=_5-[�O�h�_�U�X;.����We�裶�.4�ΰcs۪]y|0G��Z�>/8_���w�%?^�N/��ֽ/���}�2��J��ܾ�N���}K�չ�M-�g�]�1�ՌO�tm+e�/��\���y�������������'��͓��1����?q^�Gz��,[����ʈ@*I�s�������Y�hNf|���K/3
׷F��<�U���js�S����L����ɲ6xf5ߘfx7�'�l�'<�\s4�{Y^���kK�el�C�u�t��$�˺��n�l�T_C��5`��%�a�̳��'�n���ڏ��	��xa.�O4K�f�h�	�<�h����������0<<<�)-~�e��%c^���eW���.2��G���9pn��QOf`�ו��C�8��zi05�����x��u	��㢳��jW6'������:h��q�X�*$N_�mM�E�_5�����y5��������7�۷�7�����BM��5����� ���O?���~�'��o��?������T?�
`V�8Ϋ�Rb�%S�T9�A� ��~O/�;Rc̼�m��N��7W���罺8^�y��fQb���@@�v��� +Qgv�������@��C�̋�-06� o�Eo���1�C����Lk�-���[(�B�jY�����������ӽ��O�8�FH�wr�г�-��PĽ�1��h�4�F�L� �#Tj<�An���	�R�-"1d.�!vz���~��?���}L�=�����?�5pfG�P�y^ah��ك�e�l�ü�}�'3�A���'"�D��Gf~�xl�E�\V6��8�t��M�_�>�#��,hL3cm�4��Ȫr'�-��������gO������/���8�qD�o����^��o�w�ǺOl�E�]b�XfMu ln\���^��s�t�"��<o��.x#ޭr-�7;�S?%��[�S8X΄,���?y���t;hѲZ�!�c+��O�	�t���^h+؅��J�4��Du��Z��z����!��'�̭��Y�2�H�h�ө,[�N|:��1u�N���K��m�<ď�fx@���\�8��I?A�*O2��ηF��0�8ޱ臗�8��t;�Y�M�	��{�'�{������8�*��?K�v�`�����j���"���@�{���9� é���ч���� �צj��;\F	�������1�-��ݐ!J��2�)�gϺ`I&�c�W�����mو�����r,�Ļ��+��|w�o[*#l��9(�y�L\�c�֗'\��}�m&BD_�Y����{ƀ���t�a;^�y�p�{����<�߹+N��!�J"Ḥ_��
u�g���6�=��A���㻆'�RG�F��v���l_նU�)S4�j����%���+��ٌMLG��6G��-��|�z��D_�H���L��<���&�9J�֮Ă��eA�5͋a�v��`S�-��:��ຢo'Mn��H��z%�y���7�S�/�iП����q1v[�3��ƧS�%�}�nB\��M��e�?5� 0t����r���L���/}&ޕ�s1����z�}_�E�C�򘓬^k8���N�g�5�J��%���O��xN��G�<��(����������7������]I��(�!��}��:y�Vǖ�w���Ƃ:�M,�տ�k�����|?Z/퉱
��6�Q�G'A�K��d�=?�*�esD��W4�����#�%ڀ����/��:Un&;Z3,Ŀr�k��^��H�?/����`j��az��_��4����T��Y(棏�Z>ؠ��Ř9�ξfȫ�l��`YT�X�<�3?ײ"`mQ�zb��Ͻ��F�i��U�̦��D�s���y�m�*KΫ����5�Ć��]ъ��v��
ބ];�c�Ij�G�4�ag�M���um�y��i��#iOO���v�����?����=��\"����^�kB�� ����~�G��_���7����������o��z�[s�f�L�''QDEVY�ađs��-[K��X�p���v��83M��@P&P���Ѫm��oX�&��B|���]�9�Y���9���6����R8wn㎢3R��Yi��<I���y�m�N>I�'@�+�e�k���rH�θl�F[`̱Q�q[%v8�������}����/��F��O�����k2�ͧ���'�d�Rak9�����T��$�oX�eߣKK�?�k3-����\���7��l��:� 4��S^��m�ِ��y����7�y���gC��,	1�x�׹u)/�\����i���+ٜ����j�H��]}����%N�'&Gwz�iލ�2xJ��2�eB/s\.�A�{�(��A����ؠŘ�A�۔�h���画�:�k���.�Fy�r�h�O�j<���w.c=v�Y`|f�O(�!�s���	��
z���y������sWH.���w�FuԶG�л�R3 �dK�N$�:����o�#e�@����$�$چ9�(���P��=��!i�+?4՝ҵ\Mk<�/�]��C�����j<W�y�_�)&[�U��ߦ<��-�4!Y^�~��2�����|A���\7��v�2w���!�U�1ɋC:N�"�C� ʹ�y�¸�&�����V��phb��}_�r�D�������Ym��m^�����+}�|� 9k��a:��i�c�������sYQF���g��w%c�͖��s�v��:�9,�w��:��5���Kc9"������)���6�������������7^n��^^�s]��syu	���ߪ��T}+�eC�~���wD��������:߃��dĵL�������S�gZU>��obYa��ȵ����K�9P20h�����\�c�cѮ���+�|E[~��k��9( �\��>�@�U���s�[�[��!��3�b)�-�-��x�8ƪb��vr��7ĳ�D"D���|}O?(m�t���Z�긮�Z����Q�.ȼ�i�$-�bN�.�w�J�����.1����pz����mk�"뚪wn�89Ww���o߾�q9�W����(�[�Q�T�T��ԂJ���� 8��,s��'Uy�H'^)6�J���4�1v-5�2�+޷Ӌ�Z����5 ��!v�޲�C�G�]Cmy��hށc}�{9��>ٿq��O���_��������3�<ʇW�^�k�;6}� �z���g��C�/�����g���?!?�n��Mgdչ�}8-F�*��� �YU��݊��j�eC�?�0f�����!+��$��p�5�L$����v�T�菕����Z@+wI{ߐ��K`�s �?+�?m ?��fC�Jkm���]>���P��ܝp��o�Sd��� Kd�i�u�x���(n��\y��G{ֿ��g�:��3��,���}�4�<��y'V��Y�S����̆q���F�m[���Y;������������Z��n�����à�1�;P^��ɊaN=����ﵬx���l�ֹ�����|�j�F��B{vz��������黚c�)�v���~���|�yt��	��Zw���r��W�w5�>d��n�	�hT�������N=�K����8��Sy�0�rFY<��,綮�e�!�<��OpL_-���I��,K�����$�ќX���a��)9U����c3s����n�ږ�<����^��?�;�w�`�e�s�ׁyr�U�T��a'\u~gz��_NW��"���:�_�'k]�[t�����J7ㄬ|��;�o��|��ĢB�y�͜�P/��ۜ��:߭<���X!N~	956�kW}^���q�Q3�?�P�]}�L���҇R�E{+]�-������:��o�ѿ�3�:9k��V��ܧ��}�����.x	���1/�e��>P�ޯc�S�_W:(�b��y���;tC��x+��X����|'/�"�˸�ک+��.{~c�?+~��u޷î���m�KVXr.'���շ�e�)��6����OWr��{_�^�ϯ�H����wy��`nn�l�V���"c�c�M�!q��U�GN��sֽ5/R��u��d��vʞ��D3ֺ��+���2��r�}���?�$��c�o�9�����>�֝3&Z5��G����^�2S)����uJ�~�=?��Iu�o�x7�}_��?l�p�� �F��F>�\���Pl�[ɼy�F>����XZ�s�o�)�d�":+�c�OԺ�oj�����*B��<���� ȶ�ˆ{�F5�T�o*���Ni�~|2^\ij��ǡ�@*���k�"(a��C����<�������_�����'_��Ͷ}��O�� �����^H_� ��xxx���o?��?�O�s��������������6ξ?���a�1��>g#%�NNf ���G�0z��z�Zrt�"'��#bv+a�(�X��i��ǽ42$в�p�3�>���V	���$����܇�W����8�	G��' |�����_��ƫ���P�9��m�2�o�δ�и��C����<�D�s�2�� |m\�{�|�B���ٗ�v�V:j�M'f>�n��k�Ι⸴����1���*���_�5�I^} د��weX�S�{�m���<�6��l�c|t��q6�QO_|_�/��G�wF�q�]�j^X���X��)����6�H;�sv���h�OR�BJ*'��<V5�K�9+�>�ij�B.q9�$���%.ÐG»ܓy��w�6���iyQm�|�b�^~��(n~���L7�Ou���$�Hg
��w3�3�^����W��}�yf͙x�軵� ƞ~��V������o��^c���Z�JϾ�^j��b��|����j�Ks��~��Ѷ^����!���Ze8/��T^u�ּ+�}��U7}�~F�Z_�v�uZ�hnK=-��}We����ZN-+Ӌ�cO�����=~���V�RNw��}�~}h�1�����
`���3�����Jέ�"�տY�f�m�v�T;�z!�jܯ��4��ɒ�<�{��2hUϽ��NX�{����<z"�l)@�y�1H��Ҍm���+�Cp�)>��|�z�:�e�j��xN�N����(;�!�9�_d�^���v���,k�f����oek���8�c��>3�6\�<�M>F:Ł_e�|���E�-��s�m��g�_��U�qް��>.�N����uk>�ٱ]O������.���3Z���1��K��C�޺[~���y�V=�s��|Ϳq[�}F}Q/�c��f�1�0������˭�[�+;�*����h�����Km���SM�/��P�';���t�m�x����Fb�	y�Մ~����<c���ܧ��6�7k|ZB��0V�k�짲>������$�w���^�x����6]�ȯ�j�s�F�����z��YX�7���7����S��O���������O� �^�kz!}� �B��B����}�����ӏ~��۷�����ۛ��2�Nc�O.a���x�i6;���.C1�B���y*�����ݡ�������îHNSIPK�CH��IN5�ڵ0�� 
�[6�2�_;`D8�� "��$'�끋Ŧ���<~��G�����r{�@Y���!�}���Q���v��/�a���}[�f'��~��Y���#��W���>k�3=��҈@�wH���+��/��S�����x߲q��7�r��ˀve�V��|*�|d�l���
3���Ҫ��?�
����+'�U�\շ�y}�ɊǸO�f������ر|E�u��1�2�}�"����>�1�y.�I���2�J��ׇ�>e������j� ��ܯ�Ͽ$GBo��p��ƺ�v%�8q�X�W}vWn��͝.Ա֍�g�H����yE��$s�%�WuA���9V�M͟��`8�Yr���w}����n�w�м�m�}C�kq�$��{5�e��/���?��y��ϗ��<�⇐�Q=)A�����}��/of\��K�3���W:��X������+=~%gW�z���GүS�3_�It�;�_W���K��w8®e��m��GD>�����Am`�}I�A;�K?��>\��QeY�c�}a0����} ܽ�_�b�,gц�\��g�}�׹��f�;���Ċv+zsٵ�|*
�\m�J/T]�M*�V�{I��v�p�J�Ҫ�/�<�3��_�o=>���_Gɛi��;y��?���
ǆ,]��..�Ӑ������G�Gy���r�}���s>�e��_�?y�[w�g��\���f��!�`-������Vٶ��+Y�i�U6b|�p�L���R�x�@/�4�婾�O��u�5��x+^��+�ڻ��g����=�wM.e�{�n��QN��~�^/�2�!<��:&�7�Rɼ���A�]�^�X�ת��eޗ�mk�����=��J���k{t��*�<��Z�h��ά��ʂl/��θ�1���G�l���/����t��)�-�3d�6��=���	 1ך���R|��qY��������28t�~���ڌ
q�9�C�	�;����vg���c3Yތ_v�a�6d�5G��W]\f�}9�'1�U��t���fy�﹬�o?����x���?��}��<���^�������^Ӌ�Gq�H����/���s��/�w�<�C����q-ϔ# ,+^,o;���l�1�l�;V�.-�~������fJ�;Sd�A�жvYK]:�vǙ�����b����0��Y ~�����(����8+� �=_�Y���;�����0 �gE=�(���G��m��ܦ\GD�����f�Dm�
�����?��\ӹ�����F/��ۻv8��� ��a�Z'��+���W���f�~݄O�Q�f�$u�s"���y��zL%K�{��~��N�m�g8ҫ!u���Ժ����Y4�3ʢkC孜��Qۙ�!�y慞
��q�h7d!���dTώ���p4�<c~s7�d%��F<�Ey���^�a��.j|�<5�á�'�@N�n��r��Q�i�{u"a9;�V��Rz��0����6��1�j{Bw^�?���{p�J_0׻�g�."����<E��@R�ږ��s��[/���~>�pZ��\�	���� ����8���g�����1�:��W/J�m��?t],Ng����u^��kgҗI!'П��ո�~�[�,#Zz'���:��/xc�3�!-#��Zf_/d�tp���jV��\8}g��^�mQ�~��;�6����Bo�isb�����ژ�jy�o���э��v��N���g�}
>��w�Ń$[�v%m��0���0|�G/����m�Rn��1n�$���sq�<�t�6a�J��6�9��9m�::�c21[;dtG�6G6Z�Z����%~�3��S�X�:|.#�]�zs�,ϲ<����;�����Y�]� ��j�F�g�K��,�����W<U�_�m^��	���j��y�6�-�'te�v���2B�e[�I�Ϗ�^�q<k�>#Ɩ�.�
,������tဠ7��2FiyKma^�ҫsjzڦ������|�=�(�d��ʊ����y���O��b�e�f��ݠ�6�ԋ$n��o<�x �pG��zsC��>�kͳ����g���3�yC���[����:���	�"��=��u_��:Y��<�^j���/�tY��ys��G3�l��Y�0����=�=~[��h�y�q���N����&�s��b������K��}�Ϩ��}�ù������g�#�}jx����<�{q�H��+�ʏ2�]�vx�S��{�ك$SI_˼�������ð�����a�Q��|���l5w��L�����-�<Ӻ�S��|�߆/P�$�y*�!����'?���[o�����V��kzM��5���� �n�D�}���_��w~��K�g�7?����o=<��c��`���R>NPzl v���*lI�u�����E�%����x.\�msEv�kuhj͍ܬ�QfD��	�I�"�޽T�Fi([������塞ږ(�(�ϑ�ݔ�3k��y�  �[9��)+�+�W���Κ����s�+z�x8Z�F���yq��\��m�� ��tZ���G X�H�S��G6^y�����R�3�S�F��NP9�;5߅x�{�K��a, ����m��&9�$d�p�=�ۊƱ@}�{�5�}i�4qd��G���S�' �܏���{�Q��J뻄l��(��-�эz�2�,ꔏ�(��,9�l8�D����<v��:G����l<����m�	�o��R.�E����'�A0�_���F3�i�
ȩ�s�=,���<��f�Q����o�	Bӄd��%������Xa���4g3�8�Q/%Ǧ7���c`	o�c�����D����|'�.;���2�i6�N��P�c���ȃ'B��y\\��/��c�F�P��K�v�����tU���3/�w�lf��lޭ~��e�e�]bw�O�4��1,�a=9��z�����sџ�8�&N�X9��=�	�̘����+�|$��)8���$qz��4g����]�1_*_>q�Ux�gr�2og��}���J�+�}b�N����{�vl�~� 	�y.� 돕?�9�2r�)�e�ﺏ���+,��ٳ�~��ۃ|�q2H�әg7����ƁC�\���cJ������Ɍ���-2�rc~��RuΨro%��_��z�b�-�J;����pٗ��s;�{{����X���u�	�(�mG`y��� '���bs�g<�m��7��-ߛf���w�����d��j�x3��ԣCFoiN;�������gȆ*{�!?%�څ��%湊�Q.��s]��� =�\w��9��8e�v�����· ��.S1M�������H-��-h�|��1n�ҽ��_�uYN@������d�C�������,O:��z�Xf�,��[��&�\Ws�[�ʙ@�n�o�gZ�-����G@~4��|�v��z�<�qxP��D[W����-�g���,���|��CB���p�n9���Gǜ�T��e��t�
�x4�C�D�Y.�?�q��%c�o�l�)_��$��|�ģ9/b>ֻ���q��}fڰn\�\����i&���1��'�r��VA�]�0��Y_���h_�� �@[�o7�:���U:�I}u$�|���0~��__����}��w@|ME��1o�Ot�6qF��x��oc�\����\V������('��x�1;����k�|mjr������g��w�3�5�7/�����}��8�ؔ��9 �����>>Ŏ�� [����M�97��- E֋��:}H�^�����?�&-��y�<{�f{w��<>�޶�諷�ѥ��5���4��	 �������_�~����������i{������4�M�����X8v��_V�8��#"p4ɌAu�G�7r�Ù�`MۄŇ�L3���`�h  �9��B^D���:�����+V�J�W|fe���J8�ˎ��K|Οj��v�N9@#�!���*(����������u�\v��q����[tw�a��78��_v0�E��@0�G=T�qOg�8��޵�`f �4�ǳe�j�j��CP�|�ۙ�<:;�5H ���r�XX9��rc���MJ�܈ѾoԖ���m��c<�>͙đݠ��lĤQ�1$���a,�8i_�qh�OQ�Np��H[1��.6�?���c�[$ӏ�y�ڥ|���|rDڿp��w����l\�|8z��8�2}C]�۹m���Y���&�a�v�]u�;���[4���9ߎ�Y6�+p(��"�Z��$����{w� ��8>�����c�Ğ�<o���('dG�2��gS���=/u�}��v���!�l�A&��6']t�t��_=�m�&�Ov;��`�wR�����0��a֩��2�ws�$h|t�Z`�-X�c�>q����3�[�3�/�>Go��㹮hG~�,jK��(�i��n�)6Z:{�;�Ɯٸ���w�l��Ƌ�3ڇ�� ũ��<��,p�Y>߹Ѻ�"~��~���a�]�����k�O�S��2��{�1V'�9��M0���_��q�U?�1?��F���c���K�_�Zp���Ч9p��ԭ�b[tB��«b:�� �.��u�> ��]˝e�s��D[��Z��Ȩ�w.��+ԇ��v�9���H��|ص1vQv���L�w��;��?���������3H	�w�4�?�?����x��О�p&����w'5dV�E�F�It���β�f��B���Wԉ�K�tЍ�֠��tW;to��Ȳ2���1�0��X��	}�v�T��6�az�$�A��ef��J�Yמe�q,0��.��zx��s��)�-�w�v����|���1��ݞ���A �8a��Q	�Z­Qdc��4��=�x�ǭ�f": ���jr�c!�h��z��M2�F�y yg|�m��Kd}�	Xd��T[(�Ŵ-���9�El`0����_���B��-�;�^�B1��Z����*�M~������gT��Ngr���[���6Ě`;_h�17-���o��>�� �c,{��v�Z�,2�CX�m:^��>�l�Z��)_:����Gt�n�x��)4WD�E]��϶���g}��ce�b�AE�'ԂY{����-0�H��l��=Nl�j`x�!?�Ե���٢�810���	6L�Lc�3��r����d�T�B�u�㧜p��Fz94n	�r>��<�ޓ�{6�KvM��_l[
�e"~������m����e�>�b<H�_c�>l1���Dy
�qj=P;vo��A�K��g��N��v!���!�aПF��~݌�����ħ���}üf	�NN�R��x�붜.9g���B:�����M\P�Z�l�,0�E�P�ٮ�Dz��gd���������Kz���2��y���n8 �e�;�xs�'~��w�%��ǩ�7zt�Y;���]�������o�k���Ə������O��O�z�kzM��N�� �f��8>�o����>{x�sOG���>������g��w�B�ǫ׻�;�(Z�
 Sn��������E�h�f$�xժ�C��Cf��w�`�kh�0b�W;jĒ��\��^���l0���NmR:�9TOZ�. �s�}]nurPW�`t�W,��(ᨫ��6��岹̙��'5N��N�3#��3��[��E=l� �mg�w��C�B��H��|p�B�3���g�|<6�A(_��l��� wײ#�'^��]*�\��} =�SG�fg�����B�%���~D+3�>����9j|;�_.�v��W�U��		�� �� }V�� �:ʓ��(s�XU�0m2M���&uq�N%D�r�����P��R�[������ ���LN������.���X
�̽�A��=���UP��j��9٨M��$����e����kiP���+ȷZs�z�0b����@y8R�ж2�Ǣ�;#:s���9�����h��nۛ;�G� ���17��$m��K�r��a׹~(��ݲ��5�B�G�X0�S"(��2�w7��|tg���A���-�B�3/�m�s}o,^&���B�F;w�:mF`TuE��9hXk���B��~�ȸ� /�Iˎ�� g��f����l�<PB�Z�u��6�9z��k����?���(�)1hg=�ðw��́�H�A{V��񌣜�`\���g�v`��&�Pe�i��a�;�VoO7�+~ڄ����N���oG���y�<��;-@�s&��;�2��yE���m��J,�o��&I���2%�"�- �X�+̮��0'��F��_F�A9�~`lue[p[�m��OIe���y���X2�U��h��I����#_\=XV��#x3�~���iј��~�����\�w��M�;	���F�*��6,$R���уGmp#����\��`�Gγ����?u��3M8�WG���8F�"v�o�s���t����d9��/�YX��q����/��.�ⲣ+�½�]\���QY^a��Ǎ���s�>��T��m�Ghc�ұߧ|cjxg��6���ܮ'2�}�ysb�8���r����~����,�u�a��6���|�ң��X��;���� r�,�\,�����;7��L����p�@N�Q�w�]�9�aS��Ð�Zd��N�e���觮Ep"�Q�F��1�	�B��f{OvLj�H,��Oy5� �y�h6n�a����5��^`�A&�������)>9�%�S���b�kG`�Q#�"���R���F��bm�T����t�6�w3�8�<Զ�4�����֨�����������.��*�Vus{Y�FP^Љu4�� �!�ƾ;��>�z���~����8��t^��G<�|I�<4_*�b�x@9σ�7��j(�{2NO��7���&d����B��=�#>�v��n����4�%���ls��O'�>�nc��� �'v� J��1g��������.�$D�nC��;�X+��z�?QHf��/8�,e�	��u{�1���M������f��iSi_ۭ	�G�n���>�;�7h��G�7�_øN!6lm��c�4J>�T��|:Nk��D��F�r��:U�V��i�?z~�������������������������駟�xM��5��e��� �+��x�[�?�fkǏ�����<��� ������8^˜�-�<�&Q��S'�)��Pe��hh'3��ȗ���!�
̬=C������ˢ#�����>�ɳ�]a�M��r<�x��I��
��o���"򄆨�:��@b�����"���0�8��>����#O�u=  Ss%�~�������|_$�{^�
��\18���(& ך��9\?�k�_D�������e�]e�(E�NQ���Wj5ࡎ�x%�o��ϰ�?�i��Ӱ���s ƚ@���s��X���k����@E���1x ���������i��0����HLg���v;��C��f�ka�M�� �f�	����d,5�c:U8�9-���v�';b��j���Ԝ�cg;�^���"⎝Q��ϻ���mA~*�1#��'����18�r���QݔO�3���� {�}�{�iclq�c�~}�ۑ�ZU�08��r�Ǯ���?�������Ŧ�ff���X��`���S�Zo�$4��v3g���ѝz� nm�i7��/pt[H±�cXb����j�6�(ࡻ,��>�������s�ˢ\�	��6�s��"	c�;�gAeQ�e!I̽fs�v�B;tR�3�h$��=���� �4ݰ{�ưVu��~8hԻI��X�q�x���o#�ě=-0⚄}�bͦ'4�1���ֿ5�e{sml�@����G+CN6>�;;��Y_|�Y�(��{�]��sqb���Ce*�1�N�X4g���3f���bZ�=�%�p�� 	�����=@r�Yv��X�B�o��;�#<Ș$����6ϗ����C6&cl�ʮx�9��حOtu�:DL�lD�滔-��H��V��\� �N��_�+
Q���'�!��v�[,�~N�bB�?�ꘋ������7����YF�A��wv����1���0������S��1�Z�a r����;��U���������X,߂�\����<&��GP��iSy�)�����߁@GE{�}̠%�+����c,]�D>�Y'A�T�F���ܚ ��v��;�a��&4'�y��H{��ݙ���o�p���>QZ�)>7�`������g��U��O`'zv4��N�kt���:���p��g�c<�N��o�fq���'���.dQ7ق@K��FG�y��;���a�p��Oj_s�F����~�v4���L��i�flZ��8ч���C'+6�;��#α�1N�8�9�yA�ȭ�|���gO۽/*�����p=���ݐ�@!=�/Y�Yۍo�(s����A��-tI��0_;�TO�Q�������ރg��.�Ӻ�_�l3
�����f㑟����Cq�8O�`��w�įm�/D�3��i!�����g�CG�Z\���xv`K§�]Z�;�羬=�n�Jnݱ����60Uȟ8e��}�M0�h;���튲b��=�i��]��zt>��u����tGs��'��ڍ�m4�k��q$���e�O�AQ�.bmF�/�q:��t5|q7�al�l"�A�*ei^8�;�	^�8]������!g�q[�A⵳�����w;��!��*�=�y�㠺(��wl8�|8���oT0ڥ�~�E�����:�uA\)��!@���B�h��A�s�0^�m/��c�	����?>g�1��T���z�8V=�i�F=;�V��`�1]_���Pv�R��S��`V� �1�8-��>�IF'0|ȇ@�*o]n3VcZ9f��KC�ޞ��~8j�����>y�~������Ǐ�?����������^�2�(N h���m{8�������F�c��v
՝"*���Q�l�؆�%viy�`g��K�;���^	�Ch�1�0\D�ܠhf|����uT�B\P�,Ha���r&ʭ�A�HR��!��9�y�O"���M��+�9@6���g�U��}��� .CR�2�Ց�t6#0;��p= �q���Fi˴�#ɮ��Ê���ь:�l�D�M<>o��q�5�y�+=:ѕ��4^�<ndQ��c�J��ې�2]�Uv���w�(����m~�����V�/�"����orDw%���r�@S��r����2v��,����Q����h�y���e=>�}����$��G&�����T�!�M���s�}�e(5��Bk��F6��Z�=�_���Q�̧y�y�˵��6��|w��@�#��Q��Brv�O��s@�\I�,�j��ϋ�ni��b:dc��)�b��t�4��N3��ce8,�s���Ag�1�w��A��G�9@&JL�~������*�ӌ��JO���-�e�������qJ�+�-�W#0�4q�x���s�!Ȧ�sr�T�b��)N��+_��d&Xv�z6dn� /��|}���&�7Z��Xe�z�
�Φ�9ޟǽ.ϋ���4����@C^f]��ǘo�{�~ϟ�Y�Vu�9�T�����R�Vzeֽ�8]��<V�t[Ͽȣ�2ffy�Y����c��!����:����z�A�E�|b���	�d�S����Q^���S��B_�inG��Ґ�r�"+^�����ۊ�[���j�_��EU_L]҂ym�2��|sx��^�~�3������B�z�eR��M������.�+��*�0�����9֧�7��^�Љ����X������&�QǕOо��L��U�j[���J��{�����T
9�W쩋���)��~�L�U���A|\L��?�����vZd~J�#-tx7=p��/�G��S˜m�+���tiOWx0���K�z8`,�"�����l��T��>�Hl�kߎ�/��oc�([/F�/aS���]����P�t1�J|q��F�B�0x��;�Mm0�6���錩A4��]������i���Md���1�90E����ޚ�^>��ߵ	��>��#��I�t���/-<�}�/{�x��Y��1�hhG0Ƀ^`Go�=����%�]�
�FWF�l9w���7�<V�o�.�����M����Pu^�>�q_�
��롫�m|
C襪/��~�\�e�ԗ�1I��2�ԉ��z8E��S��Zg��9dk�H$_H�e��HYpVO����NɃ��Z��T��8��<f��;o��q�(c�+��zlu�Y��}�	���!+��}�K涒n"�wesIo�6�������M�}$_@�BưZ��F�f:փ���nc�#ط����Ȓ�J�<��ھ���e�<~���v�P�s�������ϝ�s+������^Ӕ�� �!���oݾ����������C�7=����n�#X��|� ��,�)�

����po~�p�Q^8�z��VI�RF,�q�	�JӍ�W;�C^D�`O��Z�E����s����і��+G;F��*�ȑ�����m�v1�ߨ0D$E�&�-s+4���}���J�X`�����Ap�0s@4��e�'<J�%"��1N���mD}��r���`��k��c,�G��z�{�e4Yn�ʈ
�OW��QC�t��e��F�e����Î���09k�Mr�ZE}��l`���~�����H$ù��:O��,R���r���%u0�1w��px޹4��L7a�v�S�Ǯ�p05��Ǒ�G�sn����l<��`:A�G���k�I�+C
���$4�0Ff����4~^�ѥ'>��t�y��U?hҥ��M�s�`>Q�P����Q��{���2�.�{���DC���e�`�p��`�W�<�#!U�;�W���1����潾8���s�m�.B'� ��CPBgyPǹ�����k�:%�N�9����E����X�� �M��L�NNo�cd���ns�;�_1��������tˏXLa��u�p{�Οcd�R�:⿋�Ҟ��9eم9�U��N}�ʋ���+ʛ�{]`ǘf�r���vLef,u��'\���s�E���Y���ǖy+��u	�Lj�ד�yx�k{ſgz�^��UyW)Rh�ߙ?��˹�˚�hw�U�΂�]��˼��i��'׉q�yȿ�'�w[���YnU�y��S��<�wƖ�c!!~��☋�_�q�������f�9wu�2�����T��u�WynݧE��Щ����_�/d<�����G`�#˽:�^J~���.<�:^��嘯����D�p�q�uD2�k�ˣ�>�\�<0�a�o�S��5�;6HO�<�n��I����Aԉ݀38[�^��W��!<Ct�Rb��%����G��J��Y}��I�m��Fv�9!�C_2��
^����=�?�zl�w��P�tF���|q��X��ƠDԉ��������g^���Q͓����#;��&�p����\c��x+N�:�PƇ�8(%�<��t�>	��}�,����&$ǈֈ�!�ѓ�,k2�Qc@$�3 �T{�ix�4��~¡�$��g��ͼ 9���(W02����$���t�2~�1������z�ꊠCȋNl>�dflm�|����e�qM'?n�%.��&8��3J�GI�[����η*'�m���o�of�	^+���~��^�綮p���/��f"�Os:�?���~�a6�;]�a��12h蟩W����kFQ>N�qt��$�o��B�U�9~#c�q���1���9�?�~���hO��_��?�����������}W�qϙ��^�kzM?�+ ����?����_���_������������vK҂j�ϻwO�a��0����	
D= �p�_e���1<����cFQ!���8?z�{fw�������^UW]Wպ�o�G�ݽ��y���׏Z����U���_�Ƨ��x>�<���˘��uLiv]�׷j��^qb���G f (�����X>��������ޙ��@Rv��a�D9���kD��Q��h��\��u���HĻ�:t���F��� L�����Z�fߎe���@�� ��EU}�d��**`u�_[x�S5`*��#l�@X�U�_ 	�v��l�Aý�͟�(�ꨞ�n��cP�z�A=��)�h�r �\0&��Qw.ƶ3�v^�{T��{��=>�y���y�t��o�[��/f� ��b`����1�ȿ��;'H��ʪ����L��	��s���\�o���h[��]��VF�Yk� �^p
���.�"����zj�x�_���X��|�97>��|�é��A7��E�0�n2�ԅ�J�,ɀ�s%m@���O5��Ƥl�] �.�>��s����W8/�:�s8�,��b�A�Z�ᔧg�����&�2M����@V��>a?���Ps���$hB�F]�Xu,c�T�8S�\��[�Gۥ}p�4���U����{�3ؑ�~��y���7H�_����>i���zO�:\u��r�(?���p�jl��;���N�ύ���r�l��R��K��NrQk��C7��{9z.;����Pe��UW]�}�}��e�a��+�`+������j�|o��c�u�_lʧ+��Ŝ�f��W�c�*��B[5�}P��S������8�����N���Q�z�9bHm_��oel_m�%��m�yD>���ԋc���ʯ���M6���g5`pw<�G�CY�5Ly䎎w�Y�:W�OcЖ�������W����~Ӄ�eANƺf�P~����3C@Q��h��rwQG��=�H�3%]|�#:��;�e�Y^d�D�I����cqԓ�3�ێ G���p�WY|�>=S]��^n�Z�X��sH��5�� ޔ����3[ڥ/�އ��{�U�A0���a������8�3~qw1�7���@}���	��>���Ee���AÒ�a���[���ߨw�k�����_�<�X���(|źF��2�`�&�s��v�T����ù��k?
��M	V1�'5=}�9�w��}�E����w�~�| ���r!���(aިk^$0Z�}�����>h_R�g����֣_ֳc�ܽՇ��-YO"��iø1!�}��S��^��}�/ht�ӓ�x��{�;��g.f���uB~����c�ƧcdV��kj�[ը�Q�Qo�:oC��v����������K��VǪ��r�����}��U�>�6� vY�cO��s7J) Ӈ�������<��
����DQ�'�t:�L�yz�H�d��ڟ~4 ښG�}��B)x⦵*Ed]����,/ ����'�����>�+��_�ͯ}��[_~���?��� ޮ�������� �|<���?�'��/��?��������Ǟ�c����ɘ8���V��iXS���/��)�F=���Ҭ�:�ޏ/W+��`�Bz�ϻA��gsx����<�[��R�@�)�3�+Џ9�L�.x��	� ���Y�)��A�^�b' �j�~�B���F;���a�~�Pŏ~�s�� f�ӡ@|Q�c�+ώ$ �	�%���V�����tA^(���mn�q�Y��-��*h��y�c*�z����g�}1�nҪ}<�E�+�9� �y��_4�P�������h:��nhq~!}<-."�F3�����ة|N:u:�3a�g�Nέ#�ǘb��a��8���6�4���9�X�b.�Y��:��G¬��O�l�q�2�`:r�$U�9Ѝ�4|F�b�a�a�Ge�'����@O������'΂4�<Σ1K�˘�1�����u�T&���;�a��$��&��  ��IDATI�B1�y��E{β��<_��U�`����9�p>�aT��s�Y_9�9��U��<E�$v����b����9�6h��@��W���i̪��kX ��{5}�;c8�Gs�7��G�`M���lK���'�u/�Vݺ��l1y�:���Mw�՝U�Y�]I���U��/k���Dƪ�`�����|������;����[*��m(7�/!��6����;^�"��vc1�Ӿ�y�u���m�`��X�]��J�rPS��:��ě�w`[{��S�������3#�}w���"�<�e.;¨7�Y�s�� *�P}��w��|�׏w�����Z���5�)ީ���P����AU9�w2����Mu�A1�E^��S������R����U^j��|-s�����B�G�����-�)�Y|���#�Żs�׹�ϡ*kv�ݕ�}��i6��,[iX�tvkbA���,t���Ķ�,;˻�[�=��#pZl�:p�W~O��oQ�P���E��ҥ}�����{�����nU��,|7�adX��"�>�2�m�����y�J��nǨ�9����Qh��z�1@��~a?�0?��R^�g-�p�ޙ�B��`�3��u�Iu�/�1x@�����v30[6(zN���:X�ʽ^�ڱڦ�ֿ�]�h�s�����^&=j`�����H�-;W�J8��gdRRj�xy�uz��T�jVT9�oP~��QWhي	�/��e�vJ���cd]�w���{��v���I?���o�XU��nW&��x�>�s+��5��lX��լq3�/f����X|�2F��#�&�s�S~V���}n�c�`#/�6$/�B��<�r����	�� �Ɋ��K7쁭�{�ߩ��ς�l� ������-둨*��q�Uǎ��� 	���>h��/�fs{^�Z��B�]},�xF��5�����3�Lڈϰ�3�
�6�<?̙cm�P"��)��ޗ�3���zͻ#�zV}�!@��P�]���s��y�r-�J������4p������������r�ʻ�|}��Ƨǧ���}���e x�ޮ��+�j ��6������O���W����3���~�O����G������+��0*��gS�fl��)  �������FQ��}�#T?��0[A꘿��s>s��	e4�,�C��  C��@B!FU�����?��c�c�*��g~����Z>���Z}�b�D����T����j��y���>�� C�3��Ti�_O�|w�`L��z�����g	��0`�,�Sߩ@��n�V�>�;k����i�ՉKc�.�X���g��5��mw�cW�?3m�ѻ�P��}��;oan��{�G>/ػ�J�:&;�^w��h&(U�_���x���t}�y�h�]� QGh�{�ެ���*_���F�@�qv=GGⰜA�d��J���N��{W��@��Gt��Qy����4����
]��8�;���ou!��;5H�H�&��a�}o���N� �:w���}�i ��s�CF��뺳��t:�j�2A-}A]d���X��x�_�Q7t�S�m�:F�f+�w�T:�?]�r�rg� ���W�ܵY���.��.���V=W�8�ɸX֏�c7��*������t�����x���Nj �|�9^^��&�-.f
��|͙�����퓱5f2P}�H�v�{9�������ӭ�]��dfq�n���Y����Ɵ�B��#?���a/�}��>��Ź~�{M?��Y���v�m".���O������n�^���]�*Nq�ZeW��b�y��݅g�����~>�{�a��],<T���ZV�w��:C�������i��S�e�LRe��mϲ��v�*[��6�_}7��\e+֮��z5w��}!�t�wX%}�}�����y�z=�p?�Ͷ�+��/07+t;�f�B�5H��x��QpG�;_�M����ĕ?t�f��m�U�	�KN�[թ����g���9'zP����3��m�d�Gw����ݼ.��]�g����2�W˽�g(3}U������us�J���;�I���;�d�8Kyd�`׳��X��������ץ>'��.�`�:XQM�'>�V�����8W�}®����LlO��n�b���x�U,�S�)I��C�Z�?j�-ڠvˁT�M6�O�&��3����U��(�;f��E�s<�0���׃��1cF;���X��<J�ṵkO��O�f�]n��].�^�q�����XAG��.]<};T7���i�>Wa{{�U�_�w�_c�%
�Ջ:o��6�o�_�CVk{փ��T�O�s*뫬j�*��#-xC0�}��Z�܇���Z��e�҆����M�	��?�|'�O�9#�2��Z���V�l*R_`�r�$�����?�8L^�y"?d3���u�cRY��Q;�n��~���w����Ǿ�����헗�_����?�zou@߮���z���Gq�|����_>��7?H�/ߝ�r�r��33�Q��U�"=OY�X�bs�~�0F�w'���؞	_��HA�
S!ǌ��T������k�ۑ��g؄�0+�;zȭ�U��~t�ڿ�u�����&}�:m�=88j{��v�u�}��
�;X�P�Nc������m��j;�\�nعc�������;�H��W�8X*8�{f���3�axi��p�V�B�D��]L��Y�A�G90:�K�+ޞt���Ǣ����^N�yߟ�:"-#xd�];�3����ye������E��3��|n��������jȒ&<Z`�n�J/�[���\5x�<���.�*ӑ����s��:G�����O2.15�河:eA���3��P�s�yb�Q��n�h�=��]�p�v��7"�	��&Ov��;yyV�F��.f:y� �I�')������H�c�����x7�0K)���n@�1=���� Zt�SPw>����Ӽ��g�_Ή��t�1y��蠼zD�Y]��<�Y���[��đ\t?3]�b8�tλ,�q-.���
�����	����+��։2�R�3Gǥ;�uLz�w�h�v<q��<�0�U
Vw+SW/=��� ̍���_��F�έ!cl�NwNq��=F}S�8"B�w�/}���W���M�e|,\�u�(sE�y�e�_��׿���n٦߹�.|!�>�#����r�}6
?�#IL�u��l�%g��.�L��S��(��Ou{�s:p�c����W���wuy��s�UN�w����5����O��t��=�P}��zAۢt�����t^��;qD�85y;�)�%��.�w����g�݁N�b���uR���U�Y��VL�:�>��y�C2� #�e���ļ]�2�T��f9~ގԌh�h��'�;�+�?�t���3LY�ݾ���1n�"��w̳z��|�i�A�x&�Ő��:V��G�]^��^w x�Z_�Sp��Ӈ_2"�L:�Z�����S��y20Bq�Ĕ2.��ϻ�~ky���S��x2�D��'*8����ڀݯP�a:]Q���^��Y3��r�w�QS�{[��n��̆',|�<���u�������W�_�Pa
>V��W�+F�k���RN��
����Y�W��4�Y>�]�n�8�+�a�ؖ=t�8��#+Lhܳ�s����C�]|���e�T�O�}���4{���
T>Bǁ��7��1�'�A�(p�8�}x>GˑrA���+pL���,Ա՗��eO]�F�^��k1C_�����ѷ����C��;��,K��8���.DV��9KN_�]��(�����r���[�D=� �v�e�~ͯ�nYW��Z��;uq��N^�6Zzq����$sr�>8�7�_�3
ű��	�'0�}�k/w���?f�}�cvc��d�W]��7��N��v>�^Ll{\��p����?��[��P�o~�×��v�]o�����G p)��<�����������������U���r�UjV�clJ���:��\1����0���%��P�b�R����r��#"wf8����RP6�ϫ�Y��RP� ���GD���m=�4����Dc�J��Z_���;�;���~6C[S��NA��pw
Q��x��k]��Dy yu����ٶqK;Xi���Q��l�j�H��S��c�,[�a_ (F�\zv��!*���*��^ �tlVg��P P��e�s.���(r�[���w�М�*�+�a����̿��CߊE鳽 �t�����l�w�o+��7>��� :�*����H'CcǤ���p�5���5�z`o��7S�Ε�;����θ��4����0�5�5�$��ر:k[��_���@Я�nn�ύ5wgNu�vc���He������=���F{a��A���W�����'��eKˀ�����+����t2Bg����?w�mr��r�����q�G kJ]��~���t��I���%S@��;�'�9�޸�O��Nuxw��/v�^Lo�\��R���<�������~�{uw���KL��wX���a���ç����{+1���ȇ=؂��1(V�f�i[ �ΰ*����z�w��_�<X��A�=���v�PBu��j2R���:�GܛVy����U}?rN��{�X(xJ}�_���}c��3`G�X��ZF�󠡷\s,\�|ʾX�Q�ϲ}�[Z30D;�Ш��[,�ܫcW�V�����<f��s d��ڥ���mgw�W<��ea�[�E3Th���$�?��g�j p�s�`�w���\���Bxf���>+Aǚh�:�U��:��9J���V�����=:�a)}�77�m�R�W_PS{��j^�O�ߜ��ٌv�3�,i]��6��g��s~wݰl���q�\�c�NB��QfU��r�q��L��m؞�ey;&eO�lE�*<����V�w�����:K7&FYM���W����U��g�/��e�����w�&�dA?նq����_�mPY?C$bQ�s�R�������x>�V����-E�L�S������FM���r�t��,b6�_u<@N`����16'apr�*���U�^�q��ʲz��?t���<�,���Gi$�|��w�in�����.�q��ӎ��e>���^��M-&�D!Bv��s����͵���'
�q�Hѱ�9�����}|�@*��d��p^`�5�J����tިvTb���sa�)�+���6���\3��NW>�a[ JksP�E�v|��W�5˳,SmJ�Ў%������!آ��y���6��;�}'��>t��.�r ��~��y$Dm�a�@o��3usp��|HC��U��2�8j��Hy�ve��Ќ�t_��A.G�ͧgC�2|�ү����q���8�R��]o���۾~� 3�B���|��_��������w?���߾7��/���7i��Dڟb�����p�p-. �_K0��v=�s��hN8Wk�N%���<�u�t}sf���\ʆ�3��%q¯��@۝85"P��P,J��E@���G=7�~/O����Q��R}���y5L�X����
0�z`ޥ��o�<jk�J5�Ji7 .
�IP2	u�T��h��i��
�����H�Ȕ��!�����ha,�����Hwec��w6�1F� ���2Xb��>�Q� n-4�f��1��:7�&.��9�ڏ#iN*���x��&,��sw�M.�B_һ�0+F�5�O�� �}��z�j`�a�q<.~Nl�.��Ry�;�0�'<bt*�8���x�B9�6I�Q�5���pX�5�՝~��4[�n���`��'�b�:/�~����9_1�d�j@�2���x+�u����c�n�zu��yą%=����y�P8
��V#y#�!��zr�^�yFz�P����Ą���a�V@�o�)t�P_(ߐ?O��	ԙ��M>闺Ԩ'X��ϙ���PN:�l�]�h�Ȩ�JC0����Q�<�x�}�o�c�T�IYx	}��P�}=9��Ig��-v���}���B��Sd�Ncu���S	g/R���*/���������l#�;d�r��xK���C��Q}�1���9]}}�6��)b�a�zuH���y�r+dD��6����'z��ĺ�4wd�;���s�uq<q�)v�@����93C���2_z��<r�4�����㱞�R�gBO�xg#�]I��*P�V��G�Nf����������ι/�����>�p�W��,D>�$��\\�w5aX���d��.}���N�#y��.˭}�{��${A�L��+���BC���~ |��TJ9/#��7h��U��F��C曰�����M�cg�b���� ��$�q��Կm\t�}����c���tq@�˴k!ω\�A|��uQF� �j�)�6�w�b	)m`=���U8�/ȸ�r�L�^��+����[A��T���+('�`��$���r'x��e��O��}��#�Ǝ�{���IE�]f�JjT�8�,C�G�����D扫��EL�e�#z�. 7�e�ؚ|���l�lQ�@:��2��͞Io���"�x�)2 db�+ ���������G���bW��O�}�M����2#�r]rʻ27���-&���)����m��c�>�8FG���Y�A�ZGg���Y�������^�^E_a� 2�x���9ff���R�F^pY���a�P��O�И�2�H�6�~�?1�y��qJ��?�&d1ԙ͌)�H"��/�D%<��a�7y�z��zŢ/ ���U�̙�K��~��F�F,�[�9y��Z�qM�ǂ:��]/�Yݨ�󷖫�KI7�8��c���~Q���)}��2��ik�]5��:�^�<3 ̔�6!��~��&8c�A���6��ǵ�ܾvd!��Š7���K0 ���z�=�����
X:����/�����ܟ��o�{��ӯ}�k��}�ޮ���~ �������o��?�~���w^���y�R��t#v`7�p1F 6�2�F���y�VJ�Pz�h��y��p��3��<��\g�=�A� A"�'����L�?P1��㝁��E�i��P����*��~�5~j�t�G���Z��O����Ƒ�=��d2�����^ۡm����$�s�ҥ���~���ҟ)K�܄�n�b��U��:׎��4:di�(�y�3AӰG�)vv�N0A��� �^�8��hYϊQ����AL#��͝9k���R��!���� �++
#������K��Eo�׌TmÏ'�S猝�ǃ�Sp<�S���0vRp�߯���A��$cl��YrSvIh�Wp4Y��8���k������Ҩ�E�,��l�$fJb.<tH'���ƛ�(�[^�r��p��\�۠�,��d�6���"���˅�x��idsY<yi-t���З�S4@���.��|&�ޑ�&�d�X��s�V>��*��'lٟøx^uW:d� w�D��9�I��1��~��a�=ϱU]䗋IYMކ|�t�(�k8_�KS�r���T}���p<q~��+zVd�f�Q��<[t����ܐE~��#<�_��&�qp �<]��t|�4�hm����I����R!�i4�ɘ�0��#M�̶C�W죋0(K�^����b�᏶��ʃ��L��/D%N��%��G2���*?���E�/���:gnw�$k����)hC�MOO
��>a���x��l!M�Y�0��sk��ߕ��[��m���	u�(-t~�y�+��ve����U%��γ���#)���yu���)Nw�:Mer��Av�>���P���:49�"Zܬ���y����,�Q^}��`�=��j��ؚQC段��Գ�=�h���T)�Δaf�gs�������_��*�e��5�T��yRu���)�x�g�G��>B��ek�	��z�9���fv*�����w<�y�R�zy�����������`����zV���ɻ��jȂ븯��P��b@	~����S�x�We����UO5;��7����m�1p�|�?� D4����f�.ж�=r�}*S�7�(]�2+ J�Ɉ4oeGo@� ����S� �n_@a;�;����C%�64��|����낛19����2g�⃚ş�c��HݯG���l^�����ԉ �EUdHs��/��i���/45A$�4�c�g����+��i9�1s{���"dHؐ3�-Φ>C~0�B�P�B���g�k_���؇4�L���3&Cץ5pѯ�w���vt8�4�)&����r����H���i=��0�ԙ�u�P��Y� �1
�7�_�>��#�r�؂*��(��C�7���\O��߀� �܀�E,O� y�ۤ�0ɐ4)Yϕ4�0ǒ��Ο��)�܀j�|���U�e �q%�&�{��ٷB#�WS�B;d��}��H�Ȝ?>�Ą�����w�`�	��\ܯ��:�z@f��~�K��.��]]~�Y��ܕ=n�����g)/ ?��1�V�v�ނ��]2Ǒ2~./!%L<g�sV�A��%��t|&�,^�
�a~g]�{b��P�5"�-�ꡲ�ʦ�~J�8d���>�I?���w����o���?�?�K�����/��ٯ~j�SB}��v�]o׫�; ��f���������O}>������,���s��z��uޕM�i�E0�q��~�a��t��,�8N	3L�f:��=W�O������r���C�o5L��� &�R���;���#h�=I�]ӗg�bZ�Y�{U�Z5��"�����:�����{^����~C�l-��Q�v���u��#���*�m�A���l禋eLY�Ιa����`���*�%S�1R���tF���)�m�3�N{8�`�q���(#v�)�CV�˼�N����l���Ƹ�W��'x&[GA5H��Ob;�1��p�����Q޻�o�#���w�c=�y!QO���A��y5K�]F��9zC�1!��e�j����(�:�#3�ҽ�<1wT=c����E�"`d9"�B8�`�q13އH�U.�m3���b_�R�)�A?��=�z}������<H�Z̛#��5�Wh��,Y?���^�qGW�^�U�8���,�X6��eoL�;i^r~1ȁ=Sy�w:
�PWc�s�4m6����Ze��2<J�V��T�\�_�X��� f:�Fo����T�:���]$��}=GM��1ǡ�N�źȅ]T�r���ˎ<B���~U�����'�rL��!��S��*]��`���z�zY����;�_���#+�PΈ6g��P�e�Yup�C��E��;���F���{���>�׵p�4����˵mp�{JY_����H�]*o��]����U:���~&8����O�,w�Y�dFy�
�2�3�o��A暑�j� �-�m���dޔU�/ߓ�3��}�O"xW�֩���	��6�, ������V�~��toC�mm����� �ͥ�����Eۇe��ћ�)�mVؙlh����{ڢ���%�0�N��M����D�NΓz�f�uئ���s�fy �X圻R֟�(���u1Q�WF+��1�@��@��y��>ς%�uu�G�C]}|��[qvt�Fw�G�V��/���O0��b�k�ԡx��u�=�]��ϹWQ��/����8��7;-_��uqc�<��B�S��4~-2�z��L��c��9=��y��\_��F��Y�Ϩ[q@��)Cv>�{���@��������p�������ܾ�*��	[ɸ��f�y,qS������;�����M_�����'>�i���2wS\�e�A~��Md�ڛ��Ɂ�Ǚ����Ҕ��c:��Wф�E�s{�����q Xm�살OS9����C�<*���M��^�����Cw���P1���J�k?��=�#�c`�@{�����MG�� �ͭ�D����\PT_Vp*��1W�xv� �i��BN�퀹=�'��v�m���G��+<�K�� 1���u�2����M��X�w���c��t��!�<�R����%�[�ޣ��`'mP�9��N�w�:�����o_}u��������4�C������Os�)�h��?�R��7���g�j�z��m�6�������S�f��`k+��Wv+���������'�������c�|���o��v�]o�����G�����'�y~��'�q��O���K(�p��MJ q)P�b|�Wf�����t9�EI��*¨h
�4D�3��{�(�����J(>ݙ[�^��(�D�����3üf�	-*��:���~N;�s��w_����0�{TZt��﫱z�U�f�� λcz�w�f:k���Oj\s��>�lX5ϓNZ�]h0u�v���D� �4,ɘ���1/�����A�+u�Y7�*���n����mS�8����d����yw��b�o��������f�	=+P��1I7����$Z�52����<�����oe����q��0����.F�����kDP��u����Z�A�}�V��"
>�c�4XU��v�!��S
ms�;�X=��'�9/Lu>�����������3�8���7Sx!x �1?�I��0�g�∙YwN�=�Y5��X�S�%F?�Ȳѿ<�Ơ;����b1�d,0�X�K��^���訳����N�)��G��Y�Ci�e�	��u9;=A�'w���(�zO�G�6�9&��&�\�ɓ��L�(�=h��U'̵������l������9HYvI�|~I��%o���um��γ�M��t	��&�0�6��e3{a����]�tN�1`�����nh��s'偅�1��X�#|���[N%���0�ý��!3~��p�6R����f\���}�;�n9��]�O�����}�"�B:}�N"�Y����0w�r��P��c��*��g|�8����4�שA%�Ⱥ�C8&���2��oE����Ԅ�̰�Ig��;-oN�:1���<wzI�I�,�xT�*�|�O���,���*]����_[�t�	�~��3x�Ѐ�w '�+/|{�l�Meg�X���6����nh�dw} |����c.�y�z�I,�0|,�Ґ��nO{߯ř!�'�:j&)V}�۾�d��8�[�<��܅��f[4��ުb�m5�#�4��8&^.�7`�?�-�"����ϩ�6�9�8�����ul<F�_�7C{S��"��Aʹѹ�����Q/71����.7Ⱥh�£�e�L���	��w��Ѯ�lp��t0�<�z�T���h,�CZ~�v4A��[}D��>7��r�J'w�o����K���h]������EX�> �^����H?�/��,l�=tю}	�Cig�b�&��/�']F���㐴y�ܒ��F���T�
�،��=�q�6x�(r��̈,n�y
λ_,�~an�^�6��l9���;rtcȒ�I���5,�J���g"s����lRZVyH}��8y�"k�Q�Z�P�\!���1��_Q��P��ֽ��Ѷx.N��1�b�f�k����!C���85h%�mtL��e����>��.?nx�<x�̓�1��#,��a�e�:_&����>0N���]�Ӈ�7���=$����u:wd��bǱ����д<i���_}m2�־�r}��%�޿]Ð��s@欷|��RI*�3F��{\w�?x*��<�)�6��INh�e��D���b+G5K�Zf: -���y�}^G <���O|��w�������������^_�y�ޮ���Z׏" �~���>}9���-߿� b?y$�M eG5wx?C�0�~~������TdPL0:����H���;�
e��W�g�ˀ^g/�%�GD�)�B�)?/$�+�_@_�$�Q�w����� ͬ�@�N���|M/& V�w����1�s���jX���Q��-)p�ti{�XsYެukt�1_��B�<�-���!r���\�{�+����U�/��s�tE�XzE�rf�i�<E�:^l��������a����!C��Lp6<|�(M��o���;����������<M�%1N`��`5��p��O�3�Q(�Wt8X�X1��/���!�$�07���k �c���gg�mtA��^���,θ'Mf�tݿ�* S�_�zeb�Q\y�<���f���9y�X�}��&r�/yb0Χ;R�M��N~���ε�K�Xeag ̇<�[t�%+.�q��m5*rӂȣ�O�;OXD��'�3��\�'�E�0x��!/���x��.F�t�iNg��D�AU��ǁ:kЈ^��K���7�T]���钽�XȟS�<ژ:B7f\��8(=�9���Zl׾hv
��)|E���ѩ� �jt�Fh�1��(�c|����q5O%lʟt0��䀡�q�;� ����,<�r��G|p%��0����^����1����c�b��S�-�d�\z��9� ���K��n�H�!οzn��W����"*���G�X�,F�i]\�ܯu&��3��;��X�x ]���N�r�LW��A?:f��D_�Y������vk��Qv�5�b����y��ęZxT�����m�7�R���$��.�M�S���Ӿ�y�9}���~F���3 ��4�Nq��QƐx�/�����Y�݅��h���l�vj��_��������*r�d��N
^|ޟS��l%w鮌Xy$q�<{d�K����2v9��C���L�s�nư2
�S�x�N�x�*/2��_>m��k�1�ʙ���Վ��d)l���\���n`���njbCU<�2@�tS]$��Uoj}>�ܛ`�m,P����:��G�e��
��򳿫x�u�҈X�������>�f�o���|�n�%����3�(h����e낎҉�-%�7��+�lD8���?N��ȯ�X3��/#�	,�_�۲�5~��-�"ۘ˧C*��s�`D�a���	�<��^u�e�
^ܱ��Cqf}�z����<{���:'��4��5o�UX�n�Xǻ�Yx<|�=89|<��◊w� "�k[=�A�a�g�6�9�s�`�Ԑq�|X�u�4i@?�I�:sNS�/ح/�3�����R�~�8lҞ�-oɃ���I,L�`�1$P�����uC20�{��=���&z��d�=f�#|^�i!�ڏhg�� y/���S�s瑠)�`��LT�x
�_O�:Z�U�`>긪���ڗp��C�̾�vI��˝�.�cV�3WM���e�xե�[���ӳg��+�=�|��><�k�����<��]_����U���ږ!~�.�K��b��ҙ����씒z��5���#��p�lw4�B�;8�=4�U�3�+�B_�7����dc���Yw�ѡ�&����=����������>:��z�ޮ��\?� ��w}�[������|�׾�����r��\)u��R<YjJWX\ R@���`Y����4�J�m��EH*�������Yf�F�:(�r�ct�S��l�(� � ��"X��C�\��ܬ�e@+��W7�����˦N�I�
V��H��3u�i����iE�Y�W�� �^/w���m�N�4l�0�����Hm�����C���.B"���RfF/�6w�ٝ�3�Z�u3w�L���N�c`���l��z��f���8�o�����\l��;�u0g@���ShF{��:}>�N�h�m&Fm�?>�5k��~�b_3�$ߥG{a�+�j��K#��ǒ\�!��C�fuʡ5`|\���ӧ��N�?�oZwԟ;���!,���HۨN��@�}��g���g� B�,th-+"
�q��gZx���G���~����i��V0'������&ܥ<�-���=��5�Z�>����A�;,�����w�}U����U�]� �3��,o!h�iY�ľ�Ö݂z,��U��1R����&/p�'��P#~�NW��;�;���q#t��C�J�>ߤ��+�k?���߸�ɯ��%���:`\tq9qY�'�ՎY�{�bT^��4 N��eIV��s��	�Q}G�������Kބϳ���2�u!��ȏ� -�dKg�Q�'�eFƂu��d2/�^�Y��W��U�[ҫ�6:nX�~����U�;Zk���ݧ�#{��!�j��>Vx��P�Gu���f	�e��X�>X7�#��FN���ԍ^�T�d(���L�.�N"@pλ�9��50�6�>a�-�^���F}^v�UJ��^RD0q�A������y��%=eey�C�[�G���!� ���ԏr��.��l��o��+�/����<Z�D��Qx@Z��h�lt����#��(aUF섆����Ff���%�����+Ϣ��A�!���虩��#�-�5Q�@.|RT��D��f��\ؚIf��J���N�S��6�s�g�v�w`O*���3ڽJ�Gf��9��v��x����NM�E���"p?�r���h�1��Ľn�����
=K�RF��?I?��?��2��b�q|u���qT���*�G�-����^�v��6}�s����qf6;dm
~����D6%v���Uyde��Ewr�>=�L�a?�}]�b�r�&�"1�fw�o��׮lۇ/��R�u,��ѯ5��5�xf�z�u��S�|������|��vT�6��/X�$6��7��UcH�i�gF���������;�a��A�G�t`[�`1Ř#y`�up���:�8l
���M=3�5�E�?�	Fy��e&����3���G1�=r��M� �s�����O�ǌ�l���3�=�~��?��+�BD!�ն��::N��b@��Un��a�]�*��#W�!�	�Ώ�!��2τ?�ڠ��k�S��#4@Չ�[w���<�>D�9��U7��+�.�'�����۪K+����<JY)4V|t��E�g���#������65$�A�Qԩ8h�q�!HC�j���������fC�-s�B9}��ݹ��;_��O��=��_���~����/���{j�]o���v��a ,��3?�S_������?����������y�w��d\ o<��j~��� C8oL����Y�3�Y�XB����;�a��
��IQE�6Ōc�h	E�vXh�P0�U ����]��m
�/��{؍�.y��Q,_w��;m���	 c}T��zm\�>�hd������h}�| ����lm'� )pe?��;�B#>Kr�F��A��ɟ{����!<:Ug*��=ɖ�<��m��6�wJ�}��:��<)Q�2������m�Q2r���G�vPNL7�pX���4�bܦ��hXy�:�)o�n�o5��A��ϓ'���d�.ݑ�rD��#E�Y�3�#���"�.�a�[�����E��(s�iTe,�`ۙ��t�����l]};:Ғ�@�32P��Q�@������Y#���۹��i8�<��>
gݍ:"�?ڇ�t�!���N�l������b�K5n�����j���<��̱�ʌ�6��&5K���N��\�	yɔ�U�^k����"jv5,
h���t��Y���c(��&�ː�tNP�\Wu�y[���c��Q�؝-yD�{�i.`NQ�T����[A	+�eV�ꔠ.�^�(��)��I=h�/zV�if���x∹	'Ĥ<Byl�Q�wGi^�����_EGO_lm}a���K�:����;Ɓ,S^ջ��U�W̡qS��:u|���0S�at����ruW��Q�BG9�LxC�̚�}F)[ߩ���Q�)�Aqz�����"�H�ʜ�Ӭ-��xj����빰��r��SAԂ<fb�d9c��Ǉ�4�XQ'c.Y�Ջ�h`�30�娆;~f���L�Q )�K6Y\W�z���7!�%�m�l�mX�BN������=y+t��n�a�Y�0�~�3���2J���Ѓm���kf�З!Ϛ�W(����&Ԑ2�(�z؋!УB'ۈ������_��5���%h	]���pZ��E��"�C���}�in��!stA�z�o;�Ŷk�]\e݈���Q<O�U*�o�\��㋂Qk�v��9��3W���2C��_�'0Vؗ+\z�����eK�b7��ԋ�_�j
�<�D��Ώn������o��t=�:|-J�fvJ͐K1�//_lM�����w<Tۖ�&�<�1�V.��N��g�������\~aG{��Z�{�8~�M̅簀�M'.�\�jF,�����K��г%� �qՍl{�wX��Aw���.��E��-��me��M=%;�1����޶#�L�M��a�]u!�:p,2����[k�����gY�	sjN��ΓF�_��)�1�s�e����8q}��v����v�%��H����[B]�n�jX���czI#��#�>���������Eg���}N[\e1�T�&̯.��T̎�
��\�yD�g�څjON��c���P� �qm���X�����+�:�cU�����(P�v(��f�.C����y���,~��/��c�ڳ��3[6��H��xr�|E�k���2{ָ����e�<
r��y<��C*�yf��O��o�F3+Ct�s)�%O���~�ˏ?��?��|����?��O���� ��o���v�]�~ �//������?�O�����_�����r|��y��{W� ����]P
;�_�+g]��2�8���c�1�z0R�G-�1� ��$5�u= ��
�PC��	����̲K;��� z�: ��_S��vu�N�h�뫠GA6���p������}�:G����wv� ȟR��~�������r8�wg?ҹ����H��Q���-3�Z织q%[��y:���f�L�����h����:��B H�m��(�5�YY8�@�Sф��iB��F�w�;<��AOb�]WM���\�V��$��%3��H��A�\Ӡ�T�5J9"�_��}5 ���V���������Z�*��̺�F�@�|O�i��˴|4�r��V�M�ɺ5�y��⬎d�߃!k�7�d�i�.��(t�|$M��$u�PL)��z�|8���`�.��ȏ6�$�4�PUf@o�v��軎C��ٿS���5�3�!2E���Vu�y�v�����u�0W���g�\�����O{<�&��)
3�1t�t�4�g��_8����+�
�T�;V��.�q׻W�y�9�-�K��xG��<F�яw�{x��|�2enΚ��12]&.�A��th^�?bG�����>^��{�RqG��IYˀ+��t"�P�5�����amJUb����TFv�A4x�4G��E=����Bwnن+F�K۫m�t�:4�k:?vzW��+�-��y�^�jt�Y��w$-Q�>�|���:6��⸾��4��6�M�[xR��#/���~��>��2>�w�T��ʄ��WY1@�#�K,��<�<�A?�,~W�g��p���6�,]�t=����E���ez66~�:��z��!��h����~�ܩ�8�*��6��S`Lð3������?e���cq0?r7ާ��Ϊ���}�A�ڧ�̍����<�y�I��?z9o���c�>�H����+`ImT��C����n�qB71�t�`���h�,e����/��ׅ\)n=sq�s�<�kG�CNG.��^��l�j�uL�j9DO���|϶�)��}�ǓA�!�ۨu�6��vTVY<���"�������o�S��i��#i�v˷�a\ޟ��Z*o�r�����vg�ԅS�E��_�uQ�OĘ�'p�I��q�?(�ߟ���P�(��ؼ=��ٸۿ� ��.l�_�Ÿ`7SB�QOt���z2!-Bו,$:�E��xFȚ�.�,����b9����C�q~���ޕ��%��GYP�w2h���t��J�c�e�_xGz�Bf�X��>x���2��8�.sHk�7|{�S�A�	K�����~l6��Jl�<w��>f�@?��Uܵx@��a�C�>�1���y�[T� ������f�V0�F�,�4����{�є7k]ݎ�G`jY�5�g�������6�[��Z���d���A�
֜�S���+���Y��������5q2V����~*��P�.�0_�Bf�=��U��H���n��2^��N`������|��|�'����O?y����}�_�[ ���v�]_q�P >��N��/�Ǿ�����k���������������o�'��Ԙ�g]�྆ݜ[������@[<=�geB�+  4l���;B�Q�h�P$�i�٥oY��ڜ��l�u��וg��6�V����/��~���F�GJkFWW��d�`��H�v�n���#�-���{CZ�������}�N���}J�u�� �fm6p$����Z�L���(�6W�|}~�R�� �D���	P?��a�)]�|��KM�]���n|)@Z�Øm�Ζ��<ӟL�,	�hF�5Ǒ2ʍx�l=+Wӿ�E���}�aHA��/DY��b+O���i�O������@M��g���/N��1�k[�Đ��Z��0GU�b1�8���{l�W&��X���!g��Qm�*��Ӊ�c�(��|$���(� ��3�pl��bߡ����q{9 ��ۻ�QuQϫ̪|s��$F�u��BSn5mj'!�?$�Ƞ��9�8��_׵�*�ΰ�#�3��х�
�,r�/�����NX�i��L�y1�&�H0z�"ֲ�^wzH��gB��wt<?�]櫿A�9����eD�e4Ʋ{��H�>Ѭ$��!gn��̱�]��Nm���nud� =���)�&�;�ztIw�J��P�{�^u���"�K/�t��^�LG[�A��	ݦ� �'?&QV�> ��w�d���G��w����W�kƖ��ђ�yG�����U_�b��b�q��)�_W�u��`7��,Ys9u���l^׻���*�y)]��f�wmnH��)l{U>9P��� q�zͱŶ��Ȼ�;�\3��y�/�	v��9P�� ǀ�b��,�
o^zu�\���jPn��k<"�ň���S���.���o�.c� ��w���6�(�)OY3�+�e� x:�<����ꠗ���W���6�9k��/@����������9��[��[��)7���A�o(�A[�.�_��wcqɉf�C�g{v���vc��M�>���Q�^?ī���=�L<�a�_�q���0}7��fb��y)��g����}���>�����z�;����xHt%�mo��g��8�Vn-_�"�)}C�9�\�(D��)��#w��{��e*y����3��Xy��_�$��VJm4�� �4y<��۹w~����U�6q;�n���,HV�1�N�>";,mp�1�(���F�3�{������A�!�%u6����\�����Q�α�Y������X�l? F0ؾ�)�%E�s��Gޱί~�OU������7�/;�$�f��Ш#��y�כּ�-��*O�t�!��_?�ӋS����5��>����j�y��_y~�����-����]IS莭^��|c��Xx]otwk�c�-��QN�Y���|1#�F�+�l�;\��,�/�F�bWwLl�|z؋���������>���o�/��������v�]o��h2 \ ��<��/~�Ż�-�<��RS/��i��u����p� �a�ay����Ji䕌��ː)� �q�gF_i��������#�g��j8�4gDU��=�����i���~�:�w� J���јQ��q�3�ʻ}N놤���2Q���?ӍGc�Q���_�)�šuc�q_��?�A�~Wtt�&��M�	�&p>3��)�/���j/���u�c��K�Kڮ���2'W���2��6���ս#v~�|F��
Dit� 5���}��r�L1��v}�_�l��՝Gg{�}ꋈ�"���<I��9����wg���x��q�#���ʊ��ѭ�i�&@��m�P�i6�	��i8�HK5����y���m{I��BC����I�A_H-p�'y��n�Lߋ�=�s1��l&�q�];�N3aI�Y
�v�Y�>�P��)c���n�� �}�x|��U�ձ�	g�т�깃ʗ�W�\�r��������:�ԉ�qm���
�;O��\���,tv��9q���ԛ 8Fj���p�@�<K�	]�������v'ց�Z��U&��kA{�o��:C3/T���r&i��Ey�eݩ�v�
����nXc���E��i cEnF�(�\��� ��k��b�d��T�ߎ��p:���1)g��&*so��|&���<�,,Ҡ��N�#���ꮧc���K�"���Ξ�O�e֬�"�L�STXd��f��9�:�\�.࣐D�5+���S���9��a��(zL냌������ϫ*�����4�ٞH;�r�fF4�c��K�`���&�ǎ�,]�)��P�rt��7�7ʋ}fg��{ՠc���j\0�!�}�����Vl�z'���(����
W��0]!��5�c�3�AϞV>��Eq0 t	�\�1���Le����tq�����Ʌ\��]�����V3�Q�4��HQ�,NHy���u8��4G���A��m�ɰ�2�����3s����K��� ���\���>�����7�9��I������xHpVN����R.�<QƇ��L��v�o̪��X�Đu1�B����c��a���$������	o�]�E���ҷ]�a����}����%���3w�>K%_w�qr^�l<���Ѡ����c�<d,���I0��Hh_�q䂥�J�*3�׌j+܈)�����Y����󯳝�v���PK:�\��~{�c^;0��E�1�P�5bcToBނ����/Ȗ�h?�йeŲ�4������o �1�7���x�*di5jS�_����`�v鯿_mБ�2+w�� "�Q�Q�LGo����9d�|OǄ���\\Ǳ:�m54툢0G�@:���<��g�^�*v�O�ǘ���w�\ǱS�@]}��(�#�TzzY�]��Y|#}��n]L`C�Zd��%�*OA������GTMy���&���2O|��d��Ͼ����|�"fʚ�-�ϛ�z�w��vG�I}w'W��gy��ͬ���h���b'a�➮�@�<'38�p`[`�yV��i�أ���O|�7�J"��3�q�u�Zh�c�9�Զ]k��_��B7f�Q�	���4��~�'���s|��9?y[��ޮ��u�( ����'���o����������O���1N1��[�P�1Β:�r7.�g�4ی�Q7�扴�m(�v	tF:R�Q�U�F��Bw����D����sD}�� .l�l�g�z{}��6L�o�����5����H4�h�>Z�b5�k9}�S����,�����:J�@Ѥ��_�F}1��� �g�O�f��Y�[����"�GiRq^&���t>:��K�K-�ո�|iM!\w٤�7�G���Mݵ�;|9_-��4�s8.���}��G<��Oֽ/�����Ù�u^(�%�q!ΜDY:gi$�����)�	���4RV���wVgd�/bp��]��p�Q��U���_i�g�]�w���f�� �l�,e���a%A��WǴ�ØF;�%5��z$��I��S�E����r���8�ð.	}u��k�����׳�0�tJ�W���iU����o�qj��}v5��z�EӺDg=�^D�:>��Fq�\���^M�t�V�0��N&e��#��Ԩc���"e�g0�p��H���~��	�^ ߖ���jc���s�x�����9W�".4�RY~�q�4b�^�w�g=��Y(n:����=�l��UD�Q˓$r �<�^5ju����|>��1�S����C�~���Ϻ`���W4l�������|�mc���<Bwa�2K�1��=��Mǩ|����2�8	�]iiuQ^�y��#l����t�'+M�2�+��M��s��\�]�I8~�{#�zb��wJ��A0��a�͠�	r����Ww���4y�G
�T���ȝ���>Ti�Ϗl�D>3��|ˈ��:E����һ��Xf�'�y�%`\6A^�7���s����K�3�Y����Y����C�y�(�s�0,��z&4�[n�*m%0_tqp�F�l�&p�$���y���� 0S���T�%��p,i������8�괏E��l�M�9�6���^ՏI�^׹b�L�,tQ�fJB�Y�FCy]�\�`=��O��.�y�ʅh��,��[��2�f�M��>�NAY��˧�<���.ns1��5��*nE��*-�/���f0�Qvgp����k��lx��y0#�z� �>6���A��8ʳ�F�'R�q>���1�[����� �1�̟�p����l�W����v#���*	�9#Uݪ�L�����9ָh��r����d+xPWSv�=�U������2%�z�=���/�h����e���;�}��#7�Lc��S\��#�XKʰuߏ��א�g�3�����>�QU��ޠ�d@�<�W��4��*�/�Or �ifqD[��=��A78`N����¶'�p#�k�J�S��4`���ۄ��8Rύ1
	��N�������6�yXq��w�i���Il>T''��H�9/���/��E�DQ��.���7������U���f;V4<wC���jc(��2[ǧl2��;��Vr��G�y�#����g�#��Fs���,�30�F3�d�>҃��46#?�W���������w���ӟ����t�{�b�~څ���v�]o�v�P fXG�߿����/����������^~�{��?��9��0*���3����������ʎ�L��?5�.ꝛ�1,L ��ш(�i%����X�3fE�� [����E�&(I����5�5�FJ0tg�nd�|&��a�'�����.��O��i���9�i��0�����р�Ct-F�`H�*2I�t7̎4��N�$�Ҁ#�Z�X�� �jU#��iH:U�(����Q뀡�<�	��:��S�_�Gahvv�Y��&F�c�������$M�J��n��|�/tT�����h�~V���].҉�}9<�V蠼�GV��4��ٝ�0�`�W9�T���T�:�<�Qq�/o7w~��TV#�`��y�Ns��������fi��7N��t�~�XF)'�r|qmFkF� >#��
�4�(�9\����z��2e>)�r\T�Ҙ	g���	�釺Iw:�a{�y���4�W����[��i��u��g>Q�D�+GzD�1),ЅTCg*�:��lǱ���9t�����<3Wy����c���@�����HF�����*G��ZƮ{^���?ؗ��1��Xp��@����S�w_蔓?'e���8!��\��W�C�f�&�$�����l;��:������\u�[>�)gcި4�L�@8;�:��*�����3���[Ͼ��
�JLt�ّ$ eH�1A�A�]�����/�`�k����SRv���ו�g���.�V^1)��8'h���g�S�'��DۨxCe ��Ή��u����t���^��,2!u�c���9�C�3�oա*�ת<��+�IG�q�1��Oҫ��%�H��q��w��m����9X�i�@#�n�zk[��:3��ctQ���^��Uꬉñ������,��P��?�O�8���m�`�o��hg�'u�	�W������B���v�qj����t!A���tq.)����1�` ��2{x8��ٗ3S۟V@rWp|���@���GRY�F�M�qBD����^�q�����u-,q���Y�����Zx4p\9�&
����MdjU��^��ZwGL�=9,�B��&˅�)ӺL����N�;���(�A�&c�AC�ȉ����0����#�Q���"W!w�HG��_}a�	��(�VL���5���v�����Z��D�xd́s�M��-�y��������g����A?1�>��yـ؀z:m�Qeu��o�Iu��?2o�D�6ʥ�1�dL��FĀ&��v�C}~U�p�X�S��5��׷_�憎�`РP�������v���"`a�М��~pj��E���'h�zz+��������l�E�&UVH������qٟ{��:vZ��^2�W�H��Gj�Z#�b��\�u��!�7en9&��!�K��3�g[v.uV�kW}3���;�^�;�6�E��������}����k�o�������~����?��o~����v�]o����뇝�o/�컿������׿���o���?����ڵ]&���"tU�� C��Q��ùn00���z� �(����K�~�	gQ��)�� �C�RG0n�@w $-c�Y1b���J�t�mM[w�PQ�KŽ��4zg9���	�Lm����c��W/k�)�?`�1�w;{�����vMY��Hg1:�A^���g�u��`�3�Lo6�\L��vk NL�0�K�F/�0F����h��β���\s����>:3�q�[��hX��p�#��~y=0�#��4�0��R��]00Vi����:8f��g5������J[�]O�ⅶ��dAD�f�f5}w]l���mW�VG��`S�1�78q:�(`�� �u7��?��y��w`��L�jOqFjߔ`�A��m��ZO'�4�Nf�C1>c]�6T~WY�c*E����С��߭A ���k��irJ-k�,����t�`��W��4u�`��G'T'����D��]����Jә� �^e ����T�� �@S��a�G��¼����c��U�V6��3ty��mg`K9�}��ʵ[�[��E��/�;��3�9����/��=nF��$���1��3���u�ҁtΥ���wzD�ΣJ���,�u�(�9Z��"��O�)7 #1�@���N'S��mJW�K�e�.��3%Z4�3�c5,��S݆��p��g�5}��Eˣ.�$=s�U�cl��W���6��O�~�Ϳ=���;:|��6�+fD]*��p���ʯ(7��d�D[g������K
�)�qO�NYu~�ԱN;�1;�a#u���C�F]���=b�-�s(�4�<���2(+:F��0�9D��>Ƣ�g�e���o<v��V��󸌤�Y� �QS��'�) <��\��;V�]��X��aY�?�Nv(粌2��O��e�n�7�u(o�6Ϭ<W��	���d\ױ��� �e����N1��双?�p��LAv�=�8-C�X�S�4�`W8���U�>cG� !�d J�g�A���Q��^k��/xE0$�3ҫ_������E@�"Ȋ�P�#��I���f�LfQ�~8K֓��,�ε�'/S�Wՙ�쾪:�.ʣ=�άz��{��f@����^w�g�'S0:&"�s���,��<����̱6|��x���v#��ns�m�`��U��"�g�%X����G,��Lz�ޞ���6����9	[m�{,��d��t?Re]�ɪk(�՞�1,lb�+�� fPl�F�}�����˯��e����Jzjo�I���#iO��L��6�#y���s:A�̸j�Ȝ��\կ��Uyj�w�ﺾ��j+uԺ��>_�O�hiӝ-�e��o��lk�;��ҧ�s�<J֋�Gf�*�����]ju?|�������!���F��Ҏ���&A5"ৄ��ن��.�X�7��n�e ��/?��������o��?�{���
 �ڷ���/��z�ޮ��#�= �W~�W>����7������=����_|��)��]B�JIv�8^������B���ܔ�H����t�Y�UL������̨És�ĕ����G=���lk륶�op��͖�y=�܍�U�]��{�dF��7��2�w^7D�J��r=J��n����~�\�������by�����hpvlG 	,����h��!+�����EM��l��xX���
�[F�8$uyw�0x�?e�"�!<)s�+/ca0e���!5<����q�P�s�u��H��RC��uZ�)� |s��3�����|�nt��^��b���8�5�G�r�#A顋O���\w�3�f�\��5��N�K�<�_� F=�<.��ϐ��67���`��T&h�����1��u��:ռ��H�	y��N͔a�?^p���E��cZ�`�7)|�|ǅ���pZf�9�S�z�z��p�&��O�ӠO�M���y�c���A�#�by�^�?�_���:�Q�:�y���ՠ��#�;���^��/��<{��R���H�|rA@� �z|��f�.o�NBYi#����L�ɼ㸀�:V�A�N��L�C��3Ц�.Sc��ο]�x�7Ђ���p6F��XX|���Q�����SS��k�uҔ�9��Ăd1mȂx��L-���@��;��3�-��9�-��F��ű��8���l<��>s���DK�����������9�w#��.��~<CM�<�<�2Z���pt�fu�g*g�x��������+��ws�㗾�Y�	��^U��zJ�j��#�P�~���զϒ�I���*��[+/�ͅ��V�q�?�*�T��}��{�g7�.�T�_uco)T�wX�I�}��|X��t�5@���暑�n�{Z.tR3˹�G�z9�����E�����U�?[3�)��8�Xr�Ʀ��u9�y��<�tp�]�rL�Sy��!���3�ΒC-�EW��ՠ��C�[x-�k�P�áL�A�Kl�tMm���A:�9�s�X���4��gp�wZm(�ϧu�S�|w�j�M�wg��^��Sϓ6��.�}�!\����}����Ǽ��Ag��Q:Si�)�e+LOd�q����*�q���B�`s��A\z�5M��0�b�{$�zf���m�����5Yy��(��}����^y�){/׌�����.>�An��-����_�zC�;�Ѡ��#6�X	��E�^6Sf��ݘK:�E^e�j�U�c�7A��X�z�jK�Ϫ[{ �T.ra��<巗%��F��0G�޽�0��˱t���G6b1��r��<����|���������X�=���6;�Vm�f���
P>|�#�����Ơ@G�>�5hCqa�]��0O�)��19�՗�>�Ɣ>'G�כJo��ho��x����2�)�2�4�>�1'������������ӚaK�����A��zp`3-S�˼��w^���v[����^}��͛��Q���/����������y��!�4��'�3�̀i��Gdp6�����9c٪K~M�u�����!�k&�!|����U��� �pY^ϗ���ڗ_{�/?���������؇>����z�ޮ�\?� �����߽|���c�ί}�|�{|�xڻ���� �B)�<���_���."���K�6Dl�7MM����� �dj-Di©�@(#��Y�����{"l�C�ˎ���"4���ͥT|n�7����5��e@�j$T���3{9��a��h�;`T˜b�С}��ʾ0�u�y�h�4�%�2z�r$���}��Ac�-�β��|�}��������Jyp�6ME�sa�>AW�2ץ;8�/�kj7��u�:[i�sޞ�B�Y��7ҸG��ER�,h�N�S�.G���Gg�;���P��g 7� ����yd�Fم�ڼ!�i������f|�g�@&�4L��\�Sh�6X�3���G(��	��:�Q_�x�K��@�:�h�9�Y,�������낛xp�DS7��a?�U���oNÙ�M˼���j�Ӕ��Q��W$Xh�lΡ;��t����#����[j�օ]�"���ro�HD~�Y���,i��b�\&si��N5.}|��� ��\�H?đ��{
Ļ3�u��}�A��,.΀�n�#�Z���V?�yutp�N�J:�1'� �F�IB��]N;��e�)�����s3v��t����׹��m8�s�,��l3�udC&A#��oUT�]����L`�h.����0�����.lGkE�-x��ڝQ��Ak.rB�T�H�ZwBz��F:O�|�s�o�?{��kے�e�9�>�:uu׭\��Ev�22~�e�A�B �BKF�~<Y�����L��`!�B�d��HYB���F���ӷ�:��ל#Y��_|_�s���{�}FT��#G^"##"#"#��Gs���#�t.�g�sR"z�Iaݣ�='��Dz���]36����1F:$W�@�!鬸A+giw02F���`���)��n�=�-([1h��������4\E~��̢Y�_�v��6��t�Hpv�wmM�\Y�a��a������]Ιʌ���(��y��<V��;�c�x1�qfG�|Oz����ƪ�E��M?ի�F���h� sB�$��������q~Я����	zP��(�t+�w�_F�is)��;��[p�F��@IC4H��|����@�2^�����,����Qσ��ؤ����,ҋ��YƠ�H��@C�9�c��hщ�`f���~��9�>�:Hx�}��dԧ�49@��k���&����=�G��Ҏq��0�}E�ƌ%ܧ������ʍ$e��Nj�����{jcH��2��~��2#���?�����Zx�ѫȽ���۸��=f �5����;��r���5J����U&`�!���5�)BPH���x4���޸�W�@�弎fjB�J~�|r�;�Z ��Ď��+mU���i.��Ң<c�˔��c�=M�7���#�Q��kgz���$�QG�D�r��5�G���y���&�'������u��H�����6�u�>��A��W���G��/�-^��R�q���i˾L��,�5D�+�m1����G�0���5�M�T���O�~q<V�K�:�q
���j�%@�����#�w�mk��
�UGT<�Rc�&��>��d�����޴WsP����P5P�x�4�AVv�jB��c?�:g;�W�r(s޽�]�]���?|�������{om�6�`�; �T������������W��e����<5[Z�onR�"Q�7LF!���<) J��nw��%&%��R\�x�ue�M��_�u�BW�P�{�}�[P�Y2Y7
� �+��7��*�T^a7j؉)â�tT,�p<��'i]1�e��b>Q�Z�Q�Pc pc�u(�e�*E�F�D����d�C%tT�F�E�b���]g�(��`��ыEC ���]��ʙ���H����;fU�N�`5�a��B�s�� v<��ݣQ��ʌ(ߨp�Ȁwu�e�
+4w��r����:Bv�Du�8=��>�8R��]	�F~&�ҰP��#wc����� ��� G��p�H�6�П'1V��p�R�����@j$���a{`��Ypbx�H�J�<ik}�Gs#�����Z tn����H�`Uz�ӱ]p���f�wݬ���RH��2z�i�kY�0e�)ˉ.5����=���9�,ۘ�FH�H��=����9S�G�:��+a�3�'�;���k1����x�>`�7�$�'Vt	CP̶B:[BR�2�2;-T'G�k�'�t�~]�2�����V�Djį��8TC�cR�qD>K>����st�s9�Vu�,�6T���1P&��1�E�[���#ޯMY�C�^�R�q�����ҡ:/�\�R9��Q�y�󭲆�����>��xrf�3���TE#���y\�*[�rx7�Yƚs��Z��<���/��;�����]��+sz��O/܋NSrC�8�mϡ}�~�����9̭�A�@#4�R�"M|x/e�����u�>��^Gp�.�>��t-��iI_���I����\�z����:"�o���(N���yx0.�|��zy���C��`Nŕv:z�Gҡ���Ș��T�.K�G��>�����8�I����N�(�-�z)��2��̙\��q[i:��>T�~��m�%W�0��yAu��4$�k�T9F�W�'�?�@\�[哮�ά����i���e�>�^�J�s����wJS̡^{��u��m�4���֔�|�>ؘ�>�gǀ�K�a��0�Ѩ����w��1�=\#־ʹ𦴬sM}zD\_�8��8�Z�=��&�?QW���ץ5�g�_���?1wI��w#m��������Yz�<ꓩ����ϕ�����0���T��i
c�,IiL�Q��g��p������T=:���-���*�S����&�y_�zS0>C=D�{vq|g\��9UƮs�u7�a���mH��2GW��v�2��,��Ie�"#�`=�n��~E�����$@8�,/	��<��(:��Π�c��+��偓H�ߢ����L\��c0������˰m���{����R�+���_�y����_�>�ū�X~�#*��:��c�~��d�G������%�W����z�?�o������)�|9tp�kp.~���/;�g_m�F_����}�~7�e��ʦP��������e��Z��{����c���R��x9}��~:�w߽~�6�`��� �o�����O}���>x�����|�E)��yJ/v�t��_S��(*`Ӕ��F�d�o���s�gLe�zz[a��e�IŻ�ٚݥ|�ړ(ք~�Ҳv�Q��}�tC��J�+��#�E;��2-u�j��J�y�WǙRJ7ՕW��>i�V��3n��?:nXwT��~��@�����rS��[�=�Qs�����*3j ��
b�!%Zܨ�)zN�0�e���ݤɕ�
v ����'s�-r�i�x.�w��%^F�TLI6���LE�����	��T0+`���\(�bl𺤯����xVz�ƒ��}��1ƻ�6�Z����U�r�7�3?�'Nd���K�s?�1�874�Q�^�9����_r���51����;S���M7���]�|�ǋ5�4�x�U92�Ԙ9P�ۮ׺���e�|��m��n\w#'(���H��!U��ߩ���$7�$���{�De��*���Rb�R�؂L"�4�F��-�K�)Zϰ	��G�;�D�͖νe<��
lm�M�#��n��3�@>���~n��;�����! ܍�17�C=�ṷ�z��<lƋ��h�&�J�N��:��}4����SlTj$�m���uό�@:���ԛ��������vZwJ��('}��;����@{;X'�w��9k�K��1Ѓ��q+�#�v��}:�����^���Yi�t����;�)����:��իk�,����/ś�JihU�	&����i0�i�{G��`��(�؃�W�!a�@f�֌4K�R������:D�(��.�w�k�NKzR|�U��t~�{&�T��^i����L)Nv,DjZ�3pb}����r�&?������4�`�����E0��\�5�nI��Њ�\+������E���	��ZTm����W��b�#�@�8/�^���㾔L����u���Ouc��J����%�U�I[�_My9�8�z�9A;�'-�m�?:Z�\P.�/G=D��-y4t��b>^���72�CW*������=�(́��gJ�3��zԹM�b�#ψv+�P݂|I�Ey5��2HI徯XY��G���� ��Jt��M��;G&K�U�k��(3U>E}jt��o1忎��Ši��N�=%��_��� ��ǈ~DZ����$u���ٱ�*2g�A�O@��̸Ѐ�Ĕ�`=a����M�G}N�V,�i{��#��H�T��eL*�����_��0ю��q�W/����Mq|���w��ٺa�7U=2�/�q��2��7]�����ô�`�\�u�$|@hv�_]χ㑸��\���2��ik|I'&+��Ap����LӸ���ǫ7�9�����\�WA&b�0��3�QH:A'st-G��R1��k���Q���w�������e\c����K[�u��'Q7�����^�V64X�������^Y�l���2�|d���o�~͔ﯤ��-���]^;={�J��n�C�X�ډ��3��*d;{\n٥z��U=�9v��O������^�r�N߷��l�� *:�����O�����>�����k��g��̏�z�2��<0ш�E^ͥȦ[5�{Sy�֋�~0��Da��Rzu	э�]�M,ﯺ"_�C���a������+&%�9޵?�?C!Ta���i�P�;�`׍Ը�
�o�1ơ�E����ax+l�YǟW�Ѳ��4 Yl��b"7�k*a����!'��y�潏ct��RQk1�a�7��p]��rG���=_���$�H��`�`��x�O_��SY_��0AqO�cs�s2-އ��OM�;�PWJ�t�]�Jk8���
|\�'���ӧ`5��)��nc����dA�)�9Y�?�}�{�4��l3���I<�s���]�crZ�u�1�u��s��0Q�yn8�q"�֞y�����%���qS�F�N͒
�ƹ�+z��_��'�U�yր����q��q`�����g��9N����xo�#��/�n�*)d,�w�*č#��6@�>����7I7N��.#Yl����{bYX�C�a��e�I����Ƀ��dp,��(�4�:���&	>\�	|ƪ���Shc�5Y#�h�ø��Zĥ�ףa�o�R~���U@��i��,L�X��-Eƕ�~ű��3~jDX����M�A!1�0�I�\��e���o���8��<,S�=��h�,�I���:S��x*?(��<�Ѳ ���QwԱ�r8��IV�N&��	�>�;��G�!�:G�N˭�<]�g�$֜��O�����K��X�4E:Ā���;ŉ3��H8��rAh޿�vG:���2k��Y	ke؝��M�k�B��09T��8��,��:%�v����0�n	퐞 3id�T�:���;�;�\�˩y��S(��ݵ ����'��{H;\K1@�CVHF��~��mc;��RI���}=�I��;�3�dWL�r��5G}�Яt?�������B��]����<f=@kK�VЉ����a�kΔމz��"��(�K�㛽4N�	r����f���:�G�@�=:��܇L<��Y��^|��7:<��I��k"��,�벢����(j׶!+A�ɂ��&u�C���ǨLL���7۳V�q@
S��W�Yݜ��C�c���spl�8�3�3&(a���#�m�:��2�9��S
�(���L'd�Wp��]ڒ��#1��F�{��F:�88���ާ(_�*�_�?"�L9�Snc,�����^M�N����G��Ns�/k\�%�IP�� �����=�ⴣ�B�m��44�io����٣x�}��`�p.4��d��}�Q7m���u��w��C��@�1��}�A�`^��ZF0�A��>�XV_W[�ʨ�RZ༔�R}?���9�R�I�L~����T/'�E��r��S/e�c&����z��_���0� ʟ1�5�p���y2��e����zS���v������zr�W����c�dvDx��� s��km��UD�ˎ�I����%���N٢���U����}��'����G����~��������{O�9�`�6X��g �������?��������_�o?;�;��_�t�E�&8jR��i�2GSFv���B��'��	I��L}��S#B�vLq�H�=���9���S�ޯ� ��b��c�"��i�8i[c��U��\�cbT~�³�~�"��<(8��Ua��BB;*���njX[�A��|�����Q�(���	�_;���DE�w{�J��+��ݸ����ו�Be��CB!�k*�)�0�Ӓ���jʂ?�F){Gu*_P�,��f4�uܤ��h�6/��%y�]�g]I6s���I�6,(q����A
��o�S���:�I��Bǔ}�la���ҽ��G�, >�%Ecx漤�黵��n������B�/�q�h D�u�E�GG\��ӽ)�s�e�2��+^f4��'��#hF�!�W[�sT����w8�3��/���XY�S�i�z�x�ێQ��nRP�[}X���l�Uwـ%��D��Y���j��:�⸁n��P�t���c��Q��L}�#v&��=��v����q�.N0���+��Hk}ڒ˒��v���!�B�F#θ������d�Xh��Y����q7��BD��u��o�,8M�o�k���r�o3e��A=[%��2��1���a��L��v6W	�u�;������X7���i5B���o�:�q%��0�F�iD�GV���7��%��n����`ԯTnI&��} oq:��N� �Y� ��Wf��2}gIvUP��ș�x�n+?P�/���2�Y:�)��U�D��q�������0ZvFCU��C��lq^���:��3=!�>��>ed��2GX�t����ہ��>L|�̓�8�.�Xo0�a�RFZ����/�gn��`�k<����!��M�C�[���K�������Q�g����>-���>����WN����y(Ֆ4�0q��?��N�ꍽ=�YL[3�^7�:Z��L�\Ӈu�dP�qp���1ȾtM�*������Ո{���Z�L�����q�����:�/S.�����ab{�wL�HC��%�bΔ�8�	��NG}�XBҴ��R������kRrx�z���8w*k��d�׈K��IN�b.��\��)EV�
�A�į�PZ�\������b�n�폙y;��[�uG>�p�Q�ש��ؿ��l�[�����x��E�r\��V?���d�[�]�ƬK[�W�zI�_'=�>�����)�u<��lq�1�2�{:��瞝K�*d)4�N�������i{�䶅�����_z_\��E�)����F��d�}���P����L�V���>4fȣM$�x+gW���(�#`l�|a�ߵ��ƽ�R�U�a��u�������Y~,���u1k!p��qKމA�䚧��{�?Ҳ��(��q�x���@��5?��Rʴ���`� {�r�sA�1�:�}�~����vI�5�K�W�|�g���eG?�������SHK-egh��!K�e�rn�6F��������T�\��Σ����̶ַ���K\�6�I�����G��٥��XM�Z�N�-���	Z(���5�s��:�=S�S�Wʷ@��o��O��d&x����̾]n��l��i�}-6)���1�3�����������3��_L�g�}�k�Ҩn��� ����r?M���_�՟��w?���7��t�7R#,X��]3:PL^w��5e2_l:��k]�)�i�S �G�T�B���t�p��Z���Rf�ϙ�jB]����0->�0:3���8�nt����7��޽e� �_�J	�4����2U��!��7�{�J@���q��g���
�*�4���)�h�Z%�;nDz�nԵ�$TW,�Ȟ\)�-5�+6ѰbN$�H�98�~S���S�gŁ�1��M��zĉ*������t<���6�=�B4������z;pf�;�֘�6��s���3�ӮY"�aї�!�On��ϣG�>��ऌ�v��� T5�d!Eo�X+�!;�o�X�����.���� x4��߲�˘K�f�A�B�4�7��q�G��F�x�x�y��_s��>�W�<Ǥ�Y����
��i�O�/򖶕���G�?cׂ�,��P����,0���X��6�um���S�xZ��:y[�s��jR~�tǺ���1�߁vX77�qmP�2�����Q��o�.����Fa\�02�y��g_�`��zZ���w�C��*�J�3Z#��kW�/��Ha�t~9�)̑�E��6�����uW�{�c3�+�����|��1Mh�i_d����	-�2��e���I�}B�Z������ɵ˗0�^˂��@*�7\���Vtx�ʅN��mP�PG �	�S}s\��8��[�|>��H�Q��G<�QO熼k-A��8^!B���D�?�fy�|M7J�<3Cj_�A��*�F�:��nuQ�WO����C��q<���8.~WYu,�����%u)L�r��,�k8V�Om-�(����#L���:��/�W�*�hvj�؃�(\�u�~�6q�t��`�r�@���(qZu�~�����I�)�+f&��g;���Q_�2gV]�yM�?�9�{������(�� z"x�{��[�F�sX�^�QXLUO:T0�/����]�}�(���NB�S���r��rZ���r�q�Fh3���Nkн΋~�%=� ���0KF�o���c�#����8W0���W��E"�R��u���'uΔv ���я1�bX�z�RWҵ�����.܆�|�W|�U-����-C���q�oc�Խ#�9
J�]=zf������{�e�ݧ�kF8�ҙz$=` � �ȱ�ȔG��\?�u.�����������6~_�!ȱm�9L�w_�U.�J���gҩ�fcYoz�ab-c�c}�Qo�5�;�DYy���Ms�����k^�2���W�@�6l-�@eГ�l�k�S�34X���D�̿��m)O����M��1^7��-x�|9���d3f7�U���ٛxF�AG\[�ڛOW��ʫ����_��>����KٽLU{�m��_jx� �
�����7>L}�Q*dFAJT��z�*	�aN�@S�wy�Ur�� �
��;�Jg�U�RF/�Fw�ݡՕb(�]����Be"ɿkG-���گ����q�u�_�s��寇5%��dn&���^���uQ���͡ΥB�(=�l/�Z_Op�|jӲ��ht�n��RꉔXğ��r�������ﱽƣc7�4D$�4��DE8��2��~Mq#6�>b���o���)q�b#IUܤ������ڄ�뮾R3L�Tv�!���lYn�q��댁����?��,}�q�Z'-)�"�������fr��b��ʆ�8R����4��%����p`�)���5��1��dA�C����g��g�JO4�z���'��6O��m�+�`��h���\�(����1�*�j ��Q6iչP�㚅�Z�Y+��E���cj*nTV瓠��o��:H��!��Y6">ux
}I#�-iJ�ʜ2
�T�����Wy�Wb���!�H�}��q���ɲ����E{�^3���r�s�sƄ����Y1��*[�6������: y�-��^��'�4�|ƹ�\��p�\����/�B�M��yeyŨǭ9���U�����P^NǮ��v"?'���NwD�㊲m4���U�����Q�T�:����}�h`��K2e��������|��a��ޫ?���V��zU��뼝�r9^�:��>Ȏ�t����z�8�*��Ô����.������*�>�-:m�s����砬��������h��k%��.�:���DV�ݴ#OFY�o�����ՇFUA3����c�>B^Tj�u}��y�ӻk2h�'�uQ|>4cey����x�`�I�F>��.�<[��&�U�	�C����3��kuP�-����5 We[��=��-���Xý}OFk�����t����G̃��,"��1[A�'��*)�+�<�{������ tJ7�8�Sw�W���55}-�ި���{�o��������35Ơ������]��33�������xY�f2�zT'��6�L9��K{��\���Ч��ݵ�X*_�gp<l_ǈz�S�m�q���)��b=��G�꾝��#��H7i����k�rB4�@�0��~�tY?�̫��R�j�Ȩ�R7)���&��;�k�������:�M=��8����;��Z��������~������u+&�.��86��.]|FR�W&sa��c�_\���e��e���F�yx���~sBQ=5�k�W�F�B:̂+�)����V[CNϨ�ճ�Z$�mO�e��˦{�#�G/�v\�	<Y����l2�JQ9ש��ޔ:�Δ�.K��4>t���Sߙ/��p��CG�)��`�6px� �W��;��������K���b~�U9\i"Ǯtg�t(P9�gQy^[�?��rkԤu�o߸yz�]��T����h�R?�!��?��4Uv<5#~ޛ�B6�k��Ttk� ���:�iT�Jx/�R�
��PD�*�0D��EvT�їu���K}�:�C�OO��l�㌴z��S���4P`mӥF�h��D�%����Y��L����Rb?Z_�0(�|j�:5�0�=�i�|j��kB�N����\�tNJI����u�=7T����]\�-�@�.9^h�JC��9����~4`^��'������_KM<j�UQRO8K([��������L��o�c��L��)J�i����B�H��y�O�s��蕎m�l<�A�<%]{Z�}$�VC�h������xc��q>���Sh������/Ъ�`��F�?�Ox��QN�{�g͑.��i�.�w�{(M.�Q4�[�1����p�lJ�A_�^�=&���>_ѥ�h�P�����S����u���y1�7ޭ�XɹF �.���Q�����4f��}�1�e�Ok�+�{
���4�����x��aLk:ƒ߳ϑn�������Y��|�BW)�p�����[��Aw��ɣd+� |Z�ŧEy��jv�<4�R�Mu��:�>���N�PV�G�����o����ot�t>��T�-����2~89������q<mK��-��<{�xV)}��x��:=�~�����hxW���!N�>�^l�G�s�����x�vc@�i��}� ���&��X{�s4ʟ��(M�Eީ�
4ծ�:�,]�[J4�á7�Q����nUNx�� �dY/���Z�����癩U�Ыp�R�<D���,��@�Q�B�����F�m��X�~�H���e�5�z ˶F���c�����(?��]A���K����ޜe�@C��MD�k'��3���{���gG�'�:���v���ė:<���O��d��Uctr^�^nJ�6FZ�=t��;芐/�o����)�^�A"�J{*zul����s�k*�6���S��3w]rz���|�_�����7}*˻�y�Ψ���Ͷ�S�*�0n-��j�k�*�ؖ�+ ���f�ԥ}�~�ʀ�x��;�͸�x�6�]���iAZ\�g�
���)�g^_�����<']�Uo���M�㎁Z�o��N�nɱq�"��n��*����0���j�'�u�H��Cu��d�2z���h�ɲ�Xǚ�CyL�}��d�A���q��e	#����<��s�|�ه��x�m�kI��?�?�ي];��?f����J�]����щq�ߧ�F�d�� \K0&�u���ǂ^Q��hЉ=f3&*.צ>��-����ǟ}������w~�5r�'c6�`���� �}��'����������{M�޿�͹�ǚ���YT��z�P8c�0�d��r�����E$�`�S� -�)�S:�M���&�s���h�a�8��R��B��M��d���Z�,��&s,���R���:���Q4(B�ﬧd��8n�T9�e�f0P���eiPI���hOۨ��4i��A�6XT��������q6*k�Q�������an��^� �=��1q]4�/��J�H����e�R���e �P���HqC�j�ώ�y������^I�=h�8���e���ROsL�G(��LA8����j����VD�t臮k��	3t��#��|�kE�4�y!�Ix��i�W�۽���/��ӛYȗ|y<]_�vC�o���6LE͍q	㱹�d��C�yg�q��)>:fs�F�Ne⦥�d�[j�0�
�i<)l��C��-ZÜ�9ޖ�p�1����>���G|��ƶx:Q׷M���Nxo�2���;�Ң��=YWk|�h��6��5��CE��@��n�u�o�0z@6�ԅ����+]b�P����{�|�2̿��˦ |�X�pV�j�@�A�Č4\����G\.O�j���N�k������z��� ��$�s�3����y�y[J�X�a�����=	��� AG"ob9�"�gս�wG�p������r�cH���yGv�8�E��.uU�kJ��ߨkG��s@��:/e��K�M����7�Pz���d- g�������q���]?Z�ر~ޥ���t��,�%i�ߩ[Q�����m˜�8��AEJjd�kTFG�by�9yt�/�&���O����-�wķ�C�$�j:t]�X#*+��^��k��^�ӌ�����g"����C�U�-1�JÔmq9�g|�z5��F���8F���g�klgt@�N�}����b�v��㡬���'UG������}�4K�BT�?�!F��:����������Ǳ4��n��_��9�����k��S_�&���sh+�5�Cqу�]��7���6��j��H��؆�J���}��p?z腋?S^F�4��H}�A6��;nM���䭝��)0�5$S!��HR�Y�z�Y��:���\��A/� ��*ޔ_�fgP��9�]�G�(]�����T}���麿~����w"�tOg8�-�L�3�\�I}��+�J�5���-t��Rb�<Pp�|���yJ�)D=��z�>f�N�=q��k�������a\��W�i�O�B�d��R�YP �����4����n��S?c�;uz�Dq�k�R���㎽N���>����qL����x�bM��q*�=�+�����<�_+�r��k)���}|6��1��ZL�64,�U��<N�+nJ��~�z�
��w>�3ָ\�xD�ZR����4���1d<|7m�~���ex9��;n�u������^�cz']�����������������sU����e�`�6�; �������/���>���}�n���C~��t��Qf0yݴ�a�3MGZ�~�D�'�p3�ƴ�{8f�qтt�םi����f9�(�f!W���ZA�|,4���3�T�R����h_�dGC�~W�C����=M��:*
��JL�l�ܠ�G�#_�<���~��T�ǱRت���7#���Q�g��X٬3n�bGE�Ԉ?5|ڳ�q W��(g�5�T�Z��q���8�0@�>�����cOE��4q#RTy���XU9����A�pNC�����)�m�>��Cq�n�пcw�ή��ͩVx:|��=q��ͪ:ruew���cW�f�D����v�k4�%��.u��k���%�<@b��8�O���T?�E��0{�M���}u:J>Ffz�Z.�l!>�;~G
O���d�G;Nɜ����ql�������P��0m�mp�r�Z7�(Q�+���1�}���1���̈́< ����m/S1���gߘ���\�1u�u����g���`aw��\��8U�h�UǴ�/�6���e�)�y�Jk�u�c�������m�\@[@���\犇�S"�C_��D��j�����y�uܩ����ODC��S�4�|Er��h�T>J\��Q7��۸^�W?E#�}?�������p��O�#K�|��6~�¿\�+J�N�)�u�`*§4�"�����p(�NK(,L�<^1����]�J�It&�˨e��������ׂ�T��^��AqF^��Vq)�*�xs�w�~�yʲ�G=Q�R�s��>�V4"Q�+@��g?y���9^I���CC;ڋ�4�_�����ԣփ�\��Qo]�eԹM�%1F�H��_QG�kZ׉�O�xEٸ��$~l|&uk_cj}�>�g���c��tL�8`�_л?Ka�'���L���F�q�z��%t�xB���c�ܣ�Z:=l�{Q�R��L��j������jf���`f��3`(��o&3�nA��(�8��z�:�2��^��91@kշA;ʇ�D�wM'�ঔb����ʐ��x�;b.�9��q��A:W�͔w/��C����''�G5���L�L�ԉuT�Z3!�z�z��蜳~�U��8�����)���'�4������t���$���9��S��uʌ9Y�i��:�Y�g��:����(ҧ�Nu���ɵ����wl]������[u�ַ��/��1`	��Q?I�lԛ�ri"�jP>��~��Ror~��z��/�Ϩ��Z�|	��{���;һ��%mr"�_).*hv5�3�feU�(��?ź��h�Yx耴^��k�Qi�lY��`U�Ĵ����[�c�v�f�I"�Eݒ�F�C�$�fJ+s[�s�טg�w�8���.�}��D= |%^��&�^�tX�G�NuZ���'ᇢ�&�p����e�5�Y�sG�i�5ϔN���k��)�Cĝ�u�klݿgB�r�H�j%q�,�ANغ8<э��c^G�\ ���꘩������׀Kݰ, ��Z�.[j�-%�r�_��x9��tx���ï����W�����~�~��_��i�6��x� N�ыO�/>x�_}�^]T>w�Lf�w�"P��ct�q���X����{���,0D��=l����4�:D���K����a��u��c�aj
�d�S/#Jd���*��Bd������[�ex�����5A7�?��
�ޏ)Zy��
�84G�3k��P'7�j����7��y��p��S���JqQd�ԏ����5ꗛ��#nոU�T�HT�}�9y���q���e֜@u��(ml+n`��MT�4�����G�䋊�h��yf�>�4�D6P?��PIeY�����P�V獂FH�)S;���O��ֶ:ZP�ԣgqgpgc�M�f���,�/OV)�Vc�p�h���r�>� 6��WI�Vw\�D�ܚ�N����s�f��a>� ԏ�V���Ε���0�\_z�w�����]v�:�	�t���̐�l
x���Sy���Khߟ��m��5Mf�c���J�<�CJ�����I�M�]=���Mڇ�x�ZeD\������<��e�#�t��l���瀞�$Y�s��ʺƈ늷j,��-�%�	\�^E��1��5�4�k#�{���q���6�X[Y��y%���o��4���48-p���x����"�(	�gԠ�z3i��h
�D&�ƉԔQn�4�����5Six�F*��z�M��X�Zv���Υs���t��h�F\�P�/�Ѣs!�:��W:���4
n����L��wއSdZ��`Mo�5�_�;�d�u��v�v�/�Ty�h�V�k��<z�y�z˸V�.����+�U�����06{2|�}4�ǁo�o�!����H��M�� �q�!|���q�t�?�\�ڥF�8��7w���,h^yR>��@8�����7�l�v8w�l���C%�*t�G���ycJ��q�c}�<���2�/��l�o�0@z���˨_0���i�Y������w��6��wqq!A�;�)g9n�p�,�ǅg6��q�>/9.1�*� /����q�A�_�����ڎ����sV���
�JoU�a��;6M$���Npӥ��N���o�g����ܐ��wC���:��*���w�@Vǹ�h��ܝMQ����^�W����療�R��:�Q(�SRGn�E(_]�at�N�����J6�LX�N��@߮z��aF�wڊ��	h�^�x�֑��J���~�kMm*��s���I@��f�w�}4�����;`�D��{��8_�ɹ���8��GY���7��e�|���K�Zd�w������b	W �F�ȵ��3--36b��O�O�^��`y��c4yH.�2r��!�!��Cy�{Y�&i��]c��.�{ꉐm�Ơ�:G�4�����F^�,�����4�7�Q.�E�p�-2���5�!�B�I�����Z�u�7Խ����iP���M0��K:�����2�n���u:��#�m��r�Sz�эJ#~�M����2O�\.�߱_&/[;����H{}\HN��5���:�[���k�{�w��/���՚� �{T6�`�<z ��W�������+��8�wSn��;c�v����W�?���u�k@� ��Vҕ��l
���&�$���ANo5��ݷ2w�c�Z�.ͳ�'�+&]�բ"�c{�9��)!���� �F���.��:�B��#��iϦ���Ʒ�����~$��y7#�R)1%}78gv�]tS���S!=�k�\���'BP� u��[o�$����8�c����ki�:�p:?3����VoU�/_]Z�rRU�nʱn�l#��v t�;�h1�e8�V,S��v#��x��l3��W%�+�5��j"�es�Wq����A1s��~i��1�F����]qli���,�T����h�5+'�S��gzW�}�
m�E=e5^��e�\7%�0�����y�����U)����[�c��/���E8&�>��xg���y"nU��[���QB-5�0uW)H��k��x����V��?
�6��y����u�Of�#������u��LK�jt�cn`<�3�ڃ�l�xb�⥊;9����{4R34yJ>Ë���f�ƺQzv�� �ds�!���sBZT@���f�D9=��k<�Yl���S�烟��f4��č^�.�Psyy�q�OC����(�� "�
���ա�p:��ֲw㧡��jw�?`���mԝ'�:RCYic�M�7N���)��1i�S�� [#�Cz�1y�}S>Mrbpn'��)F�ի�^����4?���Ѝi�]���#B�zXs����O�^�8\�cL��~�}�yr�A����Ӿ^fI�c�ZzP���Σ��.��Ic�8�z3������#t������L��>tB�%0|��)샞�>sϞ��ߌ���iA_�륝?ĀQ�e�y_ϵz�f��z��r_��X����{ �d'��S�ĄqG�8w]�Qƚ�_�x�E�\l��:����A��Q�Fݱ����L��k���4O�M%=��M�t��u��2�{�tW�"�fӳRBF�6^��k@m�\7��v}�2���^�)7���}�ݨ��{�>���h�A�Q�:}@۠���!�<��������ӂ&M�b�G�W�����IP��}u(`|,_e����8��P� ��ℎ��q��"�l����+�nyt�$칰��Nu��� ��+���<�o�GJ�؉y['��C[׶�1�_��N�
1$�<�^�����d��0�ò�^�h=	��q�K���\�;����ݔ{߯~?\����������j��O�zw;�E���n��Vf�m����S~U9W۩: e��24 ���d�4]V־ՠ	��L.��v:�s�d؄��a�WEA0]rank
|�з(c���XB���<� �W�J�_-	G�F't�`U���'xK�;W��S��!��O���u�+�3�%9_TNV̒D�C_�Э9�N�G_d��� �֏��]��H�G6~��A� ��mkh�u:?�='�����tr.�}���ѯd���M�7�&���Я�W��p9ʬ:���F�|��M���d��<�l�6�]�W^n�m�=LŹ������G�20^�wg����D��ʫ���ٲ�������ذ.m{D�(B�t ���afpNu^�2jKB�6��<�pv�Fq�i�'OQ��_���xm��A�y=%ʯ�?F����� �9��d�(os�A�݆U�86:94���d�u�#C)$�����e��3����4��AA)�|�y��es�`,�g�������И�1�sj{<�_��j�t�^�A�C���m�{ꐙ�	���A"'u]�u6�]���X�<�,�{>�E<��}Q�,�4h��D{:���|b�Y�ޯ�Q=>j܆Q��:�GY2�d�lkM��ۂ-�c��w9�M���,V;�@Fn�ZJ�����W�0�?턎��Vn�t6��z#f�g�}�W�u�U���s:^���*]N�|y��׾����/>�g�3e�6��<z �w�w�������΋����e:�G����pM#H7��o*زoVhD���K��pn�ڹ�� ���zR��r��T���Δ}_b� ��ޯA1�1\I�k}n�XF�������u
�	P%M� u�7գ�w��͞�*���_�W7St�c��'0F\!�dJcz���"N0,:ێRw��7b���66�������D=��5Dacu�=��dA,����*�8��hԧ������8���������¬�C�kM��S��˕�#�&�]L=��4�cꊢ���\q��`����\k�����)�x�PSe�:g�,U�c�?O�t��4���Jw�9;��!�� (���y�O�<�ɩm��	�4v��IiP7K���Nl�q�����NVwB�q��=�ӹ����)��؆�o��M;��j��S<L�t�i*�$	Sq�a�fG��F�#ml�7�.2��$�d�}O���1�;f� ]��e.�z	�6���A70� 뎞j���'��M�w�*O�ֿ���*����4L:�v�,�i0�O���U�L� �	�������8��eyU�+�X�"k=��NO���Rj:��U>�o�=�d��f���B8���$�eRߘ�wcK!mj�[�K���14	�C/���eAy��
����(8`r����ugt}���\:]�7��ڰ+������}�W��Ck2.�g_7QO0��|��y'.v�Ke���.�_%��ˤy:}1�>w����]C�b~�Jk�v�Kك.��t]���NWy�����-�Q�F�G���57�^N»E.8?��<��M�C����%_�s��:6�B_�|]���l��_�;����X8#䤻;v�6脔G���H���*A��,��U�ֵU�c�]�xW�y�чH_�J��N���*�,BLINP�2y�,�.���L��RA3�!�/3���x-N83t`���j�,���}�.K�r.�3w�PW#�y�{H�1xf���mK�d�x�p5h��� U���Y��&�����>�=:���G�'�_�Ų�3�����q�%hG�o4SI�;���]~O�1���ԙ۾�;��v�{��'���m�W\FP��ݾ�<�e� �z����F�]�
U9�yS:a��:<v����ks�������oԡ�5��J���+"1f�ѨQ�Kr�y\+XMz�UЧ�N<f:�1�"��8S>�1b�����s�Z����M�����������t��P�~&��5��ӂ���P��N�
��oWo���{5x��%���?��S�ʶ��
��-�ߣn3L*�d�d��j+ýY�%XՃ-�⊶?0�hkQ~৲�y�^4m��/�9u�Fu(ӧ�pGo�2]2I�|���ލ�Xآ�I�4T�Č�D]Pe��i�s��N�f#`��{/�~�6�����i�x�$�������_�4����~#��m��Z�c�,�>$��
7;���1�<��p]�3x^�*�B{���}�7���b��䑁1��������{Cm׌a�}��X'tbيI�+zt!O��݃o0"�!{���	������4ѳ.e%��2��問�u�.o�^q�1�u�[�qi����I�6�+>0�H��X..�)4��������l�
� P��g��{^����s�����~��|x5]���.���	��.!�a�i*��߹c�a�=��P1C�~Q���fD�~ꬽ�7���EdWJj���;��w�+y�9��(�j�/v��U�=��8nQ!�]9�T �/�ŕ?�6I��Lϥ
�o�|��v�O7��|����s�_�-�U�7Zȓ:Mw�T���sǑ�IW���Oj�t�A��σ����q� �P��.�"T�&el|���N�s�;R-U`i���q��:�x��z<rv�źP�K"mE<�����U7��Ϭ=*��+�a������/N*��+e��0G��`㐧���R_���S@e�^��MH�3�y��i}�sb����/�F�v:�Z_
���;�;���e
�"ͬ�56vL8��%;�M~����zM��Q�����/�\I�H	��>3v���W�3># g��((sg��\-fI{�cr���� ��A�$����9;t�����,��Cjh8^�#�ǹ�ʆ�&���Լ~zY�u�3����_K׆M2A�U�"��;�2(��g���<M�<�LfiC��@:o��υ��$<Ez)��=]�]���j�ݝϋ�z
FY��5ޕ}��$C�[�����g0 ��]'��d�Ω�$��-.<m��6]��S�K�Q�du�8`W���wĥ����Ӵ��7f �#�Ah�6a�r�c��Tt�BC��;'%���ˌX)����9&~� Z�#�!->e��,��Z9���/</2N�����Y�Q"-+�kc_�.w��<�h�Ičd��ѷ9Y��8~�{)���?�4�i���	�v:n�.$�>�8��X�a߳�$�e<�Cp�?�0m��q��]� �צ���
��8�DNgocG���v�$A��P��C�7#h9��w�.��iPd���ʖ�_���R�|J���H�{)�q�C�w��ɢK�`F�\��/d���K�60FS5'������p�s�	]e��`����j�ccƞ��%�,�W��N�u*J91#A�zu w�edՐ��b����=��W���u~;�=��b����[���G]��S�G�n��`:�G��� s㱣��
L��:&.��N��V�k���*h�ۧΒ\��<��X�,I%�O��>N��;ܠ+�u_߻�q���SQ�9��3��g+�L/��9M��g�n2w=C�ޣ�z/\G��^���qM�g��}�M���;��a�`�'�3ǹ����%��4πmҟ��S��!#�������yY��E'ЄLJػA��G���u�PUǻ��^O�[i���p�W���
� W�M^�	`�w�ϫɊ ����G+���6~vIv�AR�zE��I�k8EGw���])5� ��@[�-KM�6�֖����R��z�!���c�'�9�	z��똴�W�Ю�q΍�����B��} �U3��*,����P���s�"P8�
�q��;c�w#O�e�e1��i�a��e��g�$;d]JK����V��r]�g�;A-���r�CI�˹���u5��&<�J��ei��U;�ɲR��o�]��:G��� �D<Z+�c���N� �*��`�c�wfFƄyAu�
������Sd�M~��0���xr�p�q�-�Ay�wK������Ir�6�����P3}>����������|��o�����Y��6�`�O 0��׾�ٿ����~��_������>�]���Pw
���Kɕ7�K������ Az�
͔�72Sw�B��t.)�0j�SN��s!r�
��>���UQ�Z�!�x�|*��a��GA�hb���7�T�t�C<�w(V��h�.��~n0�G1�g���U������齯�|��52�������6d?�q��7Nnn+�37o���nn�ܪ}cv�y
t�u�46��z����g�9d}P�/��.Y�X��7���V��u��'��w��u�t/x,���r�s�lY��"⇸^��s^/wG~zc��G���}�yN7�ư�[u�u~M?��`4b�����F�ңA��TW�et>N�Q:�^�w�r��?��=��D{�%�%�1��m�ܼ#=gA���r�=UVe�G\�u���L��i�TwnL�:?k:��e��u���zөG7��{�st+�L�Q�?C�;׮�,o�g���5>'�Y���V�����u���\�˫�+�u~�O7�����y��1qu>���|�Ը������M<�daOy�wυ���E�5����i�<Տ���u�=���m������^���M��.��s�y��s�Z_��mR�}{.�<�r�X�G\��X*q>9.K����������9]~q����>�8�O�����ꋔ�_�Syu�RR�\k��I��b��?��q��MY�A\P���
_3;�Z�"}�����\b&:�-�}���I�G��f�kg6�����/$>U��Bq���I�|
��������z�_��7�ؿ���W~�>;|P�:R���`�6�ѯ ��y���߿�������������r����������3�ei�b�_:��%���{�zQ:܍1�&l�S�w��dK��O�M�i�)�שG3c��6L>2}���Sw��Ep|?5s�ִ�PA.��1Sj�|OZ��h$)�B���s��
���0����L��.���(�Q��	�V~o�W>�q�z�>������ꅕb���^|���=n<������޿/=�S?�S�a��Sx���pr-���G5����p�_��m�Q�i��=�޽y�=�q��
�.����M}�p�8��nǛ[�'��K�QV��0��ӂ&����ʤ��E߯m/%; u©t[���ӹk�с�2�E�'�dL�N��q]�_����ۗz�Gc���)=�u><~�u��@>�1o��kݎv�ҏ�Ή�W�����w�/�������{m�Kx&��������cY�c�k�v�����J�d�/�.�*�>��Q$������#�����8I���=8�V����N�r��;��7d'�Tk��K�����<:�m�,�㼹Y��f�����:_��C�>�4������>��տc�����(W�R�_�7����Ϸ_��H�8L�T�H;18���BF^;(�́����ƬL�X�0�@a�@�1�{�y|f�`*��$���3}Evp~�e���zP�4���f����%8H�T�3�^ms��n*�k�o|�G�����ݯ_����/� ��� � p�DKe^���r*�����o������W���O��?�p��)(�2�ʡ8�eԟ1�⌾̖=���1�LZu��3m^�Ţ�-k��X�Nջ�mKL1(N�T/J"��
�ک{{�>��ej� %������Q��N��+1��fn� �_���M�a���w����}�c��φe����G���H����j^;o�l���)Yߗx�����������e��|�g��W��-�VtRaJ��������Be���^v�;��o����Q��Õ��:?�凅׺ε�g���������y9Q�M_�Q��{��A��^sv�뾰��:�>�cr��;��z�9����~�ϥ�ǣ�V���Ν�G[�+��6^����.^�4�տ)�/����;)��M� �O�t��b<���=;���u�.�~�0e�2
7������:wǬ�g�/���+�P1�iz�h�k�<H!����T����M�1{��S�ū(Ks�7�Gj�Q� �_N�z-�!}��W�����~���?���_\=<�D�l�A��� � �o���w���:}��a���:ǔ�2DD�����|�i�zLQd)�#�wf	�!�j�}�/̉�������Յ5�2�1K;H�/i~�����*}o�]��8���qz:��Q#Ø�4F9�;�JXW�B��BQ-�L�Փ�`-
�cX�����U1�$P#k�����o�wʲ �N��(m�rM�{v���<�x;��ؠ��]���Nx��Gr�a�����֩[By�9���svtwi���Ug�3��ᶛ�������n:�Ow���_�5+	txf��C���x��S�C���\���q��k��u��pj��\���+~Θ[���JY)���5�z a=��q���k�>o�u�,�=A���#��r��zY����<#/>����޿�3���u�z���N��St��|a[�����}'�={nW9�g���T���:�|���z�9�\����Œx�u~��wQ�N�h���}\�6�R�{f9�῞�w��c��[��y��=U�S�����y:�_���o����ze���p�v>��i���3���n�Pk����w)<�u�m<�:�Np\ݛlMX �9�ӼK�h���^��š���k���Rz{�8�󛿾���A&���7 �{�#���c�������D�0�_'y� ���N�O�7EJ����7�2&�8]�<�u�S�/Y�s��Jl?�)���z�5@N���O˔?;������*�7�`�x� �b�Y���x�G���[��7����q��/�˜q�"�VN�k�o8���Ӕpj���}2�����0�ɿk�ٙ�y���8��^c4Y���I{��#j������z��9=�O�� �$��C��3Z:��w���6����0E����X�Ҡ­��ۧ����f �O-����	Ap�?�>��v:�y�='�3~?�I�}8���e�y�u��c��.���������N�3��w|�V�]��cz�-��^�����p��ڳ������8n37kr�����g��[}��v���_�AcE���7�c�%)ݍo���e���Ƕ�oW�C�����6e�����}�-ͼ���N�WZx�u���b�o��l�V��4�H��j/�_���P������ߋc����?6��:" L3�^��~�1h�l����I�����b�o��S��AFFc���A� `mڻ�(�c�_ ���:�����'o�ص ��#t��w�=�uni��=� ���̯6hk��c+(�i7��g/?�~��/���{����ˋw�yg���`�6X��� 0}z��+��_~������>����X�.���d��}f2E����<-Rj���t�W��Gbe��٢��������ܲ��7�����hD���k�vrݯ&� )���e������ā�$&#"���
���+ ��-d]���=%�	<q�k���O>�>�}�J�Ņ	�Ř����D�R:�7�`�6�`�6�`�6�`�6�`�6� �������j���!��eN;P���GC��?�.�e�����_�L{昿�����8턿G?�Y������҈��S(�;�{��;rH����p������_"�MS���˩�A̄P::��w��0��ǫ��e�~r��w��_������̟������W���i�6��x� �ʹv���G������}��w_�<��KS>�J&,턷��O��2ϩ����f4��:���k�`��q���ɣ�p�|����wy23�@�`���u�Ϲ��)�i��� �oc��u��֜�6��_+3֣W��?
숻$C��"��]��7��x���Z��h�J"���i���k}Ҷ�݋��$M9�Щ&�L�V�xp��n���)�_g 䚲� u�jߒ(��Nө}�C��P�����u����Su>�9(��9�[º�t����6�R�������:?��o��6X�����:����}�m�	���Q�����pN�����j���p㤧�k=n��1�^��
a;4�~����_���wr�
����d�=�wj>�d�M@���xx����ze3�0a����Z �2]���<+�:�/8���i����Yz$���ܧ�5���뎧ɳ���ڙ�>�l�UkEo�z�uW_�?{�[_��7��_����s�ϽU�����R�c{�6�`�$ �O~�����4_~m.ǋ�阍�M-��~�����"���vAT�������Dݱޣ�J� ��3J�}+`��;�GgyB�z{������Γ��|�X�U<������3ۇ���O�F������kRB4~�����ߊ3����O>�E?�l x�}�������$��ˠ��6-�N�&2�����o������B�w��C���
���c����2��eݼ	p.��)�\��\������C�}����9�����	�C'u�7�u��l���ܮ>���i���0������v��h�9���o���o���}r 0�t��\K���"�"�� �V��Ů����b����m#�$�c�_�|�kך����Ӄ��Ȝ����*y��W��ݵ�㱏}���p�^\~�U���/>����~�"���6�`�x�+ ~���/^�<��t,�t��\��Ү���W��6 r3�̹FByz|c���jz�����Ψ�.DV����4��8�3e��ǐ�H�2wAP#���}�!h�	 wFݲ쮆y<,dd�+ ����c��t�V����@��I�䂃N{뛵sJ���� �W��wy-�8�3��	Qz�1� �1�.�&��!�V߹u=E��}�u���X~,x.ƪ���.���ʹp�;�e>�O�q|#���\����"8�8�F�ƹy��X:�S��B�w����s���Ο<�=�}�{h�!�~��`[���v���M�+l��y�e]�k~�����_�g�/-�^	p��'�w8|g�0-�:�Տ0��Y� @�����VJ~��_�h=@U�Sn�0e���=��b�¬�Js���%��������D�ɜ��v%t�����?2w|��8u��1L�p&ƭ��{��t�ۙ�P�{h�+ӟ2�W�x�^�9_�����'��SJ�4�`�n�� (����ˏ~�Gǋw߻|�2]��\Ǵ�v���"���v��,(�N����9ՍR��){�h���2�I��Cp����8Q�?��N���r�4gu�ߑ����a`���X���@���I�8P�� �~�>Nro�ws�$���@�d�߮�$p��u>�LY�2b�����-p���ըµA�zp�x�Sήm�>�6ծ��6��������v����$ ����S��3<y'�q��j�9yx9���V����m�w�B���^��6���ރ�{_x����o��p[�����љs�,��_^$���Z��Doo�;<�N��A�o�:p�������)����3�����൮�=*<�<?�X�k�߇nom��p/��:¼NN_g�NN�Yڋ��F��c�8����\�}�=���y�4�>ܻ���ӣ��e��?���ȟ��n�ە�5`wa>d3��>:��5d1{p)�?����溡�"�!��=C��$>��M��� ���Ó�A�>��f���
c��$�XG�Ь ,C[��O�� 8�i�<���|�<K��v��U��CI���;~�S���g~���o�R��<2<z�+8~��o~�o���������/>���ޮ�kّ��>M5�1oF<U�L����3��{TJ�)��ң����ߢ���WU ���Z�S���`�Jv�ۻ���K�C�x]����'��J�08���Y^亀rc�� #Պ�`kO�9�e`@�呂��$�(�pқ ���q���u��yz�}�-�����Ը:�����T�}!��{9Qf[����]�N�Fx��7 ����m�w�:?�u~����ۮ��7���7�`�6xˠ����Z��տ˩e867I�ZB�vu��3��ٛ�e�@b�~�Ae�Sw��@%�'	w0�?Qrr�Å���6�����*,`��w�9%�k��<��ܝ8����DG��ċ���$���/���\���~��Ο�ӟ��޻�>8\�/�����	�������������?��}�[?�ſ�w�ǟ��+~�i~��as���Z�����@�,b��N��nw�0*�$�'F�)�\�����Z�l��2�6�w��� ��d�&�&0��5KԚ��e��@n����e�|�q��q.���R�BL���Ա_\��[�sO��Ω�\\�S�]�p����S���؏��s�z�	���t�[�C���M�~�<i��=�e�?6�ۧǢ���Ǆ���c���H'��Lxx
�����}�~����_|��󧁻��m_�o�޿����+�:��9�k���w��2*[0@JӾ|t�3�T�����ߦi�&�>����|�>X��*�ݧ�����K�>���'��޷��b��Z:��A5���X�2���ss��!N��~���$�ĮD�W���.�I�\�ynGfk�����|�g����7������bz������I�S�`�6X�G �b\W��̇����~����?������?>}5���2}1�!���A�N�7���}'YKc����D���pU�>���c/��Ιɂ�<�v0Uh����>ϝ�C��L��c�3u&B�/3�B�V�����/f��x�F�ݤ�w4@�O�����eB��O��B��{I�x{�����V���O|��њ+~��=v�)x�9{������%<j;]��'^���3�׽��b<8+egzbx��:ٱ׽��ү=T�ڗ��=S�-8�
O�zk���_�r�Y�
<C����m�����Ro�}�w�׉����&��k��e�di��u ����0��=�Jh sNyq�_� �w}�	�эS�C
������!��4�ʮv�Lp����⼯��0R�ٞ�4?��z�.Տ�����>��ز>k������S�CS�#��!y
��\@�J������I/�W^~�_�틔���?�*pH�ˬ�n����S\�.�`.���3]�������qu��S�5*O'�E��ȷ߲K�»S#�&��b:�B���J �$�k���Rxn�Y�ۃ
�� D۵�,@\N�N�}������8��[)���U�������H�(�q]�eHX���~�,�l��l��l��l��l��l���|ÿ������˝�-N��!��"���aޛ�r�.�E�;�yʟ��E���I)��,x-�A$]���UvxY|YŲ�3!$=Dj���W��^z�L�W�.�]�(��~B��͑��\O p��v��w�����/��/�?y�eK�n��sO�ң��9�)O��/�^g�5�
|�[�s��:����ɣ�zLVH,�pu "�<K�S�3�E�͔C�f�Ԁ�I�D�T��	�ȈŦ'�S�BQd�3�e3�^	��E�N��zV�3f�w�x��X��b|��n;֧��m�xH��u�1��S�W�e^�9<u�V�j�1�_��ӹ���曰V��ˉ�O�{��P<��$'�tx����K�{��E���{n�J�s�x�����:��	���p_y���q�o��m=m���_�u~ø����/\� F��u����`qr��W��am1�e�1��Dh��B���_�΂�|J�n�X�f�S�8�Y�	����_bPA	W[�S�p<ک��?+_U���d���K�S~��U�_���x�8�/���z�il��Ix� ��.qO�����˿�3��_��?�����>ϗ�ij�����}�ӾSn^�IN�#l��st�ϝᛀ��T>��7w�kt���<\7c+�6���e��N&�Z�{�d&y��G�@A$@�����`�R8��]�48+i�)Xc���D��X:�l�n�\���k}B��ѕ]P���o*���I�<>Z)s]M� �}�'����<?�np��9�?��kc@�c9=���K?΀�v��/o=<���-�7V�&��C��'�Ҹ�0�g]���k�y$+�U5Vsk���~�٭ߗw���N�j��oy8�sk�Ӽ�K�ڥ
�l]O��s������KwZ��D�#��m���s�?���F�����7g��9c�/bO���N����Y�7T�<�:x�}����6x-�\i�5��F�����a7C���e�y؁�P|F)�&������쮥�g�;]���7�)��h�Sl�)�nW�ñegF:)W�Dq߼����Ғ���{�+�M��Q�����v%�dm!`�9v_�G�?~�����;���~�w���ŋW�i�6��x� ��|����o���~��~�w��.M��!����n��Y��]�I���Q�cO��'�%u?N��չ�|�mtG{�uR��*c�8����:�JlX��s���8��ЫLpt�4MmV�R�g
�iPV���ʫ�[��܏xQ�=fǉ�l�D|8n�����^�JA����`�6�`�6�`�6�`�6�`�6�`�NQ�aA��B�ꭄ�Wn��T�>��!�E�E}Á�<[�^��$O��5�s��#��=����R*���͙4��gփ�%Iow��k�є^��>��>���������Z��>�e�V�Ҡ����K���~�_�����?��'_�����W���z������ ��o��������'���W��7�<����\��+&v�(����K	����S{6��F,VQ�?%D��d}��{Q��?�b���_)t���=z�������to�}�8{]�޵�MKǺ8���o\ 3�8�c:����u���Qg<���hAA��z¼x��<#CǱgs�Y��5ܶ��!\wD�T����~�3�@�|�gO���No��mˏ�:�`N��.����N�������8wr}ܧw��߷u~Ν�si�sp_yw����n���7���sy�c��q_Z:�k�����r�i����&��p_n��nm<�u~.l����<wy������`��<���w d�O���1�"�k�\�(���(��B���M�:��@=d���d�z�7V��f�8+�����$���}��<ﵯ�tOO3ܱ�@�� �\<�bّ�Ė�(WE��|����XrE�%��� AD�`H1&�0��LOw��ޞ�9gWeW�ZU�j_N��9�<o������w��U��Z�8��{|��#+D��� �a�~k�i�~ʣ o%���GY34�ԉ��)@:��.o�>l���l��.OƸR+%h���|[nϞ�w_���������ď���*�U����GFFFF��= ��.�W��5g7wo�ͽ������HxsC�+ �E��@���ּ4���-ͽB�'�Q�n��)��>�F�D�uʂ�jgYF߸g�n������1�.'6��3I�<��� �8��G��L��b��`O-����4�6Ń��d�d�	;��'6O"������FJN������z��@�ձ�#h�=�}����@%�I�D�Kl-K��cI����_{�7~0��M��' c��������$�%�Z��"��Y<�������s�F}S�ɀ�@��r?�������{s��	���yJ�]q���}����c��|u��{%�ɴ#�WJ=���QZ��d�����ј�׭j�p��M��6ۓ���S��ii6{���<����C�?�t�}zo]��� |�%ql��j�C~$!�������B̡����q&�1�A"\��W F�8�[�����y���gd�x�?���g�W�?V�&��
%XY(�㢸��Ջ���ŧ���5c7c�'0����8&fW x������L%�a1�}�s+�Q��
�M:-*oFO	����Ir���_��Z��y؊s �K�qE�ܝC��(���q�R	z<��jx���x���d`蘀 �gn�	���Y;���D}���b����9}O�^��F�" ������.��~a3&Ź�U�~�)A���w�r�����/��qcd��{a�Zx�z��W8p?_jWi����4���8��ET���|�6����ա�X98w~���χ<��~���|�~���O�#��}=��h��yJ���p��%�鴑�ޒbb����=g����*���\��m�ͪ?\Ӻ�?�{�a��b/�1��q܇.�#����q��\�&ѵ�a��8�_ �a�^����

� `���*D������~B'*�3�d�#B�g�m@���U��l��۟�o����JC�����?##�s+ (�&�gp�{�x�����o/w�u�>�� �����O*�����#�n�<m�ز>�����EC ��	pw�C,�/�� �.3G ࠠ�� "�{��e�¬�@��U�K�D�|�0���'c�L,(w����Y:M���cE	��4���x�����26�C��SA�q^���S�워���;����SoSwkY���\�ه�����J{��0�L/�2D�;8�~��a����G��s�M�ۗ΋&� ���`����yF
r??��+)}0�O�>;�?��gdddddPp�isH~�0���8�o�g��و�8���>*	p0�T�hf�mr<r��� ��p�����BX�F0V��8h�A�ŉR�bHdo�S�|q鯬W�4�I9��l�:�ز�z��U���zywG|l+�ŵ�g��)3222:0��
��߸��o��'_��w_n/7g��*Υ�����	ntw�	O׉r�����,�'�i<�&�j��U:JOTB��xm���>�y��9rÙ2I�$���h��c���b]n�i�.ԟ�<�02������������� '�u��іKv��w�n��8�F��w'��Н)��ԻTb�Wް�(#-�%��������.�5�AK?_����!��1h��޺~���N����"�����q�/^n�=�H���}�q9���sN?ћ�_z�>��<O�
2�4h���z�Y�~�/�z�Tzu�����e�3�zH2����w��%ѥ+�g�P��������4��ޡݑ p��,-\~Bޣ���j(5�bKHK�[���f��;��ru�����]]��WeYް� �����{ �ѝ��՟���=u�����s?���-�>�G$�E0p���u-U 7����������Iv&A;,���w�0�H�c��7g�0B|�=��َ�,��&͔SZ�k�A�I�[3��=L�g�BBc*�Y��6�i���<�F^� ��rØ��>O�,]k�����|�u2e��k��K�3����-��h����$%x�6k���R�ɱ�q̾v�y*���U���y�w"���������9bh=�ƯIԷpzv�ԉ��q�F{�d,�Z�e�F����/�ԁ�\d?��=��ϗ:�xX�ړ�u�|$�Ut�?�t͇�+�0��j$��(G��w�Ix���J H�1(��`�h�I�)��,L����F`޲��kJ�#��U�
X������BI	�L��ks]��?��
�7k�@�m��_��O^�������d {q j�Z]^�?����/�����w<���\�];��^���� ���F�z��f�(
eg��,.
"D��<�<*�.X�ݾ
Ҡ�����a�tD��� ��F<���Y�K}j1��Y8���6[�S�����)�wP��k��<����iޣ+�CC��,�q '������������M��kӦ�)�U K��{S5%;�:t[Ro',������9e\C�̘u�\�\�|O�GS\s���C����iBj:��;ޤ���J�͙>o��Wf���T�������Z�M7~&��~��~>)�c*=�����1��K�K�r���0,U�&�ϓ�����'��v~��&�M�� ����p�§�<q��<;?L�|J'��,�]Y�+�}��PӦmHyM�E�Y�w*�)Zq����T�?���@�L� ������G������y��Wo�뻿����B����-�
 {0�@%�*٦�?R�y�_�y����w
����c8r#lw����d�g*@��ZJ�9��eG!�V���#���M�㙀�&F�Q%J��a��t=i/�y ��8��gR���{M>���d�O�w}Rw#�á֠;φ��o#���=���������������������������"}-��sa��K@A��$��[b�n�E�S3�G^�14nD� ��#B^�������/=X�kNE ���6gM�#�hD�U�vg	D<��>��LV?�ܕR7�P7j�vl���¬
 
��J��nv�{��s?���v}Ul��.�p�׸Z�Z^`Y��_u�3�h�=kE������]��Ƙ�������j_:���a!P������@�fd3\����% �K��X�M���h������mh�4^���x��>H�z���1`4OT3����?�퍀�\:��6%�]
��I�� IQ!e�4"����ƯmH�gZ�)�t�i�%Y8ƘϘ�j����������o#�~ē뤌�>�� ���Z-��U�W�.χ��Z�ۼ�hK"��q��fO�MbXm�=��I	�^�%�i��1O\c���D�I���b�T�uܐ�K��|��}�s?�*�e!��t���t������݊v�Z?�8��o�x�:�<5c���W$&�;9<���_�Sk3�E��C0O?�~�?6��{U+��[W�kq8�_n�?��aM��	��5���g8<��x]n ڱj)��<Ae���?H@a ꯔ��
�9�[y)�u�W�/q�o���:]]�ܖ�� ps]�VlWް��R�[�k� '�S222��C�7���?��{�_~�_}͓�;[��v�.�u!�=�d��<y�]�(��ڊ\���v�SN����+�%�EQ�����t@��9����y!��r��O9�����K�}W�u4)�V�~p���Ahx�U���󈺖^H�32�z�8�(-� ����A[-�{M�.A^����.�<���>qj�U�|Oy��'ƶ�!���u4d�v�no곇ޣ��|�Xz���\'�E~7�p��6/r�urۑ��p�j��~������1�a����s���QP�&W���)����u�!�� ���{��� Q6��G��&��1ޡ�Bķ`]h�Da���0��A�gG�7B>��+9�1�E �o��x#����g��o�����o�����Oܹ�أs�^ٱ|@FFF�V В��^ɻ������.�7oo����L�9��h8UB38j�h��� �p��'�����M(z^�~P��a,Io�=
)t���v$6����Qe��)�.YX���O�#���.�� �F��z_��T���mIb���<���5E�;m�}lI_6%u��]^�9_>[�Z9T�Wv6�e_H��R�SC_�7|K����<=�1;թ����n+��;���nxǯq��ydr������~z�~>&�S{�qJ�<|�E��n�K��q�������;o���a���)�U��8�ҸIL�v����o��\#��9м�[��E˄X+~���?��F�X`�	t�F��(0�l�ry`���%�$]F���(�(q�E�#�c�K�z�6���#��f�g�6���5X�}kD��H��bs��g����'�������z�(޸{�.����XFFFF�@<�zr�������%�+ϵ_�m!�F����L9A�t��>)m�֨B���p��,x����B���)�d���Ù�Q]p�^&ϠIf�u�l�t@	:+н��~��"ʗ�>�`:�/�fG���T������u��z�~r�#pLm��%L��� �<&����M;�l�}��#!�����H�8O	�s-�2; �ۺR]�{K�v���kRF��Ϥ8t?OI�P�|�mi�$5oc� ƶ��u3��:6���t??%nc;��<������|�r��v��~~\�2Ę�u�2�:�bL��{�h.cd��A�5㸕�o���P�.�0�X��7b__�'QO]c�,�JW?���B���w.��i6�K=s�M.c�ܚgr���.�) y��<F�q��g��0΋ �T^� 9� ��~�=we�j3bţ��s����O��O��� ��.�����ޣ��>��_��������*�����сCx ����`�\I�V�R�k�+�Jt�m �(�6X�ڞ�㴮`d�e%<^@`@����".^@S@ɒ��݊`���p�\2P<� �� �(1��Jg<0) �L(���`p�Aڱ�|h=���䍀����m����ug�����r�bF`�Iw�^T[N}_u��O,�>��O��O=e���5U���y���������{a�|����\m����7ݩ1���1�=4��N���O������χ>�������χ�ejܦ~�7ޱy2�_�����ߌ� ��aXj�-5_5���&Ğ���b��zŷ���i���A|j��(f	x� ����	m&�xH�%�Ai����`0*�c�1�<��p'�[�b5/�C����>�e�"�ޜ�w�[�R�qL���x���i�R�F񂳭�
v��gg�|�k���;?Jsm^#####��
 F����7޼y����y]j� �����sB���P�,$ �^����l�Hw�*���'$9x�J�5Aҳ���`��4-#�U�ܴ��PR��(�� ��HF�Y܇d{�˰�<�3Ts�\��^�:��XW4޸�����x�~���MCV�z*�l��r��wJ������0�U�8�w���PHM/O!�1uݤ��9d�m�s"\�Mϒ��|��ؾ�%���#�������O���#��1��ű����p
y�ȸ�8D��<�Q�~�_��^�-����p��Š\\6k=������z��ȍ�����M�g@�O҆#�� ��X>_¥��<$!��P���X~o,���A_�����R�J:��d�  ��IDAT�U�cgB���[꛾�;�*\�ح\�eddL�C( �o������̷?��w>���UyS�Y�;�d�\���c�m���^��e���j"�mr8�h�ވi.����@1'� ����4�I�if���
�(5ب� P�Ee#���&B�Z�׭���b���>o�z�l�?��z��0^��*sH_S�{�<L�E΃�"�����%�!q�H�e�u�9�\/�����x�3cTU-�L�3Z��r���A���g��9�T���a�(Gj���2%Ƥ?�}L�|��5r#�'�C��� ��u��@�����!�'UV����K?���>3��A\���mYIK�o?��������y��Jz�-M��Ǿ���<9�Ư����0�s,`���n84���"��4�x�R�����ˤ-� �m����r-H|��|ٰV���R;~���a�O����s�u���D�<�]�kN%>��qE������e�]FI��@�q����G�a�b�{ܧa�F��]��
ēp��?c�ܖ?��c�4����II����cw��杷w��m?p�.�����yu����]�[@C�VW�O�������;?�/��7\�T�;/
���Y'��̑�80yW��C�@��dq�O�}$��15f`��0���]�W_K��
��"߸g!��u�LZ� �B2��2���5�ċ@�@���~?l�Z|����~�4|mu`S��J�!��1s�S�߱s�!�c�S��b�2�ŕ�0UGo���cA%�;t����c�ݡ�z�>?4��$!c��R0V�[�$)�j����y���������Ԁ�O�͍��gdddd� �{����Ȟ�rބk�"/B��c�c��(���Q�!t�o�ށ�q���K�qI����J �>*8������o���(0ƫ���F�9�
�����[��;<6�,�SlY��u�c�9+��<���o��g����n��b��fU �H�(�������_y���;���_���_�y���}�+: �%�ϸG�tu��Y�3F,�U�^4Ӏ�G!��!� ��N	9��U��4g����6��q.^0���W�{�j����1��D������Y�s ֽ��s���0?�5�B�6-�~^-u-Xs�32222222222222222222222�#�uo ��ӓ���%��}�P�<FH|�բW6bm�s�|��xj+�����g�}G�{���=�^�ѫ4z���QN	�J�D30�q5�/��wAJ�D��=��L�ɶ��������={����gB<�s��5�
 {p l���
���|���R7��G�W��,��'Z�[o�.�V!��ߜ�~��Z@KP*(KcE%���r�]�o���B1&�Y-:o��8��5pao�.�/C%�\���?�g���f��Y  UӰ�0L?<K�� M�E�v5��L��E��?��]q���q�8�T��^��~\t�c�,XA<<�4��j�j�Nz�c�x�ђ�Yҋ����a��?����7�x~4T�є��|�d����&�ί|�So����RԆxׅ�6:UIar���:Hr3<G?o�I�G��Ϗ	��u�{�.�1w���ZpȳImqL�l|[\�8jyOSv�[�}���k�)�~~�j���y>��t�~>��{n��sL?��0G?gi[�x�c9��/�����-����r�I�]��0v����O��-o�F{�p�\a�?�Ξ1-�&�]s��)� s���|O�K$�4� W��*��	�nip� �p��I�X��5!o�O�����P (�d^i(R1��֋�M�;�D�	�=D�!�������qI��Y�/�f��ro��=�����Կ��H�����1v҂,##� 8� {�ar�;���_��x��V�*# =����~�e�%��e9�_�]�_�a�=hh���w#�!�`H~�8c-��4�ᠢ���/x�<�\�4���3 l���������Ð��t�`.}B4�Qx�L�|ғ����k��B�Ċ�f������������������������������{�d�ws�>?�� A���tG��0�>Z�c(o��|l}�bi����E(
�?�4G	��9�I~�9�E��56iܢ�iF��3^�sX�kEa3��Rް�x���Z����R!###��P ��O�Ϟ�\��k����7wWwo䥐Z�	8{�ʆ�x�
>��eԐBaY�<��,��G�+$��u�7b���r�Ϲ������ü�ڄ�<�y)�J����E>j@ZF�+UQC����P�gP�m�X�~�`�ާo�������Q�*/��e��	
�P��0}��>���k����{���!ϷŕR?��6&|fj�	c��|�w5e�������t�~>�S��c��1WL��c�O��c��6L)���=�XYG�����~>����w?߷�j>�t��<������}0����Tx� 6�B�5>Kx���i[���K��U=�M�D�J�c�~G��VAG!c�:�<=;�T�e>p.��*���!h�8X��G �.Q ��lãjTP@�
�G�A(�]���R��Nrvnt#�_> ##��* (�A�]m������o��o���=7Wo�]��F-��w=�#�y�9���� GQCt֚��3�P�r���,0�,�1=���p&Ҝe;�f�����Q,\G�4�);����9��`�����8=:1�J^����h{�0�X%?X�"A:ȃ)>ƺ6�R6IZ�9d�n�n̈́3���e{��i�ݥ��d���%4�.��h��������> �~���a8��8.��=4�%5��)�8��"x�x��9}kRѷ��N�KC�gdc�}�f=�����]�,����^����t�c����;�1w?�+����Ǡ�M�)�)U¯��.�G���|H�R��C^������GlsG^���I:�`�2����;=p@=�a�>|�ڟ�C����w�c�_�=��]iJ�"]�L'G�����ɷ��̄�D���s��g��9������wz&�j��+�+P6���Ix$cx��R��UL�e�)�#xU�����n��v�g��4Ju5(=��x d�Tl��]�$�>�tJ}�dO������_�����x�������3�V{�2222:0� -���N���_��7���߼�{RI^*ɑ\G��T(r�-���ְ$�w���]I�p���=]�;+sO����jWF�Ki�)���Y�5{�pr�<��'�&�h	#�*��D0��1���@b���d�+�!O����m�x|zX��ҟ�Ժ�柹������<�=.q�x�[����,d� ��]R]�]��S�c6� 8t=/�R���Ǵ��.�OC�OR��R��)�K�v��9G��"��y�?��s?������S��fdddd���*�F������s<��!�rĸ��LRS�F/0;.�r�B6�g�G���=��l�|y%��Ps_X��R�h������WM���0GKY�J9�	cA�ھVUyح����/��+�����˿�<������ �� ddd��G ��{��/=}��*_S�<ߖ;�5��
#0��_?܄�h��.����������` B�*�YM.�_��na8h�W�|�`5��/�{������K�B������FW�^�`��f�G$<^��0�a�1��fz]y@�똗&E_��9��]�Q��mc�3L��8��m�09��[7Þ�	a���t��_ܖ��c}�BJ��*��)iv��}��l���?�ݎ�G͕�ظn�88f?K����]��|>,1OS��|H=��}c���χ�7e��2�%������ۀc��#���4̐,%�!a�|�'�x�y�{.������,�.�#�i���h\ȸ�a�2 �l����A#od=
��gQ��FA@qC�3s�g�{2�7	/�O<򠩞�~���E�p��z�b�ͮzX+=.W��y���_}�ǯ����?�#�}P=~U���!������p 쏾��B��3Y���r+4��Pb���p?"�����Z<�d�s�����9���	`�j���/��K� M�f�^�@�l�����i�h�c�>B���V����ppI��Ao����nߥFM4����*t�xG�`�F^�>��cc���A��%���K߸��n�eD�2:�W��ER�P�����c�Xˎ���Y�;Hn�3	����!�r��p�~��1Ͳ�K������9Өs?�ƭ����HN�"CҞ{!vl-±u2"�(5�81��S].I��~�L��)7_����F��6/�QJ$C|�3��"&��|���0����Ӕ���54g�=;E�	��hL�x�V�)�% ��;:�gY7Ro�g �N�x����2��Tw��E��W\����7?qv�yq�,����@̭ `$�'_�x���_�~��h��F(-�vL�0�UZ�y�om��|$��w�±����5��`����S2 ���Dq.���[RRO�1��7F���P�ϰ�AP��oB���$�g�� �u�@�c�)w?}��x��}���b��@;.��՘�xxݕ��������x�@eu^�ddm��#v�,22&�1�y�B,��22���#�?t��)����M�M�p;���%�e,��O�N��=�n2yHy���}�EX��~������� ��h\Yc̱�&��y�G+�M���U��yw�����3I�g&iY��G�����P̥��s<ʚ���=��D%	�[��x�TlUe���0�a��+/�O}�3�s��u����]8� �O|��G�����?�����噑�\
-Ñ�V�m�y5��u{�A��U�Mc����>��(h�(�����̘@��Od�Q����_Q� �4�~D����	�� g~0b��1u�cHM3�*�
��G%J�����I�̿���A�����h���s�,�Ɠ���Y���A=d�5O[���c��pLǤ}
u;%RʛZ'u����K!�뙥��)�1C�U�r\g<s�sƋ�����p��>�>��xs������wL�#�4q���Fn�ܼA�Ƅ�C!����J�H@�#Sq��<�
x��x��f���r�`�%�	��9��w�<Cˠ.� q�ly���]Al�
ÐI�'U��?W��s}-_������_�9��w]��MA�2222:p ��J\����/���[�<���}�Zߨ+C�K��ﴽ����/J����_oIt�p�"���,�t$�����P��%��A��X�@����J����/
} ��q���;�hE�K��mXQ=t���[S�lW]�m�@�Kֆx 	��@������@K�q���b>:���zp��:8@����\��i?��1׺i^
f�e�"��U]wR��M:i�����:ٗ�!0������&*��{�;���m��*o��R�j����TG���6׏���h��>���2&x����$O���=�0�w>�c�ܳB��{m�;e�J��}dÐ4���7�����lk0U�q�jl)�H;���@C�w��ef��J�����[��op?o���|_6x|!1�T�}L?Wm�T��/M϶����+s1bn���4����m"��v����~l?�^�Vr{�0U�����0L�v�T����H#�s���X��>3u�O�o�@6E<���$T����>��Zҝ��gj�g����hc��m����%����'�δ���w�'��>�s1ǖ�?�s�	G�XDRJ�����&���s�<�5��ҏ��/PJ&V����6�af�Ф��i'���X���I?/�,0ePT0@�P�': �KϥCT[?eX(F�Dk�|4�#Gp(�x���e���7�3��<:���]Q�3y�^}|�|�������z͟m/�׌�v�(###�ͬ �]�h��g7g���������~�w��߼��B��p;x(f�����SPj���Na@�#��������|�~p'�^��睿B�c@tkc˩�M,�M�eM�ԭ�w,ǘ�{�}���ԉ?�&.;��i�j��p ����@ik�`��[ :�~�8�}�r�4���x��g'Øt�<;��SktMi�J�+p[~Xz�mC�<�d3�AÎo�w�~@zC�L��شe�^��y�3�|�#�U�)�oF�{�(e����~޷��-S�|�un��y�ʂ�K��ˁ!m�'Z�
M��!����q�~��׷x�'���~�E����k_���r%BJ����z�phS���#�]kz��iˋ5����%���aM��5������ޔ�'��0�m����C����������pl��$p+q~0�&�J�$5�����K�
q���?�g��V�x~��߰� �����8@�e�����W_�h'����L^�-���$[��L�9�Z��H��25�<�\�sO^S�w�g���y���Ϳ�����4��fUx
��j�B�4�&HʖY�+�@�1pa�6{�e���AI���Z^Ox�@��<�\�Y=ĺ?�����䥏���d�k���ЄN��p�O�bL������:�ܒw��o����=@�Ǧw,2��'a�l�35i���>G����ōr$j5)�2���)
V��&�R>����}u���fh aY`�i$QƤ=���^���9Yڜ���L�V'{�u�|-��e�H��p"p��ذ�9�3c��3�k�~0ǰ6Y;a^N��'A;��w@��=y��y[a;*���,�O��l�:!����Zи��0���u؞4�����a�,w�O�9�Ly������e�(�ګ���'a�i̘�g)���zg�v��NP��,\O}�h8R�����G�zشkHn{�L�o&��Y��@h�t��K̇`��.9�G��3#�Fa�v@����ʃ��i �&2k_��T4�;�w��1 �ꕏ�y����mpV|P���/�a:rFF�	�
 Z��R��;�}e���9�º�7n�U���F�����P�wоB9���<B�U�0���^����(���\|tB�����ߧ�|����>(1_K7L�Ib��PFs-�$��K��P�5,A���:���gj���$�?1޾�+���d����ܑ�=[�n"��u(L�[���T�<{�����)�X �m/p��@�n3z����9�̲`�^��N�T�iPFp�(��J�̻2��Ƀ�͚:��^�"�W�\�넑�d]�e�x��f���R�L^'�@�|߭o�u��CB#��~�[�i�kƘ�v���ɾ*��*	�z'#���S�z��=�^L���h/㘠d}��� B�����+@�_¼����!��?7pq�q�'!��4B���ވT�����WD�E������M�z=X���`�eSA]qmY*���������Fqu�2������Y �r������W����f��\�;�
��ǝF.'� #�S
>��}��� ��`��*B�;e ;X8ǆ�S1�0 ��]~��S�
V��Z����Q<�xe��}�@<�6��hU�4@� \����b� �e�[W^���c��^�`��Q�d#�!�"�~���f��I��I�� �,𚑑�>J{JAY�$��T^t�{��S�^F�c�dBod0�@�v@��t��=,dh�q��[^�וSZ��:�
8Ιp����d�۾p�N�\�
Y�\�Àr�P����s���v)�u����L����3�ŵB��u+��>#�aD���TV�U�����V����j����sՎ�y>;����+wh��\vp��m#�Hֶ����#��l��<UF��	�������� P.�޶1-4�t|Kl���['���n�><�
�] �O�F�y�>���c�)(O$��-T�d�'����)e`y��6�+Y)Kv-��+O�����f����r3���؋Cx �v{�������w~�K����x����z�MCJ}j>W&\�r�������>=$������z�׍��q7�����-��A�D�5nȣ 2p�!&�C2��o:�k��8\<xן	A5��8~�î�y]Q�uս��3�6��:�T[���!����V֑HR��&΂l��F�2>.��s����4�g����A�����+�-ߡATϪ1�V���VC��~��W�6�.L�Wqb괒JK? M`��(AZ�[n��Ŗ����e�u�p|�Z���_}�9�e!���/�������0��@2�7��`�;X�x�s��bq q#��CS9�,됸� ]��o��I3�b��
��pCZ�LҦ���}R6��\A�r RȜ�v;��]J?T����79�f%�C��	Ǩ����i�{�����T��,��̅����dl5s.�F�n�PE �W��l�r�����S��S���o����Q`�W�FK�^�@hDz���eoØ�K��e��A��
>��c�c��T��+�~��������-b���#��^S�8G�sΩ���Z��}��f�Q����6���6!o��"�j⒞p���ƁL�wχ}�y/�g������Ҁ���Q�n��¢�x}a�1�Xo~�>��XT;��gU��z��~�'��������|����g�z�����[@K�b#������W|�-��՞Je�;ʟ�p�ϓG���GaI�e�x��V���1�	q�bg~@�np	�Q^�1DY��JB��̊Q{L�	(5���)%)�/[������; 
�1����@o��k�Z��.���G��),ԏh-��xx��n�dK�d�5���&X��=sO�b��YF�܊(������2��dx	X��[w���%�g��?ȅ y]�
S����)�����)��A/(�h$u�RP��^Sag=����m\�����~��g:�,�v���b�u������YH���z�s�T8~�XOVs]wD�< �Ke�],#�Y'pR�����r�nw�=��,`X�*�_]�ۜY��:A���Փ�
�nn��0���d��#Ľ!��׶,��$й,:C�%��`� dun�i���sY�v�/���"3g�+�P���Y�������c��
��kqZ!�r,��o`z!T cLx6N
�@�K�C�]W)Ga+��"@�bX��)��1�SX���[x�./��+_�����?�����×���/�߿�2222:p ���q�����} �<��]%��f97;"Z�
 �����M$���ʸ��J H<s*4��QE��a�w��[>�N���[,�ݾ��H4=������( ,D�6 =ǒ��{Ժ�+ĚfnzN�ˋniS'B�� ��>,��M���c�������*o��Aj~�ܥn����aW��\1xZ4=�DA=�F委s���P>HQo�
LXkjD5n��Ha�yvঈTna��{Q�v��ᆩW��!�^�Ω;Za����r���*��~`�$ZX|��؊��-Mc�4�6��F�2�B#Bۨ!O`a?�2�,|�,y� 3SL�&�\�t]��iʲ�k��G�#��$��$�X�K�������<	�2��ΚH�@��в�nK?��N`h���n�V�ι�Qo}��)���<�YE�/ha�B���#����Ć�|��Yk�����7nL�<� �ĝ�:�cU���;y5�^�0���{����܏�rk�c� `̊c@K�F�����0��1��zk
�G�t���,�t���L�^��H���򚃛����\����0C��qF��&�?�4�?#o��b���|���#����xG�Z�>X�eg���U��{nv|�!`򈆦���fJ�[�*C��y��sOʥ�u�s_0��wU�r�oH�����fu#��{~�����ۿu�ӟ�z����:###�� ������W��X񫒯+!^�k��ٍ(�p6�|  �p$�_"� FH����ߚ�*ϋdz挽g�`���
��2>�<�4����:�I��R�{p���G��,��	֑W��t���q��@�68S�>�)�+V~we�JW~����Δ�n�0���ps��/c?T���4JE�2�ko$/&s����Oъm�(�mT󥃬�_d��[���C�~��ȁ\���+�pO��J��~����mi ����/P1���F=�k:��m��V`���s���R�g�\�=�F{���w�����3�pk�����țà<�H�/��m��y� ���.��{���']ƀ��}�*{�d��&d_��Y�y`y\���x��q���N@���
m�ՂA8������P)&V8pܒ�:��<ߤ�m\41�+o�Vl�[�={�7Ϊ�4�'��m�f���� ̭ `�1��������/]}����O7r��-5i\����Ds��}�U*A��"�3
qL�
Z��i��q��r�
}����	j�[���c	�৛d&]JrCN�+"xY�aڝˊ�aLh�1c�hݗ)p�H�&�B0:�����������(r=�����l$����{��ƣ�"�q9���nN�4Ք2#^6����ɑ�t,�rhj�%�s���T=�
����hI�1�"'C�&I@���:W� �J�)՛_AO$VX�ׁ�w4��	���	�1 j���F�}ۼ�qDP� ����4l]	 hxGlX�+T�B�J��>����j6��?���I�U�d�S$��旃Y��esdt�q�'i�2f�"��P���q�5B���R���r�iN#W"]]Q�Θ��r �L>�����hs�hY])%�]	���ۿ�{w��߾���X��{p��㯽z����G?x����/7Ͽ�r%�Y%�vZ�
�Ҥ  )��1��3$�&�F�:z�
0�%�L'�9<���eh����@�B�P�<�Xs���� ,(����T^�yg�neςOO܇���}L��5�B.���|�2������#���k����<~f�NĊS��
�]�f����j���v�,)OUí�l{�m@����75r���g@��/##��#�<���#�Rs �*�D�3"�����je�`����>['�ylN���}6_) Ϊ�<�\�t�c/ ����N���}j� EB�@I 0:�ֆ��A�PmL)ei�Iw�$��Ɩ�a9�E�9<1UQYc^&V���$I�)ઘ��J�w��7������{~qq�l��^ݹs����]�[@C�_������}�G����~᧿i�`'�+坡)D'�#�J�6����} 摬�ಟF�c���P�@Y���+~��e�i��w��`�cM�h��l�r�4a��ME��-3*�yǢ�j�5y�3�6�?q�� �ǣ��Ǣ��J��Dzu�wn�/��C�m�!�0f�^X��O��譢�����uz��=U{��>��q�~>`����ҴNͲ���N��T+����i�y~�hS� �P���R�v�|������X,�~�`��Uk�=�}��T����x��ΔX�ڀ��qoǮ�C`����ֆ>��i��;�M�Sm���7~ݏ��C�§Z�]�1���ujj}�U��e4�9P|C��E�2�9	b�x͢^�qX��"߹�W5. �ߏ�@FC�&���m�(q�<�` N���^ 8E7X�7��䭝&���i&�[��ce�q��CQ���Գ�l~��c,wuV����~߷�ɧw��'gB\޹wo�����Ȉ0���@� 7��%/���Oߟ��/����_*��7v�Q��9��������rZ�� �.��A��a	x�}�?w;�~WD��Z�a�K��2Hs����k�5�Fc��f*P,����2�u�M���31�{�u�u�������3}����̷u�����xR'�s ��ǌœ��x��m#_�Luޮ��7�0��|��T�;o-]�I��Rى���c�Fp<O���M�_�q���8C�����yi�ߔx��ŧ�/�Ye�Tm+��C7a�~޻SP-�)!jӬ�D��'���RB5uκ�l0!/��v~�چVYkn��Wj�����'��>d���=TBL�dbKJj3���汙�yWV�r¼�{�ĪWVcw�N��O_�4BS��X��Axj1���㐚�J���=�(Q_�]�Ҳ�/;s���z�yA���^���:�o��ơa7��J��r_?eV�6�Y)@KM� �QD��k��m ���В^�<v:4�	O��[~��x_��)*��ʄ�plj��۫)k䮛j��C�=�9{��(E�H�74�A�1�&�bE�.n�r�y~y����ޝѳp�%Z1tu`9<ĈWg��J�=��ͨR��2�@+�֓%�̀���
�=lJUl�7��ا�V�#)�Uugǲ@FF�� �n�������s!�V��E%��jg�X1g���nP �x+(��-P�M,*L�7���Z[� A<�~t���F3���8�����uۢ��0+-�%Fk�e���
�`/Y�4���!��V����"$�I7;� �YT@`nP���B��?k�����I!@��uE]�`8�k�6��m}t�IU��Sr��2h�lLq=��xTK����=~�:��v��4
�#����F�&���k;����œB5�� X�+�5A���~ϟ��)�kK��quI��!%j�D���_��u6�r>F�uX��J�F�G!=���,��t=j�T����:���g���YB�&t��o>��x�K��W3�&�Kh�;B ��͇#��Frk�6���б�<Y�]M��RN\J��d�7R��D��_�q8�]y���x׭Ê �(렂 �*Up$�N'�B(�O�G<�� .$�~�*) �� �p�#��F���X��<x�4�S�n�S�[�����_�w\��J�f�1��֝���dD�(
q��Y�����ٗ���y�8�^�JU�sś�5JB������*���1JBSAm5AX��
Yo���8�V�tS��ņ�
:���R�]+x��3$�f��s@c}q�I�o�M[|q��wX��N*���;��Sn1׊S�7S��{N}[�-c^̵�y��w���e:D���wpk�S�����3�-��o�K��E�ٸ�2�5uc"/Ɩ�E��Cc�u{�9C����udSc��n�j{OY��ښ�EF~WÐZ��N2-�۹�~9�vۇ�џ�D�����-�Ϋ����_�(�ނ���Uw���!�!�˳3�r��1F���:4?��b�;U���������*mε��j����}���G����;^�3������h��
 �2�|�^�?����/���>.�w/�K.����;�����Y�p��S_@�3�3��-��
������"�_�76~A� �	�6c��	H�3��K���G�;*^42��Pq H�A��)]���B��h�z��@����k:��n�L�C+����L#e��+�C���!�Q�\J ����V8�����CrF�	�YD�و���Mz�A�r)#�dh���m�32^�Y�:/�,�P o���'Z�G��/d�Q`Ȼ������Ct�O�W
��Gޜk�:&�h��c��cp�QL,b�򜤫P xg �*��"҄n�?:���*ύ��?x�$�uz`\��L+w�]�J]�ֻ���ɿw���/�����\\0��mYFFFF�@</�{?����ӿ��O��!�`Ei]�G�1ݾC�'���
�?~���VPۣ��� ���d `̻�!$�sè �4���^�!ҟ�b#T.`p�wN���Q�v8�r[�w��<IY������t@� �A����ZY��7&L8�L�&/_�g`����i]u�&��ù4K�Ԯ�j�۳Nڲ�wqq��{�oYP�$���f���?�8~��3,龚U���2|^��e�=W^���{��/���M�����ukMZ=�	�Rr%���l	���+)�<�����v,hS�oV���k��r�~��ڈ��<n2�yT�D�v�/wJ
K�]K�y{��ؗT���	�fKq�mAL������[p�+�&kW聿Ȟ&���(�z���M���K��q�� λ��p�GZ�雁=Ὣ�>�H��9�`7�lZ��8!=��#�!�w��\����>�hr�<��n�������Jx��u�����,�誟Y��;�=��N(>x���KA���p�g��Z��q� �� gX����?GE�c�ia�	�Xh��>�y�ۚ<j���W�|{.Ͼ��_���ǯ������{z��������с� ���MY������Z�|����R��N���+�~V��N( .U��RY!H-�)�n���d���f7�ި�����{L1�����`w�9y���80e�y�A2�`��,��'��W$|X$J�7[���ǁ�m�E� pr/��o3�ߤD�'�-��Y&���A"�ڗ!�Ge�Hr���w��;�6@�����Q<��J��ڡ�g��H�֑6��$u�;�5)4�g�p=^̹+�ז��6O_p�k�i��'��)�5��qި�R�a�_A?oo8t>�NO��GS������-��@��V�qX��%�E�vσ��~k� �;�&t��$��>��k��@��M��@�=���;���T���l?���ᭆ����C'.�^��j��a�΃������q����)�G���)�㡡���}�T��?Vݥ��6
se�&�p�3l=�����ȼ�w�d��5����]��.�ה����=��	���/��K�7C��D�R�}�ڄ���05􆙡W�0�x�0/02�Gd�w�֕b���f�*"q#���ʕ����ѣ�Dǣ�y�p�51l�^�阥H���# y�y���`j�
~W]|���{���޽�̧>�f�edd���
 �0V���/��������C��k�J��W	Dr\+���X�Cpt�Bf��m>Z�G;��d6&�����e xaP	Έq��i��n�@+7��r¬�|j�&\�ʹ	�ue.ρ�\B�5!QӴ1��d���&W:T[-<?�i�J߁�*2�z擞�zdd���@�V(6��]:��۷�/D���<�p7?@6�J�B���*u��Rn�V�Z��a�pe����pYA[��ٌ����H��\�w�H����b��mX���=Fl�'�Bgh��y\�|\��g�0*
�/�ة��;��wJG�g0{d,�+_�̀:S��,���N8ـ�/��K��|_�M�;d��d����T8_}8瘹o�9��*8�M�+����WP'��2�a�ιo����:�1�RǮ��C��[��.	v;)��<
�'�I�ߔN�}�
���<��l��>,j?��A{�)�I��1G��}eU׻i|����%��u|��޾Gpb���Gȷƹ�[���yZ�d��p��1н�isC���{��O�=�A<zg�A%w���5�\Jck �����3�2�g��FǮ�]�� IB� �2ZN0�D���~/��.y�
����-W�ؖ�W�������4�U@FFFF�ُ �d%�>�����9+�R�Ti�nV�#J0����%�a`t�i[5���L6ɏ�eK�2<��mnK�I�7#�k�&��p�� ֌�.�=t�H�&�S�=T�-��A^C��:0N�ݏ0�ߙ�=��9�"')+�#`a���0�������p .w���8A��PÓF�DoD�n�L�U�%�JLp���,�R´Y걳��	�|̔�(8�-�l�����lP��pܨ*[`~`�ɏe3�i�M.�X�ám�%q�yh$m�Sf�����Ը��8�Iٜ|0_�,��u��A<=�ndYQɋ��Vbз�k����xq�Y�+&�<��3�[া�Ϣ�@��"9&��C6��\ I����x�JH��_���mo�W�A�?��񽷴%�Ct�,[ȓ.�J�=s��<�T�&6��")s,�#�'�`/A鹻bR�=7#���7n�6$�W��:�^�R眵恮��2�[��L�s2\�ի?1B�ܾ0���-���u�q�{G�}��=z��:��b��T�]5��t�����4��z=�˅��_�̥
BOѯBbM�#	ۮ�e�ЊŬ���*;h�	��W�>��P�ε�w�"lzj'��6�~7��`z�f=8������ǸC.�]ހj�C
�[�wƼ���M=�
�GHz[S��Ѧ���g����OQ	�uQ��͆m��U����z�;pFFF'�V 0[���uo˷���h�h{ys%�z�d����E~5D�;�G7,��W�(�/guN��c⚺��i��(a�ԕ�[��cd]���:��A�F��`z���;��� V0W�ZEv�Np��-�� �X׹Ϙ� 77M��X��HXq�^ �����n# �vv[�r�>; l���k�\�󞛟�R������$Kh]�
By9F]b�'"w���	%��x���,>�>~�o�P�s����#zcQ`�v�1>c��z� �e�֌c���OD�<8������=���
��*�C��6D�q:��|f�r^���7��t�6�)_�����^?�4�� �\d�r_�҈t�1��M]�Va?����Q�e�ٽ%�P%?��c�n��y�R^����c�1eB�����2 ��5�R�.�g�T���/
�t��~Wl�CW_���V��~=(��TP����-J�Xjr�gɇ�?���)���r2��N�Q�<Ev�
����L�m��猌��-��G��(�U�(<k��������<ݘ���9Sa$��Q 5CŦ���5i��5��Y]XTh�0A��\�i����q�P��h�IUa�|��vS�EBm�J�c᳻7�xk#��fddd4`v �'_����g�����?��}����OV;��k^�v����2�.��<�T`{+��~ڰ�Zqd"�'(g�J�8��'.]�Tl�#����	H���MX����ʐH�qמ"��`/Ɏg|QCrߖ�(<(?`�Sj�ă����w}�?�I3Eʢ�-KCDs����ۥ���Q�Z�qn;S�n�WN�eB�Ul��՟���6lnM�"�����k�N�^��Ǎ�g��l�b��cʺdv��l|�P�Z	��QQ�A��K�}%���y�waSQ�N��K�l��2���cg�5S����-�Mݖ�Z
�Y���Zx+��Z����K�)��%`�; M��e�k���)"#������юQR��M���nRkBɀ�:n�œD쿢�XY��B
�M�f�9��'-w�<�X���]0G0�݀W�%�Yӭ
�D�y3�����Q<� ���_���}o%*��`�$��!�9�U)Lwgц���\�<o����9b�Y0�r���qw(Jѯa�R�J�Z��be�O2<*g���1L��\Sg���~� r��!w���z��k�)c��ol�t@���Xf�3J�%v��@.��w���W�܄����M�Enb{��2�SY��+z�N$Z»$����@���ͼk������q���fN���䑜Q$hx��E��:V4> g���Q	>�O=�5}����&V�|�L�����HЦ%I�>��C&�h�-A1!���C�N��]�S�����~0�n��R�]w%����yP.F��#�F'aR��_�u%L_fwv?�?q�}��}��B\���6�(:edd����[�}�mo������[���ϔ+��M�Į���ܑ�TX�u��(A��B�cX� m'��"�u�F��/¦�d3"��(䑴�ݑ9�Z얠4�׬u�sf�#�D�c��J8*w=(AK뿽"׾c��O)�]���d�ާ���N]i*�T�!��ݖ0A^�{m�qK\���N�]p��}�R�K���q��,���/vټ�385�S/گ�Jv�t�n��l���̭�_|ul�L���1�M��`��`g�sO0q����H��l�Nv�߮���d��n�K�]�Z���|��v^������WV����_TN�@eM�m�t���76w��X:�����fc��[B�RpRǰ��	����^UmuS}�M<�$7�K���l��)L}�M&�����C���AdoϪ�?2,u��(g�f���-l��;6oHF�����.'�=���`�r�؜q���m̘WɌ#ˤ�eZ����4E7���+'U�s�
3�T�H5�]�F�Li���;��X?K����:۱�g;Swۭ4�'8'�c�;���@�N�����z�e������F�����x�ˀ�E���!����i��0+ �J�Hw�����^Gڹ���j���З̚\x�um�����x�H��HZ^`�\s�fװz������^Ksd�Q$�5����`l�JI��[��'Fk�Wz�^����w[	K�Ŷ�
��Q[�_i//�ΤY��\V�ݛҌ]hY�9*ފE�]]�Z��ו܅��>���Ua�>3�uJ���I����4�|S���g�Y��N���̰����Խ�'h�p�۫^�	�>�<Pq	�@{�J�
�P�oK�N�*���
,�{�QĠ$�AA�eڙ�{�+؝��0�V�	��34\/�\�Oӯ�����t.펺\j��C�q}�ېtsp��^�tLŪ���	�'x��y�����&»����+��� �u3)�$xԔ?N>Co���fz�yӌ*-*�G�z�E�$�9�q����qF�-$��i��Vl'���������L\Ƚ�kS:�ɣV�\���X�B�.��������B\<�������,+ ddd���
 ���䛒���ZȽ�����_��_�������G�kŹ׻
���X���'�>�@>QA@�2XP�@x7��)�)��6nt�oS����v`ry7�9�%�e����`���VѠ��8��.�SH��d�&�����xw�4��͎�D��M6���uE�q8t̵��E�s�PF����]�Y����vzS�dOm���;v}��bl�͐N�	�7�V�Z��E��ݓբ��oZ��sVR��ߕ�ʸ����(S<�5d�&ε\;?[�;�V��˫ꙕ��21��.0_?*B��cz#��Yɞ?���V�/��3�?;���Cͪ�������`+K��1u�7Ym��MQM���}V�W�`��Z��bj���VR��2�Uיm�z�P0�)�:dLg��֌N4n��='��Ne6��m�B�������a69�;���|!���OT8��\%%asB+]U���G�JN��wi�m��8A1��nd�mi��&�w�+�$�����Ж|gw`,9L�%�`_�9�&�6��&OUcۓ���r����xTّ�(]��:���]�Y_��j�ez�~����L�N�cy�}���Q��b~���&�r�n�ו|��9-vS 0�L�kf�����R�����9i�u��� �~v}k%���2�UU�O?*��͍���C�Uv�"�ґGt�k�>f��J�w
v����+��u.������Y�<�hE=׾|����zB+�^�N��յ�U%��1�ǖGF�V"V���{�����Tm�(�	N�LcSKk�*���j� ��zfk�+v����v��s�u5G0J�z�{m�g����MΜEgr��~�p��ٌ�`5�z�Į����F���Rә��N���z�����J�Α���
�\ua*�+df���n��.?�ZW/q���zt�h<p�f��B"%k���ͺH{��h�	�nkڰU�{$�Э�^��ێ�}�\I}a[oþ|��p_���g� !�r%�v��22�[�?s��C�4�ci8�[�ф�y��5�KT��#9��2�C��m<r3/�n�L�|��7�zRI�'�����IMFFF�G T�j���'����>�V��|%�i�u�ϭ����_"�.�d��9�-��0�B,���[�97.~i���%���M\H YQM��\��!�,7�YS�A�Zx�J����`Pu�f�?H�*i���϶׭WR��GSsH%�s3��iI/%�S��%�n�C)����h�I��4�/�!�S�hv�։��%�5�{�\���9wm-�UYo���6�x���b�2cu/Q�pK�cx���'�	X���N�,��ғw��S���+v��5+�+άՖ��hA�Y>��ld0r<�^�_���Ѷ*�ִ�٣e���+wkc�sq�j���e܆p1���Q`)ͭU�V��~�3J	��ĺ�f��e�VT��[��Z�M��Z�J�m]âũ����ť� ��L+�˨���	��t��	Z!h}��)�a�9�|
�)��)���h�k7���ӏv��W7F�M�2��T���W� ��9nE�Rh9Q�!���]o�b�ignC	32"9 ���5����V���@L�^cɻ��\�/�jJQ��Z�=xym��Ҋ�_0�pc��?������?��1�A@�h�U���Q*�<yqs�
 Z�j����Dk�ϻ��T��"�xAˌ�;�!l�48����v]�F��ʒ�z����n[��������qP;	�l@9yj�wm)=OsJ��c�Ʀc�ɥu�5k�Ҭ%��M�keW�xe��ƏUx��b�n�ܐ�w+Y��;�:�kW���L�zG��L ����n�,�Xv�\�K�L|u���%;�5�ו���y�~����!`=�=+��3OP~/a����δ�g�7���&�_���Z{YYeBM�k�F�����j�\��0f����δU]o(�7C=�;����@ӊ�>(Z48��\������s�"��7�k;W�J���b���)�WH�/�9�-�~���t��}ᐰ��*��Yo
F�8PH����`�㞠qlL��Ԝ.=j�)��4�`JBi����TNj8���9��ʙ�4o&��Z5	~��o�	ܳ*�g��pǺ%rFFF��A �
���������.?Z=~iô���p��g|�ޮ�_!�l�;�/"��X	a�]��B���K��� �NB�`е�s��$|?��g������m�Q�P���غ�\$f�#�B��pM^ω�@�3���?GdB�h0oycv�+Q�@֤���7���D��W0ҿF�����b��V��`/͆��3�o{m7�� �R�|?��]$?xYw�f�~ΌՎ՜��B�>��Ղvk*�U��������|�ejg�2�=]��JM���0���zיͿ���]�ߡ<��������轪L쌇� Pխ&0u�､7�
�	k7Gm��V$R&�'�\�kK��\Ԥ�n��:J�Ӝ�}"+h��7D���v�2��uQ��j�"J��n\��6lF�(S�I�4h-��@�b�<?d4H��C�/��@0��g�H�і=���۲z���tk۷&p��RJ ������c�IXׇ�)�����ru]j%!=�i꣯ް�|͞|�1c�����)�"�>�����ؿ{_�8<g�_V��62a�]���p��^*�U��\Z"��u�&�5]�F�n�F�u+̝�?&즽uC}�����������/3{���*-���L:�z�Nc�񘲟��C�Af��X ZBZ��~���u�5�[χ�i��#���+���Y�������ҫg�x�^U-��:k��ƥ>��=n��?�]Wm���Mb�����J�VU�j/ 7� 0��X�bL���k���-΀�_k��3{����]��1�;�b�RM��\KX�YBU�]�{�Tն5Vָ6� Ɨ�  ��s���K+v���=�@�9��{��#P���o�w�j��%X������c�*�����ϟ�y��(�iYpj2\��4�5ګ�g]3OX�O���7(^���61;O��ȵ
�Za��p�TnA��=�S�����q�e�V�ڛŪ`b�/@
�:���)��"��Si����V�T�_h�w�>�����#��O���ZҘt��&g�HY
�@a�dU�{�a5�|�5c���j���w~5�
�=6=�������z�fH�-���C2��x�y;k��6B��'6}o'�)NҧJ�h�i��(_	.x�o���Qi�)B��� T0�V�J�u��e���Yߧ���*?4��d� ���Ґ ~�+���r{V�򼒮z�B*����hĬ
 ��·����~��_��o�u�P>��Ma��5rd�Delx������TԪ5�����N�@�N�L�3t��� �oC�����lW���H��}H��\��=Ϋ9`�x�V�A4*�eǧ��ݱ�W�� �_[�Дĳ��"e�� z.�&`�>����w��z�$��m��21a'��!_��L!��ڸޕf���X�[�e� 2���E�X��%.�Bq䆴i:��'mы��4��؍�os��:5
z#�rgε7�k$V�i��n�����s�ZCh��l:�1K�5<;*�U�+���n0Y��z��P���T�z}>���%�� ֛�lmI.��"�	jAb��܄ �%m-sc7r4Q�轍��`k�F�F��\�Z�wTe�>���C�ʰv��qvR�exp�����;����`�� Ve�k��"�٭�BG����t.����1ַګ�}k�#��
�g�w��p���r��OI�@��#a�!:��\�T->z��l�k�v�������ܲ�օr�BP��D���ƺ�E�s6�v�ӄ�SC�i���}��k���k7�{(%X�M�  ��',�ջ���zbI���w
Ӯ4񯭤��X���Ȍ�܃���e�vAm�%��������҄���U�9'^��?a��.�u�t�A������Da��p����W�0��~�~~ $�LM�C=]��*gY���������u}��-��,z>tu�6}�g�I������L�&W��(�&Ѹ4��\M5�i������[#w?��ǯZ�
Zf�c�F�]5R�R�mk���ڃ���l����ͳ����/��%9��'�`�83�IZQ���z�$��/ ����Pl���vc���5^LF�"�Q�X[5W�W�0�ت]z��ucn���Wʉ��{1 ӵ²�L���c�u���9�������A�Z��W[��f�tn�+�.Ř3��}�zs�.1�5�'A����cS�h�
;�fˍ�����*�8 5��SA�FkN=�Z�[�s��=����Z��pu���P��Y^A��s�t��C{���?w���:[�C�/��H��y[�J&W�p
\�\iۄ�3F�oܞ����e��W�lU8�5���_F��ю��ͰΧhW���yꥸF�D�չh���-(m!�n��U�2{U�W³&���.9x	ht���\cx<��)�=O�3wD%L[$�����8Xj��/����8>)
Q*�8���6�P�� ���,��oͷ�������?��_{ ��3m]kH����fdd,�� ��my���?��/��߼�n��(��>��0���VN����\�3R'�An�sVG��	@�v4@B&���?� �hƚ^���>�.C^�ہH�񦜹Uq�AO]�c�:��� ]�N��{�e�?^kװ�$�*�$��W
�
�ٺ�?MѼۆ�=0儸i>ż6�~�۲t����;��-���w�1��J:�|�ML�?��s����-{�6�%A�[Q�Y������(�M�� �}� ��|�7�����¸���pe�6gu�l�t���2�iv��^3ۭu���T[Dh����Ao|i�z�Zu�έ�����B��������);=�w��X J"���zk�f�B]��Đ���JzCt{Sz��O7����+�{`}����n��-�}Шy�^�����b;����/	$D���	���a$�"Y�Wx�/�	ށ<�Ey�B!� H��DV�p$�˟����9����=/���Q����ٷ��{��{�}����Y�fͪQUc��o���<�g9�&��d���B�Np�Zw�fq�`F	�@��$ E`�ò�"wY�� �3���.l6��O�������.����N��_��0<�~pG '��@*�Do+5,Cr��C��ے�}�UV��m,��.��ez�v����@���eBQk�)�-�)��D"s1뇑�a��Ɯ�u�G.MmD]�ɺ#q`钕��e�Y�ΦY#L��^��0V��	0����=����-���6'����b� 7N�����~�c�s�cJ��+��/����/���Շ�'�8\1�%�F�(l�[PۙB�����+�֒��R���T��9��m�m*RSN!����n�Q��h$� 	G݂)Q��/���7���Xװ�4=�u���[��L�=��:�P��z} _�Y��s;�6.K飇�F0n�+c�f������
��X-eA[Y���KvW�d��6�NT:0��0����gp�bn5kn8��vs�A�{����3� �� {��L�� ������h���G��,�8��w �3 ��S��?F��$� �X��Ҵ��eκ �]���7c���i�zeq2�;�� �Sh�����)�\�l h۱�sd}���!�w౨���mH˶�K��>� ���C�&��;�X�ԍ�:���g�Y}�-�@{��7��N�y����3K9ꋰ��%ٻc�J�O��}��M��h�4}�/�F�P�l*m� ����z�pO��C����O��B;�o�����!��G��ġ*m�m�;�f���d��_�����w��������Ҙ����2� �,�] x�S���|��/����f{r�zM��I�_�����Z�ј�H��N�(��(�:(h>ܭ8�KA��C5�h�eu�/%��:�)�8�hM|�su��1��Q���,�k���%GP4�G��K���/��C:!�Q���]fhĀ�v�V{$��خ�z���ථ�K��vD�i*�8ΏW4���f��lt��U���u'1�&,��o����]Ǐ�aj���;�!�aTw�k���i�����9d�D��8�_~kL��kD�ج�8GIsxU��V�Aw`%�4�[��\�C��q@D�Á#-�sn�L�q����t�/�|�ց$�3�#(}� e��b���F>���&�q(I4,  �/s�-�»�lH������l`��t�>`�C�(JrВ(R�G�U��n>\h,]���L�<µ ݂�V.��go�^Bߦ�Sg��;�e��k�ں\� ���8��QE)aF�EJA�1�o�u��0��s�)5v�Ư�j��[3���GЍN٠��0JC����>��Ӓ��������Gt�f�  ͩlkIi��\ʆm��:�st�T�&�BC�
g��Q�\߸s��%�ɼ�l
� � @�{a9�z��m�5�ɞ
m�Q�,�Jm�vӫڲ�w��|��e�F�v^%�)��~� �U5�7wH��80�8t' }V�k� [��8��<f��S�	�����^�~홒���nE  io�R,�<;�\�t%`���#z���%^~1��W9;��hep�9��J��l	����Kj��Kn7D��\"��ޡ���mS�[*9��`@���i:A���Ř���M�{y!�^"z��C�X��b�_}&�S�������c���x����n�*7����q�� ��U�E�_�W/��>{���Iʬs���R��?�\�F��װ>@����x!@$Mۆ��ݵ0"�U�%J�����7�9�BӮؿ��X���1��j6>0	��de���T�W¬Pk����Gph�؀Y��:�2�����L�OF���3��Ӭ:r���!��tܸ� ��`��z;k�Q-�+�Q��D�y�Jm�H�����5���2�y\5��V��MJ�T�c�]���Җ�os`[�����z8v�w��J�8�ۿEu����(�1>���m�ʈْ�r�ةR���)z���Bٱ�g΂�y \,أ�,�IF't�������?���N����
�Q��2� ����.��n�̨<6�͘��Dт��2<�Έ<���e�H�oP��M{٠Q��ņk�91�:@��wR�8���)�[���=MRZ�n}��-~9���գݵ��b5�o�aU������z����%,�o/�^�;꼋�y��� ��C�a�q�HD����N�Z��	::ɘƷ*Fΐ�(���>�I�.b���0Ph6��}Ƒ�0
�]�(=���(c������V;Zu� <�9�(}��*��٤�ǎ�=b���eN'M;g._g�E��M��@�y_r�;��?2Mp�r4=%���{�'.�� *R��l�C�([?��-h���ώ�L��-��Zm+e΋n%�4G��<�P1D�`؂c�*�=z}�d�qP�^�����aԅ���d�� �N˔Lj��$v�N����2����D����(q�r?v9��)f���
��X��9ϨD(c�w0z��9�t��)2J��܉#4߈H�MKGY�jd��q�W�T���{D���#z��q�3��ʆ�TX%�ԯ�+]��U����
��Hsֿc�.�(�HYa[}j�5����NI�Ug�?���O�6�=5�Ǩ��C�=>7�G�(?�08j7f�>�ZN�{��)���o�O�9���=�y�T���� {� poݷMT$�@H�81��t#y�+~��-��M�'��'0�%^����G�|u���9;�%�:�����'wm��8� <��c���q<�u"r���a�x�+�%��ޕ��Fc���  �L���=�e8k�0�}�+`-0a`Ō���Q��Np�g�sj<��9^�%i�*:�� �/e�����1}��W8�/�I�q�N}ľke��YW+z�~Q����e�`ɶ +�v	�����.,)ό�@_U��Xea����8��{ܬ�]Ь��_��5�� V����1��`�=_߭[xMe�5땺��� T�L�/�+�m��E#�uR�K���Z��=�����$�.���|Jo�x�)w�
i�3���w�OBY�r(��}�h�S�U�9��W���e��h��l��	��ʄ�9c��n�H�$��$�N�~��І���߇^�}�mk@�M��u�}0�+����+ߋ�~%0�U|��Z��$���S��~��^��?��Ze�AY*�  ���=:ed�� u���W$�jcD�S��j�ӇIeމ�dZ ����~y��9}^�H$e@����!ey�@�Rw��ӊ*�_��^�o���#8�#�@O�ۓy��I���s�4���@ �:�[n߱��Kh/��M��}M��\g�1����u7���Z�[�;��-���� �(�p9P+R����1��w�ߺ��.2�J6�1}h�q?&�9*��
g	:3��nE�?��\��Q?>�8:���G�K�����:Y\��'3�XG�<1�pT������ѯ��
��u}�F[U�>�7� .S�"���3�ҕ~�ؠ�[Q��Z>�a"�RB1G�:w���&�(��lt~���Q��ca|@����H�');����*6��1��}Q0
�l]�~j��K�^l8��9��#��%��[�@
�y{� b��KR���<�Ҷ0N3x�b�b�	�')҅T{ҳ눑yT���4��rD�0�}��^6�A��N�46zУ�����(E: 8��E;ø�N�$a��i�{� �Y3��^�{J��LL�>E��
�8�&�H����HN2M�$k:�UY";p^������Ab'�sH���jU;�U�N+�kq>��f�ꔏ� 
�PE��B�c����~K���̼������y��.+�p� m���� C���8Ve�sQ�&��Bd:;Sߌ�q�ѹ�O\��y����ش�X�����J�A������R"��N$�
t����ֳ)L<e��D��	��-,5H4�X���K�
��A�\ȶ*�Ҿu���K��� ���8m�܊)�G.�BҴ�甇���+���p�_:�����r����W��Q'�r�9��`Zv}�U+�|Ip׬  �	ɸH�"iHF�.�vH;�w�����
�����7������#:��8Ě����{Sȣ�m�84���(k���f<?	�݊��<�^Z�gw�
�$����6���U��/�Қ�	�����y�&�)sT�3�߿�7=�e�ݣ����ڋT�S.�u7���������o��S.u����-ɬ>��jk\�6���G��7��ڙ�uM�zDR>GeD����!z�r��|T��G��
P��qz�Y%��)I�m2��Y���������x��MC�� ��Xv `-�/�ǋ��Ο�~���դ��L��,L%Q���#;e����2	����c���6Q乻��si���t��g���ue���Q�}b���0I��V7�����B�� rΏ�tS�5;��T-㥀���b��ۓ�|�k/F�u�Mn��j�嵏o3���	�}���S̃�ϋα�Zc�#�\�=�^v�u��I{FG��C��D������X�S��>�o��g�k��I���`U͆��}�4�c�	h�2�0�\H�* �ڥ�kݞ����Q�	^�~�����Yr�a�U}���O)>ǧ)�=?�H�����&��08�,l�M��Y~\P�.T �/8�����&���v��e]�36�W�R�n��u���d.�-���׹8|F0θ�Լ`p"�8ڤ��c?q즮qu,T�J�Sŋi�(����Dˡj����}��
�yJ���K�I`6�s��#&����F��J�*���J�F�4��1���x���]�08�0~e���Z1�<�p>�}��C��1��T�_��ۥnP��kƭ!0/�Nk��٨����/��t��H7�[�Qh��"��0�=�'��I�{� ��ep\ͨ
uܵt�	n� ���Y���"u�QX��|L9RN5
��S+X���<^�hLꞂ��uF���Y����� �6��Jo��mH�m�ԥ��yr/T��;[�+nݥ+o>�!rQ���٬/ 2<:'��Q��on��mM��������VD �kE�/\�iS��X7\���7��_O�wř��&�������'��w&��.ak����zG�6+���%�,���H*�(<W0�A�%nc��׆A��ź|��i�=ᜄ��XBd=�_��A� �@� g��>Q���τ���K�l���F�U *pZ�Ή��0�a@���2��5}� � q��m쿿�`)Xc��o �;�0U�y.=��V�:�}-�������0<4�~��@�f9���A��$��]󼡃+z�)�S����
��)�M�&���0*H*.�9�6���S!��_x~8��k UV(!�8����"���iR0h�`l@��q�ް�}�qL�L/�� �v�`���	}�G�l[�b�B�����3Q'a»����G��H��u�����(a�&�5�c��������$Ng,/[GQ�V׬⫑�M�ՙ�ղ��؎;5ܚ����~�W8մ���zW/��8���X������V�~�8�޷�6������6 �����i���گ������d��3z$�� ����> �����?�������{���W��wIe����?;�� �t���ȁ�d��W�$�y�]a>�_XZI[��F�{ӊ`n�-R���ä�N��}N�U`ş�¼r��=�Q�4Z%�I�K���E�8XL� wD���Vz�5��2�Q���8�摃����s�ю��u,bÃM������`&H節t.iv'ɒ�W"��s=��a�P��6�Fh��Ȥt��)~5 9�0:�t�z��� |���Pe'��s
Jdl�����S�%���a�F<��OXs{+Hx✳%�?L�go>N�a����I�4\f0xL{'��E�c*�r`��~{��d�O���b�a���lϻ�e��J����<��FFM9�7�X��.�h����nm�:ԣ�
:o���4��Nq�q��p���W
6�c,�/p�^!U��mt0r�u{�<����į%��EK~�f&�2�r��M�h��!�Ց�l%����5E�L�[��;�-
�d�7͠�<e��K�qTA1s &�_L��ށ��j��e�ᄆ��Q?"Q}��>��}�Y7�mpՙ��� W��tF��5�ry~G)W-ǧei��Ij��>���Q�X#��G��8onS!�Ǯ�6����� 24sIj�I�f:���S�}�S�}�Lb�� +还kPA�j�T���n��믳�/$.�^���T���Z&6:�F���3�����w��z|�Vd����R������βB��qN��]Ю 8ù���:6�e�0�m��;������nO�w�݂�ρ3��Z��K �G��ĎK2.��"췶�t�=��Ւ��wge%N@������tz.�%�>>u��D"�~ړ"� �p�cX��㳜��l��/���s������gU��%>M��Ƀ�7L�>EP�@�d�3u@ �H���Ϳ�<��/��Ti���:�{�q�� ��������ūU�p�m��/�+��J�Z�\ku��Y��N���V�u���u Y�|�v�,�d5a��pe�՘���x?(m�U��]��wF��+gg`us������-k�f���U��W���x�m�Ԥr�A�0���e֭�ȧ��~����J-���.���3f�������f��.8XF柔'��viX){S�;�^�=~Zv�e�]�m��>�C�9:M�r�Ƿ��!D>7�����)*�����3}�����?����OT?N��
:���fA�H���w�"�:+P�{g�w�䕝�g����������e�K?�7?�S?w����������Ad�%�S  (H y�O�8������/��sS�7u���6>#e@E��e����`��:ޕ���m�c[J�+d���������S��<߮�Z��C�_8j���D' �̀8�T�`�NT����&��6n��Z�6`����֞�u�%�^ d��]Ȯ��,א��t���h�l�a\~�lp������>�-ر
��3�����۝ؐ#������J�[
)U�h$��<Oِ.����snD5�S�^g��U1`
�;30���4}!9n6�#��6�!�u+W�o�V���'�F5�B퓎��8������^�0���$��ٸ�G�����y���occ���
u6�pA��
��rD�s$W���r����
Z]�����l���3�����p! ���$ ��6��0�Z�����4�`�  ����&\w6 �Շ�����8%���6~��I�y.�����ĉ}pWӵ)��ڈs�ġ���5i9_��<΃�Às}���`�҇����`t1p� �S#�K����&f㡝��'[ �����޸���0���+*U�ṫ>�˃�^Ġ[�_x.�`01<�s����]���]�F��x7�5�� �3��r:c	�6����,���EE��Z(}��˜���v_bG�qFK+N0D��	�4\`5��kַp c������Zr-O���-��#���<ɉ[�c��5tW�^=��$�ҳ�r�qN6�b�R�B���������nc�w�K4-��'�_���&M��|�Ӊ)5�>�.�a"U�X
.��Q
1���B��˭|�� ���D�i6�7�kX���h���8e����N!&Ӊ8���_�y�:pv�s�1?��y�xD�c�Θ^_�
�F9�2g���|�40��hu����ȋǆ`A��Θ3x��L��y�:am��ُ��
  ���=��@�ME�z�'(Z�;N��.�UT9N���У����R��_ʾ����03�ZeC�~?���T���r��?Ю/3::K�0 ���B�Y��:����~s�aE��1H��K4��]��R�a�)�]Hq i�)�G����2�uo��Lx�}fYj懯$���W0��T.��{�P���d�t;I�Yo���D�w��_��gqdb7��H> �f�W��0.`TKwW��P��#?ET)�.�����w���߭g��t���Ɏ��.��ML���)x�C�g�y��d�h��_�g��$In/�m  �2�
���Ͱ\K��'�����/�������ʻd�C]�JUR�(}��(��2��f!V��ڻ�K��<M�Fk�}�}\�b�u���k_G=�F�_7fVSK��2`#X��- �$Y����A���>��O �DמT�s�t vsF�e�����eR�[H�M��٦s�2�-kw�x���j�s�b�N����#�5��L��Bu�(��pD|3�D?�qL��\Sjx�<�X��7�����T� `����ɏ0�t�q��h�9�UY9 �R"�ضoč!�v���q;`�<��I�c�%^�������Q���X��s���䢭�� �)�vhW� �}'օ�)��(u6;� ��cEW��)�0a��s���\�Έs$F��E|�`u�h�u��'��	��i��5"�`xB{����_= ��9Ͼ������(J<���y�7�^ m. C ̜C����ڪ�y�l���\�9��/���a�w6�  5; q�)���pF�.jG
��ڶ�[�u��[�G�k��l�8�`������mIￖ��/���.�E�����!��`@ۗ�ޗ�	�[�����Y������Ǝ�u�ȼ�ъv�'��s�n*����\���v��o�����x�PջMU�S�'��4�	���%5@nw�޽z/k2����q >�ۣ��ԋ�}�:��k�u����!k����-�J�|o�K�Rgp�7S�"�|�g�ϾY�Y��݋�����̱��=�eR�������KY�΀�Cps\6��9>P�����H[٬��Fv��z�{ k�����) X9���3��~�f��U�\8�B"W�^�Ի.��#��>sm 6y/A�}{��+��Y�3�E�o�����J֬.e�-�d`;n�>n��I�yz���v?���lx�L�s�&��R����}�\��p�x! �Z"g=�D�����f2�^�0�q;�u�a�g� ��G|'f�����ʥ�����}k�s7�� �s�I����b'�믋���1q����bўLU_�&W
%}.�'�e�$ ҭ���N�Vn]�����%Rh���7ca��L�VX��Dͱ�>x�t��������2��d���MsI�Ѵ�����(��=�.u�ɩ�s �${y�	g����^_�y���8  X�3�`3_�;��v�̖U��w�햏,g���-��`�k��������p���t�5;�)���g�6���K������a\���'���`�H��ǇX+���/I��M'RYvj�B*��������̣R���ˬ������ꧾ1���β{����T�2���>  ,y��&�����WTg��2Vt���y �.U޾��(D�r�ET���CgL���U�[��<2Fr��� :�%�hjM# (0w(Oi49Ŕ2θ��V'��W�(�S�5�[���8=����T#Nq�2�h]C1kr�V{r�k+A��E�|V�PFL)��>�h�G��w��Y�����"�Y���kG�f��f����늍`o8 ��SG5*��'_���'?�ƪύ�t3*�zN�gkq^⌝��|�RZ]FE��m�f��Q]Hl(I�S6�:�C���p��ǉ��3w����Lꄺ�X�R9��͜za�l�]'�F|F7�36����F>vrɉզ��E����i�y�k���#9h�V��g�,i�	QR�gr���<$iw��C���JT	�&���q��!G��fp�̖ s+�_a����.��m�(D�9_y�ޜ{8_a�4����_�#�.�3��<X%�����X�`�T &it�8�ۏ�^T��*y����&��w��DԳ4�'�/�N�QH������q-�y,��0��~F{B?#��k���|-�Y�5�@����\%�,��Go�K�"��F\��00C�sn�f�p�
���;!��vu�-u�(�`lѧ�.��v��E��9��ٵ�� ��l�G �ss���v�����QM���Ȇu�z���u`-���������N8Zs���95r�U��t�BY��]�i����c?���l�8u�2v`&.�SE�=�m��{�u�ѵ�ˁ�k�f]}��0�n��#�X�͐7������� h��-$��֚��v%^�{�s��\�H�w�"���Ǻl����� )� X�J �8q�5}֑\�]Fw��!MC`d^E��̂w�A��h�r��`7�����q �f�A��wu���C��N6��a<��yA?@�.��\�ku�N���fM`�p��L��I-���p���$ז�r2���H��J=X��Q�Zݓv�Q�K�
��F��X?ja4x�~v{,Ɯ�<�%�PQ�&r/`��i���M��9�>�tG/��Ǝ(c��ɺ�E�5����5��uz�*�?ӊ��aW��n�@�'�ە�݄�yw�b��a�9�ǩ�Y�7_g��g2��7Θ�-���m���}1u ����c`6 0!����]ʒf]fļ�J2KJJ�#�5�K}K��s�^5:�����3v��MB�pc��� *H��bw�&cBX~T'��ѠP,(���nY�H%�'��$i�^�����Q>1�Ls;m&�Ѱ�d�AV�^  Y#������o]~S}8�ש��c�!��C(��Q�% �"QGx�U;����K^���Q{t� 
����x�͂��d����'_��\��ld��H�zB�jBii�jZhz���Y-�U&bԉ�(:q苢�2���̝���1m��|�js)Ď�y �N{�<�( �=*��+��}������Ls8u�!���Q?b����3 �򕉀Wj�އE��>8�˗Y�>c���Y"�m�XWQ��nz� �s���t,zp��ٛ�܎��ߗD�9X���S�T���h�?sєW	]_�t�qDg�%.�3�F1��`�wOI�B$o�>`��t�E?�:�#�%J�DM�_fl(C�E��Nwm��:w;U�Nee�� � ��i�����c0K�O�O����ǈ�ݨ|L�Jy��B��?" �9z�5���?޿|�SЦ���c���q_��nr�KPW[�N��+��,�9H���A�8���0�N� ?��c�i���c�\�9�Ҩ�H��԰�q�^E�Ɛ�cI�p|��Z��X�-"8�oZѝs�2��<�:�Θ�8��is�S�ʊ�)u��
5������w�[(s��C��`61<?�q
��9�x�`92��rz�E����g!��]��U��洷�EJVy��~�s/@�s<g1�"R��e�N��S��'�ޭ�~������$͑�ł�Д1j;�CQ�n�e^�,��fR���s��SM� :�T��u�\��ѻy�C�?��`+����n�:m�O��`�q��m� VV��>^(;��y�s��󙘲��9-o�	��5��_S����l/$�����jN��Qrc-�+8����쨙C�� ������:6��X�ɭ/�r󳕹ij+�����%8eי0,�O`���Q��R��_S��c��,���M��}n�'�/ �t�tE;� ���dL�'?w֯N_�{���V�������?vlmif�9^�|��hZIz��p���^Nw��/��XK
+^���3�m�uø��8�U��m0ߙh~�`�,�  ��`���{�K�r@�p/�%�g��������|Y0������Zu>��+هUT;�eE_dn�[@RP��ڪYÔis$�mQ/+h�)�[~��������8�|�W����&ql�,�{tE��j��4��R_G�Y�9H��k4-B�4���a�t*MS33c3�ܴ� ���� `�>)�������;������?2gS*ַ��s������.��J������<�t�yZz�n�^qw���x���i	�i9%f����Cz�x�8%�Al�9JO�3ù���Pο#�/5zx�x�e�ʥ�����m�h;��m�Q�c�a2n�'P��D�c�� +E��[ې�w�6S�5?$j���I�6(*���b��dR
�/6����T��`��Ⱦ���zr��k�z+�;J%W&�M�Kh�cK�ΐ�9��p�>�K�d�s	�N�P�N�CR���LOk�78��<H���*K�sjӛ��wѳ�E�1�4n��>���|,%?kL߸<�0��n���1Gu�I�e�۔����_Gimx�j�1
�B��-"eJ�ں��hb�W�E""
��AK��w����\���6n`Q�sL��%�Ɗ&~���Ff�_y�HO����\b[�Q �(�?p6 �7�_���bZY	�d��)7����a ųS�kg@���ɺ �jd?�ᯕ�&>��&���kg+`u��b�.��X'P�1���X�� `w99kt�F��Y�:�՝D�3��u�{����U�������}�D����6�,m��Ǹ��(ԙ���ok��$�r�-M5y'��W�!8�FNv�-�d�Dዾ���[�zg8���G�I����K��_��
K [M�]�(�Ŵ�SM��r��E�P�#�fA��<5��C��+8�X�� �h}�^�tO��B�Ly(�7��6�����I�j�SUځ�b���ֺN�b^@T]�Q���}�č�����~���t.�I�����������Ѳ�WH��f/v4c&���,w��T@����>u@w���6i�꿩�����S��fU�*��3���(�v�F�Yv/k/����x��9 P���j=l!��F�W���t
p�c��Ž0��.�~p,�H����N����qǏ#f>j]|^4C���Xy�>R��o�����Y�̒��n,�Ḷ���`��f��J�+k6��T��d��kGD����^����"x�dB0il��S=+��;��i��� o�$�oչO6˳ ڌ��FJ|�c+<�Ք�X�fh��25�z3���������?�O��˳��)�FMфd�A�Ȯ ������������o��'���0Hy�h6�6��I����� Z�<Rʸ�;E�l�� ���:��zђ���xu�uuJ�H'�8���t
p��t�5���%��uA�Ԃ%}u��Rk�y�gB�di�k�S�.A�?�f�;��f�᡹l�w��=ᶥc�j��t�[,믷�	� �r�u�Yd�[�1K>-������Zr��&@9��[����,,��e�y376��	C�8T*n��E.��❨ܦ�׆��1mf���2��R*�Ӯ7�����=e���i����o>�����˪bp�
G���#�q�����B8��Dx!@����J�Ն<Ѥy��� }�G��}'9�b��?��f>ʏR�s��bL���\ը7S�Q�vA���,Sn?b�1�N�f>A4\9�����V����F�DHE������[�����
=�lC�8�E�w���m[7��`��C=G����FZ�5��:+�G��pYrmg`�	QT�U�c:Sp��9}{m�U��m�ǡd8��� K�P��#}�d��j���"��z�{��ͧ���E Z��� X#�S�pn�cx$�Q�vy4��	2KDa�T͕�qf�n0|��ɤ�H���ŉ�;�r|`���g��wC�o��<�������M�:n�ȩ\�<C�,����?r:�V�@"�*em&Q��Zl���:��[սxϭ/k�utɢS[c%�H�������±��xP{SU����Y �@G0�Q&�L6^ۄ�������_��~��O�^��d�W�ky�Xy�8�}��E ]��"�m�K	����FU�i��n"c��_?�|�+�S��Q�u� й�'
 ౩)�6n z�X�@O ����U�m�@b^#�F�ߋ �����YR��"�`�����-��-	ϳ��U���k��p�u [v��6��y��}�C����P���w$� ���c��K�͜�i& Y����c�i���j�2ev�L<�л�H�j��{0��cJ5���-��"6=���Ǖc>_���V$.x7�J�.�E��`��ɲނ~H���W���{��l\���U%%���7c���.�(i�i9j�v�XHl�x/5S?�|���_FF��p��/n�<b���~M�J��f����i�V�����9�|X瘴�i�֧��̒�����~�;�������_��˗/����s�V+d�AY ;O���������L�/��eY�c�P�Ġ��w���3��L{]�i��r�F�1#����KM
��6����5s{�GZ�	'�ȴY l4!_��B%";�f!:�̩lf�̦����ͬګ�>Ь�(i�g6�Ѻ��d#�L��a�(
?��ͳ���-�c�eC��_�`�	�8���9�M��!݅���eC�3���;���j�ޫ8�R6��r�z��A�"z�sz�䢕��+��P�[��Ȼ�//�S<��6��=>�����H��6�l
،���N�sτ"�}����Ԝ�Nj�!tFJ8���~�{eCyڊ��8"^@����?s V�_"�Rȋ���3w/ތ�6uN��w��a�f4��q4�Ķ�����3q�c�U� �a�Q6 uD��d�w��f�Wc���Ug�{���P�����ԩc`1��3Ո/k�(j4�u�%�XgN���ظ}��sA�w[��v!�*�IY�r"Fif
j�3��V��la��Q|��kRY/3���Nu���m�z��!�3��%��a>�e��AFB��iUܳ/��uT��*}�tM�s���mK#���,^��.[G�,�)#��qX/_�ȁd����L`�31�J��a�k�]!q:�S���G�[oQ�a9���z`z���!�$v�u'��U�2 �Z�YԦ��f����D�G�X����w<w�n�A7���.lWD�{#ԛ�Y�[#p~��S���n_=�]}�,�P�7���o��:����U�C名�N�V�hͺ����.�m�\�:\1�e�3(ß�&h��Y7d�UЉD"sŶ�zN�j*kl� ��C��nۓ8���3�S��u�ܡ�s��g#�& ��w������o���
�A�U���Tl�6)i�7c�߾���R�6�3�x�W�)��9��t#w%�WHLB�X��!��VR8;P�w����li��c`Μ�ߕ�N7@Q��b����(SW�>�Ҍ�*�3{q5�y����:}����pK�2� Kd� H�����tj�ܚ:��J
=�ZIv
:5� �s�$�=��'U�mǵH�t�՝ 1����hU�y��|�޻M��ݽ��&��`�\:�>beoDqs'I��Ԩp�h&����ǆF�gt��n��Wd�'��?��oYu�P��i;��[1��Yn�ڸ����6:6DP	ӾNH������>����4b;ox����*2"�Ԑ�cǒ�qMb�Xu�F���d���W̼M�#����v^"��9����;}�:g�=�R3�;RB`3^"F'��O?���tv9�(�<�ʭS&;��i
Տg
JN��E^d����-��B����J5L�
���eN/s~?>�(O�	��I%j�4ګ�Ce�~���;���E���i��<@���o�d�lO,��#�845�y٪#��<&I��Qjp�"�9��7������Vd[:�̋���CA��ĭ����ǏY'��LM��"�՘/�u�z:*$zӷ�^�>�SK�c��S[%[�mPG$����ߖ#�â� _��v��|�?����v���R:�L�v�/-����X��߇�ђ��1��9��r�������ӵ�4�A*���V��μ��O����ҡi.zY�F��}�r�k��*�N���|�?i�� �L�b:�_m�AQ�k
:;w���W�'�>"7� m�/=�v����o�����TׯN�ZG��:���a����6�	HJ��:�����'�O�l��&4!�k��v	i�J45����e�+��,x�K���D��j�b7PM)"���������1}H�T��GT| �7�lBi�~�� �S�#u%N��M��ު���T�]�F�����)�-��~r�om�un�����Lُ�@U[6seI��E���o�w��Ƴ$��L>� ��Pv �?����U��(�{7����,j(��+`uLw�҂�_G��(����;�������t!��o\���S�azV�]�?�1��Y&R�ZUg�i^E�d�C�Q��Q����������I0R��\ϭ1�l�^�ns�q����Ĳ�ye��>{;ߦ��E,�S -��N��V\?�'��N���a1�:�Yt���S�Bؘ���ƃt�F�c+���=VmԻ�w{����Am���f�}|��ū�Ӛ��J��G: DAV"sT��@�	]�i2b ��ˀ���y�]
N��{4���"�
�PF%�9�W%]�-���͵%/E�0���2o^#~@�h���.�x-�M��/A׉@�O[v�6%�3cpTi������qς���c���L��['�۟�hn��E����H��1���.���Zk7��/�ֽ�Jj��v�9�A�ا8����.�h���Y%�\���Y@�L�y� ��E�!mfb�"�ݧ+�ֱV�v�wT�a�Ǝ��a-��F�[�����C�����kN0�y�+'	h�Ykr�W���y�u����m��%;��������ۛ)�	�r`��f�-��:�8�~�t��1Mj(Е��g�h��k��қ6J�B��H�Ω��������O�DJ�&v��虘��=�Ӿ�.}�, 3/I����Y��"i�=́͡+��'[��^;��c��T���q�����f�%�];���c�ჿeW��h�=�zm(��||�b�{���l�1]��o���� ���7���i��WrJ˓}I�?�yEU:a�3l_k�s~%�L�`��� ��M�ܵZ����_�]� ���ѕQ�}��O��_Zw�T$�?_eRTg����R�� ��Y����������G�M43� �|��s @����������o�����ۛ�d:>>nTai*w t� �]���\�G�;u�����^'=E�%�߀�l9�Jڸ�Ztˏìl\VX�[-��Z��4��J\��7Ln���"�Q�2����T����Usn��6`"D�w&���&䙱��4�� �S#���}��'lӦ���$��}6�"6�ɕ\kD��acw�S�\E5�T�	�l�������L�/�� ���.炷�e	ݼ+�1rV4�$�x�2��� ��U�m�En�,yq'���/骹���YS��i��0S��'��?)���?>�h4J�PV�(�z�`����A�6F;H��Eg�Ƥ����χ�G���!H�:I�ǧ�Ld7��F�k�/GQ�@G�]>`>[e��<�g�ʲ ���67�ot���i�V��+�͑B�K�@�Fk��̞��������d}WV���.��Zwk;ET�f��P�kP4(��ș�C��b>���C��F�M���f�ᮙ��A�giD���M�.nS#�3���������ct�6�h�ɽ�YO*���+�R��-��s������{�F؟���J��U�Ƨ������������5�ԲcQ�i�\N�����HR����)`���A O��^=Bt�^�.�a��ϟ;z���=M��>�`-OJ��}�ֈ�FS0۳�0QoJs�
��}�Q)�Ebi�4��L��{��bz�"1������-��gh�u:����Z�����Jⶰ
 ��$��3�/��,�C5<%�Aj~��v��ʿ�uvrt4��jF�� ��Bv ��/^�ɻ_�ſ�������ۿ��_�ߵ#�V�6@qi��W�^������<�TW[�>�Z^�����??,R�!�:�}���g%A���g~��ˏ|7UsߘԔ�����f�eE�ֺf�߽��y9��nJ�T'�N;D�.P�:å1�h�C���[NL���J�F��J���,c-�/x���U<T{��.��Q�g��]/dr���6���j�9�a',)'*��ҕX�� 7��sD�W��M!��+eQ��I!*�*�����1?�㳴��'4kN>��K
�Xz���U�a'�䶢�%}x;��_O C�s��	q^��qJ�/2z�fL�_���e��a�mQFi����������~������y�X�ܘ_%~^�3 <B6����*+��D��Q
�$���[��6�0٦�_���|:]`)�������޺X���ֹ� C��AO�� ���zw�#n��6oݩlr�e47�?Y�C֯gv�v�+~��3��|�TԼ�֡;O3eU�+�z��q���>�d\��
�9�W�U��6�v�F/�UP�׆�mQ�ۦ�%����6�q� ��MEE)�!��gӊ�2:�J�� �������
i���F�X����>6�A�T$8����m��n�s{�eX��-��������˾uFŗ�4=*i���_�E�F���C`�&�;�R�g]���C�,i:\�Տa5�Q��(u��o4�|V���VP�hl��G�y|r�n�%�y�M3�c=�,4��L�Ћ�����_����n��ܝ�Ni  2� +d� �F�YV��ɍIF�����_|�������5ʻ���ԙ��q<a��`���b�l+O'V�����Z`���ߏA>Lk�n�&�-�%���#�e�Hd�j��R��`���%����1U���Q�w#x ��I��WtA.Yv%��=�}�!�������{Q������>�	TK����枽��N	YyQ^�zռ3�W�]�$�,s��>����ck�Sv@'��0;1�8�O�OO�jDʛM����9]~1f�}l���H�� �?�T�2 玎:>k^��|dBk���?Eu����5�P�������]�/hrW1A|O��>@:��˜^|Ѽތ��	�oQ�j�a?�������0�O��O��CWw�6�Z�ĭ� l��y�� +dݙ�.��1%��O.��d8ݯ'i��ڮd�i�I�>-��詝u�P�]y�C/���18�zdÛ�8\ɦ�w�OK��I�T�a-#p��֟j�����
O ���ͥ�H�y�u��"��F��5�����]�q���zϺ��8��I�Oa�~��	R�TL��I
�}���A���x���<����c2/�: �s�`t�ҿ�3w�%\����~H(�]�"7�4���c���k��g��sN�؇PۊA 	R ��iz�NE��޺|u�FOlp4�ڻL�!��RvX7ƾ����7�p�nM�/Ķ�Q�d��\NA��JCkx���������qM�_�Ǌ�(��@����!MJʒ��_峟��?s5N��Mo�_�Ad����W���W_�ڢ��G�Cc}dR,�/�$�f���R��������)g�����&>��-�n6����G���稸��඗�҈Y��k�	g�pO��1�2�22�ŗ�F��H��;�������6�N��/r���E�*�C{³���3��^��l���	�x�z�  8��KNP�h�2�7�Ӛ���4�ӋfS�7eY��b��S�V�P<�uj�^��7;� @��ۏ3��ݺ0�al�����Ft�j�@ $d�C���;H�I�.���yP#����ֹaL<;�����
�����A �Aٳ��Q�{�8�6�a���<�l�,��3��$����&jVX���:=Gľ�G �4�;*%�_O: � =a��Y' ��S��Ӳ�Q�y��ȃ�܎��=���/� ������D��>h����)�7��)K�u���,1�c�LƁո����G#_�:��Dş��r��<	�
����l���݆�Y50!�ߍ�kb�L���1��7j���u]���O�+?u���u�Ո�/i�2�
�  ��䶺�����wo���"i.lJD�S��ĕ�r�$�S����уB���A?�Z�G��i�\�\L���z1�~���Y�@e��_-�.O��]�0���0�Gշ��c��[��yW-M����>���.H>S�?o]�ipciu�A��5u�T|G�)���ű��ջL(���8����8޳����=� ܼ��쪢�(�cl�s����%�W����OhPL>(����i�o��_�:������׫��  �F:�Ns�2�s�al�+Ϡ�U�v��6�&?k� ��|����jd����%^;=p�؞ع7�쪋�zNm�Yjӟ�4���H�W{�2I�Ug{�� b�����@c� ;�B0��X��� �!�v���>��鉵e'c{q��ț_Ȩ�^Oe���۬��4��HD�u����4ѵ�tu�k�}�g�s�v8�g�GT���я�s����!�ρ!#
"s��F�o���˷}:���њsAO]��,�,�m�r7��e�� �2�J� ���P�|���w�{3��n�Y��%�.9�#���Ǩ��������r��Q�&�&'�B\��;��V�>�h1yg�N=���\9u4�%�l�o���)���0q05L��ۊ�iE���S������3����bdh���l��f�A�.���[��m�|z\����T6��ι:��)�Gv�J{m�ȩn�C�U�ʃ @��l�/2v��^�t�.����i����������Y�׆�ߗ��NO�s��6�f^�k?$H�)'V�\������ft]2(�����4 ��.$}��/���՘����b9�`���)�n���_6<�,��C��<��y�oW���m���]T���B�Y�$U�W�6P���v^;�� Os6�@�h����{>k���s�ⷧi���?nv'��e���l�{�G�y(:ɮ��9�'ۭ�Y�[�t[�qw����s���>b��6�$Kht�r�~�7���뒄�,Wͦ���{y& $�eV�_K:��ӋW�5N��kXC��K�̄O ��i}Zyn{l>�b��q�t��j�L,�G��-�ؙ����S����_���w�}����DN��7cئ��b㧖��TwNp�Ҵ�s������A�8����ax�:N?ڿ�����=��mT��}L���N*(����*��������d��ᗏΒrD4����Ad�%�S ��d.dn���7����S�����M2{A�F��:��-z��X�s�w�B�U8���� RFW)����"�U�0ө&f�쾾�w�n� �S�Q�{+���^\�< 0.$5Jhsz�G�|O2}��0���c�Iv���b1-T����oe>A��Q1�c��PV<w�W8��F�!bc�,R:����eF��9�S����f�Z�s�`fizƀ������M�����7�N�D  ]@�D��0�GS�t�������n>4�TTV�W5h0��EN/^���͘�_�Z0e��;v�t� �2��d��P>W�� !C�d�A�B,���	���@�g�>��U-쪶������t ��l��`p �M�`�E�|�����+h;̗0���q�;��?#I�bG�+�A8����oV��[��Ǵ�&�JXTc��ڋ��ծ��;x;�A�/�#z�7Y;��J`�kE��nC-��+*)OF����o�/�����7��g~�l�a6�����uI�A�s�}0 $_������������V5+Ouo�Z2u9]��$�i���}ޖ��'��p�q�"�lk2�����x��)�'4F�-��qu���Ӑ�@'6_��N �F�w��
:?F��'b���z��8wd :�M��͆��w>'N���W;��u���1�����B��܅���k��<K���NY��&�t�a 6�G')�^¡>�h|8���23@.��� �pW�����FG	_�t|
����]���&����T�lʝ��U�uS��[� (�����}Eu9�B����g/3�|�:�L��Ak��ll~*:h�}<`�d�A��dPp�|��ӵVd��yNxl��Ixǧ,Ϡ�?�*��v�Il+t�Oأ�pԧI�]��|q�!����sMn+�M��� A�.��3�rLm3�S�m�$8C[uف��.:HK���������}FHM(Qp��O����D|� ��;�d��ع��v0c�$�WHS�>��9..B��@Axj����w����?����Fv���)ꥪ�]4it_��8Z�U>�n�����.������Ϟ4�N�WA�2� d�  h��̓�]��E��F�/s�<.|�U�:铤�Ĳ�O�{�k|�����}]��Y���w�~G_������oa�⃢�w��f^���sH�����cd]���	��]t8�o���UQ�݉7Dꆉv�2ٶ�ųf@�{b����x���!^�]l�P�V5r�v���OE)�q�qs�{�3��=?��:6�Y�0�>(�g3�T������;��u���^4z�0 ��2���Fǆ�\t= �  Ё0������oN%����%��k.��p��6׹���e�z5�3D���dR�TC�a�6Q����@0��ra%4��}���ѷ�N��v��\����4B�����I?�ך�!�m�_���5����S{�N��l����Q)�H�=��'\����+�ل�V�����^��8 1�k��t4���,J�a��m6g�����59P��=:R� &?0�H_�����F0@W�v���l�\h�r������I�j�#���}�Vt珗u���aV}Hd���\�_7������ۖ��I-��c�6⻨�Z4e?Z����v��v���̳�4H3���]�;2��8�k�kî������n��N�ѧ��ԗ�@��$m*_��:Ώ��ǫw�UU�5�\��ۘ��1� ���> ���%R�6AبM¢���	(/�]�in<
�U�ghO86z7��Z�����x[i�S��;��)��D[+�N�|g���2�,勺��=�]t,_�,�v�=�/e@` ��,^��]�D�� �,���ڷlj=[�����ڱ��o�����s��}:>8�/^���/��n>Vt�l��U�!��~J�ё��W;㏎�����I��g�B��:%t`sD�#���ۂ�]�����7�T���n�<i�N��BR\�̛�\ȏ\��Z  �yۓOĀ��[X�F��t��m<#�D���w�<�1l���=ȳbϦ������{���N���Z�V'���^�<��
����k��m��<�M������>������
 �Z�xHA6?6'
 p1�V�8�~�1ir:�)�H����LIj(:j���0� B�M-�	���r� �d'}���7K~[U�J���졵|�l{:4�ߨ4��.$w�b�w	�j*�h��sn��� R�aZ�����Nؙ��G��zCe쫷�X�xߐ긊��Mim������&	�i�AY!{ ���Γ�,�	˰�lVRY�P�F��%�z�����gCar��	C��8׊�p������'HC��}8��}j�����G�uҾ��`�8 ���
����?��}�w�ZmkQ�'�{X,������g�6��1��L6m�M��;�V�������F�&yp{ڵ�j}�r�WF��O�r*_Y����vD��⌟��Gt|���+&��o@۟�����.g4>�?g  ��{���D����ߖ����]���Ms-��������3�x5j^c:����,��arUE��A�؞�O�F\|� ���O��|ɸ���n��y��{@m���dɩ��o}�W9���L��蓕�_�L<���S(ۡO2ȧ/��z���T����H: 0���9����dW���
8�IP��d�B�^$ՠ�b��
�ݖ��G�w�`e�q���_�=�����i�� O�!�2qi��s�� eP�D �^E�I���jW�O��T���n:�(�)-hEӾ~�@�Rfj���j;�����ܟ��rdmE�L3� ���] ��";�����|�{���}3��?AYm�TpX��ZU����`�6�A
-��$�FNEG5�7q�[G���'��<���{��E�_��)�#���}peh�<�v�?�q��n���ZLi��󦹯�4*�9M�e�������iu�d>�[�}@�y1�s�:�c�$[�.�k�	��4��8�qWF��i7ҷ>���^��AK�����r����y���<��,:��i�];�Բ��Mv�, �F�*s�xU��/J�����y3^;t�;�9��齡�늮��$�Qʛ�<�)I����C8}���۫�>|=��  P��|���������#N0>N���l+������d��Ӷd����ݲ�<��3�����6p��藙@vq^,�[���{�]����E��v@e�<��V�Ǵ3iq~-��=�u���mH�e���d��G�*��gp8��qs���Ta_�в�z6���>�&Y[�]"���|L�߃�/��>�|������n�e�t Ӛ�ή����ss"x M��v�����/��o>�?Ey�<���1����.��{�h7R$���dWTU3>�L�}m���r��F�9�1Q͌�T-H�N�4�T��u�Q�墺$�,��i�\Xj�D]Z�ڿo�SL�;	@����F~kZ���Қ�ߪ���ET�'����w����7���o�,�o~���Ad���6���/��_��?�����?�'��OWYa3(}��E�<�͟��x��5A��8ƀ:�'��!J���6��w��n�{p��H�$R�ZU��O2A_�9�}�d��D��`ˌe0�!�v]��q/��5u����j�c_���r�����*��n��{��tżdwN>?H$}���e���(Ј��!2Ov3�w�Uo�fJ�� ,P�傖����M�jF��f@��T�A��A %],�蛌F�F����uGb������͇������;0TL�FOη=Tc��	���#�|3�T �8�a�z�(���c@l����?cQk���G��'x��v�G>�M�-����y��O��$�i^w�r(�ܞ�a�۞V�Ysǲ�?>:h�����r�#a��:��Uc�Z��]��~�剣�OH͹`��{N�WRї �����!Z�K1Rp�` 	4a��'$�~�^:jv<�{�������&�;���K��y�؞�:hۭ34ͧY��'��Z�M�;֔e)�����u�\��1����Y��1�"�c�N�VM�a�����2_����׶�}��ub���{��-�e�����ww�6����r�z������w���1ه���-�qI�2� Kd�   ����U5;6'����|�;����㤞�ujL%�ĽZ���I4�*ն3>8�[
��-g����V.��{U��.Y_n��{��6���UT���⾎�����E�#��f�ڴG����p/Xa�(:eg[Z�X�Τ��P��
���ڝ�hiLx��O���r<Z�^xv��6m��c�>��R�GV�P���v�����y��&�K�~�҃�z�q��k��7��㓌�_�hr_3���MA����I�h�B�ڟ©U���򣔎N3:�@�~�i �vUES�mS�ǒn�t󡤻낦�5 $�;�4� �'/2:{9� g/rdi��>�N��������.���.�o�ӓ�k[�� q6o,��/e��\ À�S�h���`�ˮ�6��䓑Ey�<�s����rx��|����U�+�vo�1��m�L�U)k蚝�Ξ[�����PI���G)��?5�;.����P`��e��|��٪h�K)�~����@����>	��~�{>���~��=efe�Y��_@��l\�h��������ħt&��'�~V���� >�t��9~���z�x�FHML����H�A �C�J�= �RxF�QrF��Q��W'i��)���lJ���Ad�9� �eY���pv|������:{W۪N�c-�CTOa�iS�dTוs�[�����ɓ��bF)_r o4pO<5;�u��#�[ W���	�x`@L yj��>M3~��qPKUHY`�T"U�냴	�]�Ox�>���m}^-��WL]������y�AH��9���iӹ��ׄ4���f�o��iW+b��k�H��A���*f�� ���'��p���U�h��k߾������@d�鋔f���o2�z���c�|nt�Զ��Q�!@��;��Ӵ9?k6�	N���R��|,���iS挙 ��fC_Vs�֯�,P�_����eƑ� (��u�]���S�\�J�9��1x����(��L5��|���ϖ:p�<�9��0U��Ȟ�x��
p_U���}��y����QbC���D�� �5���V����_oU�f��0�,�*���B���8��5��q�ѻ��硧��Շ�/��[,�3q�c�@4�.���6��>dɕ9���� �G�H��;�S쾻2+U��T��L��L�)�F�`��>� $��؅éo��zR���f5��}����G��_W���c���^=l-���͉Y��a����񀞹b"���B��.9&��?�O�;o�w��j؏��ЉUt���������l������.���"
�$�Qp𨏢���c�x��\��Y�=����m���E� �������2�,�|&�;�v� �[;h�K�\��vRd&�n
��Y�����)d���^  I#����������*��q����X�S�q��UU�sD[�/Nu,Ԕb�r��d��FY5J���+K��I�։/��BUG߫��A�+I�rY�L�~ʐ�y-��J�Iǁ�_
��c� �U�\$�!�<����"�k7��~�9������A��o�۴E~k��Qt�:�Ц��S���3�OH�aXۮ��g����Đ�FG�6�RuBdL�z�gnA�g}��㳔�YN�����t}Z�����-�P`��ɦ�����.^�t|���(�q�����ջ�>~3��E���� �h�l�/2z�jD/^���ň�6���
PC� KĬ�<���Y�|RK���g�Y�C��Ua��t�@&�'t@��AV��%����zx=6��~�S�>�|�ͬ��dw����#������?��TL��fi�g�M�:I: ���-�U��$�f1����0�S��	�����.���cƇ�L���,��>������o���5$r�|,�B��$����G�2���,0¼�pړ\+�u"H��]���ߍ�� M�l"6h��\r)��L�:-�f`b�cDv8��<�L*C�bB��Y2�j4���,3Ο:�d��S �����e�����o��_��]>;�&e���K�D�B	�^l�����k�^������)�d-&�?Q�p���]��\�"�"�'�����%�&��'3$!��'<D�	 ˀP-�@ޡ�oϱ��@Qa�U���#���n:h9ש�ڧu�kk���ջ��o���|�q�hg�a��E��{z[�Mu9gײi}?U�[�x|�F�~�ҳB{B����.��AF�u�C㣄N�R:������S8������X���SE�7�]�twU�����&5L�w[�͇�>2���STe�[�,M��t�/^7�W9G��)%���M]Q�j{n�+]םR����YKݗ��z���]p�&�hRA�/)���.�p���}r���g��<��n�����:�z�R��l�C�Kl[�}�*p�)e�4�K#���֋����m���>a�ha�0H�n��hp�1=�5�ս�v�:�d�������ƙ�� �OR�u��9�52GCLI嬦����* 0i~�n��F�c�����Q����p6�a��H�Bh�;4�_����U{�����H�>@ �Ԕ6��n����u͎��Z
;2E�
2ru����2�kl�W��)�7�X�H�[0&�i�[����[�); ��+������A-IRԆ��.Xn-�Tw�����_�������[?~B�>'z9�Ad�%���Q�ǿ�?��n��w����W�e���̬�����<|�۷�[@[��2L,$��el����H 1��0�!�����0DB2B�Z�Zju�i�ݷϽ��=����o=""��jgծ����Ժw�o�|DFF�X��o��mu{ꭷ�m��(����&�u/��a�I�V@v��o�<�����Z�@8��)��@���iɀ���"�ZK`P��пxEt� . �~=�d�s�
���>���$t�I���|e|�B͚vV���:=���ݰl�*ˀ�7�G��>�50�?fj?�������̉����2�b[GY�x���Ztj��v����c3����6��);�{*P�_������L�2*�@ ���|x� ����O�v-?�������g9Q�_92�M�.%�_���8ʏ]v�L7�G�^�}x����G+�ﾽ����k��_{0٭���F��'Pky�'�<����%M�}Ę��-���?9v�� xV�J`��h������X����^��N��|wh�x��YaɏP�� ���(���+IJ�ߎ hr�rY��&Y�I����@�Ĩ�V���r��7�8S޷Z؉E��`  6�dS�@�o��H��������$��1�.�S�"�|-�wŤH��t�_X�+��;/��}{����t������s?=9;3����(G9�
�7  j-���ӓ��_���T������E��)�XI����9UqR��)M�I2�x���������0
F`�������U!+@�]6�rq��R&A����?���}�x�X�P�:kS�/��Z@.��k��m?G��Xg9��o�+".��E5��!����i���G�Ϸz��F=n|�T�(CO^��꜎�%���W�&���-�i`���Ʀ��ߙ�S����8Y� =UA��Z���\P}����GcgN/rs�zd���,����**@l ]����5� �i�AHa��~dp����K�A
�|p�Q��嫑��bl.^@f 9}����{qT�~��E��oW~i�:��o${x!+��!M����~Ԟ	��I���(�*��6��V��}�%��:i���3x���P���q��a�n%�� ��/�n�E�u;��	���R��ݵe�O�c]Ҳ�����8�tY���+>�C�����9�x}HY�;qǷ�~�Y��?����5u��7�D??��f����B�u��Jտz<|����`W��4�#RO�����n��?��G�C�1���U���| ��i��q@���7<�S%,��v�v8��;�M�W��?}$���V��Q[�PJ>Ѝ��kf���ą������ 8������h6�}��$�>����Jz�G���æ���/{��:ٹ������I>b(��JMe�yBv�I��v�S�
��=�/�h�C2�)���s��q��$K�
���f�K[|��G�*��ؕ�m��|9^� ���8J~�ɭ�����k�����̧�ǳ�wo/��o���W��:k��\n�=*���(�r k2����v��;�+�?����2˗��u�N3�u3FY����G �]:z���Ԣ�� �4߅ �փ�~验�c�#ٴ�*�7�&�E��]R;��b�BӮ,3��v� �<���Bl�N���&Q���Rڇ��YS0%,�r�1�n}�g>��Ό,lu��镈��X��|������sW�\�`�xu ��D,�r�^�y����ӺZ���9`�߇�Yw�w1��E4�/F�F���7��NQ����A��:� pf�@���j3�o����"��o�y���3�W�}�s�rD����2���3ÞZ������s���,[�c����u����|Z��w�d>l|�' C�*uJ�n:o��" l�F��q�=,���ϼ�R�f�(�F>�	w����Lbqb��zuy�_�FOzNf��ӿmrȎ��iփ�H>�� ֺN�ޣ�JTC��g׎3�����fk�'�뱺�B���Dc�vC=���w�<�2�AҘG�~b����y����_�����e�i_��(�[�`�\�_[���~}���_�h�I�Dcզsep|��b��%�z�l~��+���w^��F�Ej���Vf1�L����%h���w8�d��UN{^$�s~Y�'~j}�S��Y>���V�ҟ�����w�K��H�4K[���1�tTk�cHF�R�Y��Q ����*,�J�$�e��J��ĤRb"���즌��F�&1�Q��%iF�~�ɜ8^@�<O�ȡ��&t&1�4!���q(�S��>ĸ�g&hA%P�ʻl��؍~�g�R�	 OǙx��e�  �O���v�e6�{k�ܺ�S��"v7_Kp[a���c��ʞ�J,[��WU��wP�{��LH0�ܯuA�����������J%ԯQe���J�E�6��j%��9/ˤ�Lc\VU�ӱ\�8]L�ٚt�1�y�A��M��1�����cYR�`�VϷ�_��؄� �^��(��lql��?����c�|�  �r�zA��P�m���*��	�Hh�j��O^�[�5�7�}���A� v����	��+Ԙ轢�|��#���ma޿�������H��h�y_U�/����R>�\p�=|�w�cd����J\�(��yN� ����CV��зyhэ��o���w4���#�noȤb��ӫ���5�9��,kty�T�����m��~���Am������u�䱗
��3��`�7۝�̄l7od��9�9�E��sC�$t�P&"��3q�����s����>*���'`��)�m>1��Ӗ���QF���Y�Ϛq�~��`ۙ��o�u���0衧�m�3H���RC`U�����U��"�~�$h�����t��X��L��C�n���={�����غd�6�n&g�F�Ģ}5��d�[>�g���b���Z��ݡ�V|�����I$+�I&f�ߛ
}*�"�jEg����L��D����T�� ��|�&�����#���u��?X�ּ�M +!�g�����=��x���e�C��u����1_��	�	t��iI%PV`4b
r\7������XK�4��o��8�AyhDJ���,I-�D�pս��$v���>UP)+r��R�G?��_��@�SI�{�� �ˑi8�YN'������1��o��ލ���ϴ6jKP_��'f�X@��
@��I@@z����{�V�>tT��$d� Ʊ�n�!�l>/��s{�����/*?k<�TG�Q�r�C�  �Z��w��g����j6��/2kA�D׹wUf�2u_��W�x�F,[(ʚ��S+�U���J�er�L�\��@�Q�w@�9m�dZE�����U�Ւ�yig\����VV��{2��m/6.R�t?o�nL?KL��馫[��.0�Rf E�z��O��T�O��_��4j�k%���r�,��6���!G�瀱��i�O2��q��t�ѧ�Fi��JP� �g�n���m�n��GӨ�x�_"�_P@���B e?��G&�����ļ�rlίGf|�'��e��G�0�[kh,�S��>��$�G���&���N��~�|�8"'�f�<�W�3��#��soV����:)8��K�y���$W[Γ}�M�g�����|�7Luz��`�X�v�����{N=�gϼs�h ��s�]幦v��w�z9X�,���>� x�rG���m��ؐ�!��Rƪs��_�.M���	2g®��v���p?�9k�y���\�9U1�1P�v�{�BKg}��ГR�_��<��ݬc[��Yۓ�q��� ��������5�'���}�Qe�ߜly��"�U��S�o��ά���5�@���9�%��V�v������7c�'�"X�۠(�B�����s��[�{k5A;k�n�k���:�7��uQ��JR��S�P���ѓ/����e����Z��j��b��T��UΙ�й���,���!1�>��ѽ�緆|jܐ���-���]���-�D���n�l$��nM�\ng�h+�0��RE`�M���Od2H���~I�3��TB9�V�H����#+,��N��~��z2�̸E�x�:��Vb%�^-7��XP�f2�������>?9y9-�bf�{:���(GY#� @�_�~9����_��o�o��/>޼���bDa���ֺ�����%���$�?^>*�� �e�.�S��e��ƕ�A��~o�@2��.F�[e��3�iuk���a!A-�JjI�(�L��
r���|&8�u��U@�� �"��E�g'�H����RTdh��c&H�6��޴��>�|��\�1�9O�lpF'�O�����ڔv��f�V��GvD �,_� ش�l�<�\s �X+�O�LJv�l[��>�-�#���RaC��<�E:���{��bd��<#�˗���0"�����D]���	6�X:C���8=9�	dp�zd�������Ϊm���̹5��oK^w�;K��8��nc23�����s��Բ	IM0��U4}L��7:�sf�Q>���nrf�,�9���E��#��x��
�y
%2�c9ͻb�Q�S�U4�o+ÏLz�D
v��G��F�Gp�Z��*
Ǚ��x=P���DW���d�sa�5�y���&u+��O�u����(�Y�6�r���\�X�1��$
\�Xg=I�l���\���0�߲?L����4g�̦�H��n�	��	���/�,P���>��c��vu��!Vl�	g�OX�a���s(�}�l�!6n���M"4䆓G轣�#�W��Π�����r��~*�����>�h��$���]�B:�-��a���O69�it��b=s�b�b�¾k�Պ��ug�.��U��}{�ֽ�_Z�6�@�j13��V����Z�$�QvO����kVd�� �i�1}�Ko�ⱍ�PQ~&� �aPm9���q��4U%v��9�E�aƼ���pz[1�`�bϧ�By��r4b�J:/S�^��G��?�����uҠ{H>	����L�����n�@��6�U� ���rL>]���1i���qZ^�6u���6� ����Zb)>���F�������9�b�4|j���~l�5�Ͽ��1�w���n�[[����r��e�����y~���_���������o���-Q~07�!�x�|u(���H�3��r�TDy�ē����]#ۋ�un՘��9�w)4d���
��`��"�1�t1R�5���'��aYrq���2�/��T5��� �2
��w��BoLjd�f���k�[�����ވm9��O��QCs�mϕq�M��,7病�����ӻ�,�L��'��n����`]���j�Ū*N�`�R#�I�	<�����[��WV2�=���ϟ߭�=��F�i��&�w���R�Z$XLl%
"�8B)�#s[�j�ͧ�XZt<�+.����&�acH��������/G��eA�8f����k�K!~�G-I�Q:6�	@FC�ǥ�}��	�|l��_u��9�5
YNvje�'�A39��/JatXл=� v {��>/ښC�'�٪k��%�!�s����':�Xa��Fv�/@�ִ�w�9�5?Eӯ��&����A]����ӑt�T�ȥ~lⰊ��
��陣�5��̌�����65���ˁ]�O�x�;�By��TpD7.�~�:�������`���Fc�9�ng��dw����Ě���y�#2�XQ��� e����A�@~ͥv�`O8ѷ�d��7���F�WIucҶu�}z��ޅ���	�U�-�?���Q"�U�ѭ[�`@^˚�z��4:�伱&N�ʅq]�L@��z���iJ����7�*)7�7�|�Nd} ��|
��'@��߹l�����@u�{�f�66�	��9{����N�Z��t����G�������ۦi���|B[ɏЌ��˜���f�M���� c�|Y�1ڞ�]�_[�����o��q�Ij���N~��]K����❶e�¼�
۵(���WʰW��ٮ��Z���CD�٧�&�F�?P� �ZY휙ݗ���@��t	PA�����n�T�ך��ͤg2�?9I�Q�ǰ>$BE�>�������;ϑ��?�7�$0�vĮ�Š�����_86��Jۖ�_�0�傯	?f���,�C�ƛ�Q4�ڠ�dBm"; ����v�	��t�y���{q�J���$q���s!$}���<9����������ח��99Y̍1�>w���e�  P�@��f���������O����ٷ����1��;[�,t��\�8�մ�*?zB�Mq���"@4,-kW)UR�Xt<S@���X��m�v�@�b��D����7FK8Ap���P�<{�����]�6��Q�`���4�6]t�,�؇颜�w8���c�}��)bM�MF�����g�ۑ���绗���!�� �3��)�Dq6��@��7�"��T��a @��1m�RTw�j����q��DǢ��Q�eV�&`����ظc':Sذ�����>L�_%�W�U�p69���4���F��j�=tI�Y�K��N���9�� ���4�3uY-��Z����5�%/��X����e�oN�l�qh%N�U�����b˭��j?DPJU�0F�:3�gZqP����JN!h&c��&�����@%4�ElgG�k�M����+�uo$C���UW�S_&&�z��[���s�Y:9��(=��s��|j�=���T�Ʒ��5�����k&�{��Y��̿|52/���W#
�!8��T~�_���/-�ˆ��1��F���@mt8�Z&�=�/�5��XK8x*v��񺛞�LTY�yx�(H6����Ȕ�*���;b�2��+Yt���e뎲Oi�sl�#ϵ�N����m�v�a�ɗ� �+���THU���N%��-dKt���'�y�9ۈ`��dQ�7 �࣒m��l�T��w�D��U)!�]��5������УE�c=���L��.��Ecǟ�3k�`{�)&��Am�1���Z.�:fl�}x��pq|�kڸ���xI>�����h'`@�0xf�m�W��sf�;9/�O/} �;t��^��fX+W���j���,�#V��]��:����فm��v�4�\�s:^/���/�   ���8���s�Wv���ץV/��>�ǐ~͹���d���0V,�	���'����9e)9 >CT�L�Ϻ����\7��� [3B2@�+���K� ���� �]^�wK�O��o�[3�+�Q	�m ��䌓�Y%`��e��a����	��*i�ƒ�`W<�j���Z�����Q���5 �T9p`l%�ٍ���e�?��B'W��=��}���=�ǹ��x�;	����r.a(�kp��1S���ɍ��r�Ĭ��>'�=M��
�5� �Ϯ�5�s������W��P� @���*AS��������@~�F��v�O������|��ŷu>�1�� 8�Q�����|����ﾛ�i=��/Q!#����ȚNh=j��{� ��.:�Z�	��K�]��`�k&��*��o�Ě2>������yA��3U�%,P/����[O�7+֤��b�F�7����보��|�t�HQv�,�|�y��Yڏ6�Oj���7��v$C��[;�q�2��Bc�v���?�A��Ħ���0�KC�e  Lo%�O�c*s�A^8�˔6�'�6�Q�Z���nƛG����NyL�h���8�@��k �Q�C&8�.6�h,
�nŦ2W�謝f�w�f��c�\�s�Pr& ��,��ؙͰi�h�gI4�{.'���q�넆�Nn8c g7ee�POp���G��ͥl��� ������a�ʢ�W�t �vr�������+�{�}/�'/��kd�9.�z��ku�i�d:r��o��t$�V2QOe�\�c��	T4����X�c�^��xBժK�8ĉ�}��5P�/F��ϱ��7:�ŗc��+   ��\��Q+�j?
	Ƃ%�n�S��^�u>��a-A	0�`��_�Q���e�����Ǔ��9�`�Ν��fvW��j�
�@ ��DQ��Ƭ{��68�ۦ�Q����S�y���l��d�U�
U:���>3��,��iNپ(�݋q��z>�����a%B�8�W���kuh�P'(d�Y������{�[��Q^����qe�#�����s�z�ň@�h;:��ӹ�A�?YQU룯�@������`2�TN�U0 ����x-�/��Zo�x7���͍�`�vr��#�:����	��ňi�]B�*)���������V3W�`+����`�e��f��eMȦ���=a'k�,�L1�Z�E������-$��BKz	��k �����2^O,`u.�`�;�b��� ���M�k��%�J��Ƣ_�Q2�W���K��2���x���������ѯE3���ڄ�<��k�sy-�57��w�s9����2�b�3��af�ˬ��p��㢱9Ic~��k{К:q��u��4go����UњJ%��~�)��ϻOl8φ��s�m�����O��;�w
�јK\�����,���2�D�>BG4+?m�M��	Ax#1�\+�q�OJ���G����A��CN����h�D��l�1��{u�j[(�#d�.�3(��R�$�Y+q��Nl�ůB�5�Y4��x�\dVx�EK�r��e� ��͛�����������������*r��9-Q���:��D��{Z�A9'��gr/+�u!B3Jߚ�����4 �W��L!�п��E��#��D�X����L������0q>��"ۺA�Ѓ	��-��gk/��K}���]*颜|����!�6�(O*^X�i����F�޳�����}��FPc��@Y���㋕��; !��#�3��@[N�3v� ��'6�ӛ�~@CiP���XL�D٘��sOl��j�i��]�zv�珼>��xO�RU��f�|�07oGf1��ymR#_ѯ>���Y���;
ؼ*(3R)� �����,_F6Q@I/�1%����m��P��p9�v��>���dCf���k�PR㢙Kp�b]�XF�1vA��?��G�˲�����A��;��+��!cB�"P:����T8|�{��ȼD����h�8y[��\�&?CE�_��I�?@5��C�N�2r�+�z��u����\�@TN5^&֧zړ���КI}�3����K����@�|V�.B�a��^ӧpD#�{!����"�a��f8�s�i�#�[ɴ�\��47���vY�c�mv��w*����l8~��#6L&�*й�],��/f�+A��H�V�]N�*3�V(ܷ����]V-�!�N����۲L��+��knKwNb\�NsY��\V�3PA�>�g�%����(�Ϡ+
 
U��=������1kY�"��5�[�M�b,c}���������6{M]�����8�,�e���ʭ��#�U)qɛ?�k�����@w��{t�X<���)�'�7lm�o�WD����F�=���?���˹�������=��W_�2)��O. �-��&-�R�N�m $��~=g��+x�d���`�9�r׌׻;C�P$�7����l�#et�EvV�5&��#a�[Fn��~M�t�ez}�X�r_��G���W/�['�嗬_Q
 �p���6�v�n�2�Y��(J)U�˻�=�٧��f\�s	 ����tX�a^��}S����2���/#'�HN�[��i�P�m;�]G��$�"�c ����0�#c�ÍlG4�����٧��6�>_�u_̼��5%��	Kk��b��Z"�τ�����5���Z~ ����1)���'��"�1GKZ�n��j�U3�ƹ����9v�X���r����+ �{�X7
i���o�����ͯ�2�pq���*lZ�0D��
i�@D�>�$�E-
���'�H$���F���P��q����`���й��6I�q]g3�����ELƮ��NX��������(�����K�E��Lw���E�u7�򉓰u���8P�&���c��-��o5�AY�H��sΠ��r�5k��Eb��$^�Oc�3@�mbv�Pz��k���mv��~�儃</G���fϪ1�7n�vC1#.��1Jvd��q�Yv�L��&Փ��FI�ob4��	t�L( ��(&G�.\6ad��*≓�v��R�`WA��;���D����\�}p��x=nށ�:{p@��4Oe넚9q $��b ��r�,�?2�@D
ݣt�[����l�ܑ�Eɑ��ﾝ�7���Ƿe3^+3�s�6צuއh��E�gK
*�c���9�3�}8RN�K�R��J,/�q���tS�Gxuv%��v�7�?<�5v��x���uD�Sv���({��fD����cx��ȼ��'��W��}��R�rfN��V�`� ���������`�0Q_��Q,���X��|�3�;���@��#c�)IYRִ����[Jv;�zJ}��Ȋj֕�� 0v�A�z�vÔ�O�ߗ_�QaB��>�kc��ղ+���c�\]=�}��c,[�̱�-c�A�)C5� t��5�)�:��H���w{�ӱ��K�.=��pd�-�SY�]Ӎ���R��.5��LW�u�^��ht�|L�0t�Y, ���F��Û9���1jS��cY�_���`S�b�S��i3_j��Ĉ'{��o�H�0��}���&~+�i��aj�F:��U���o�����Bĺ"ޔJKo���.������ūB��G�D��3"�
���i�1'�nB65lwɦ�?,�����2�}��1k]%�l�&���6��-h'�n�񜘃'�	 Yb�=6Xˌ.�6@#3���Ʈ�>A;XE���x�-�g@��#��w%��
kO%t3X���T�KO}ݐe�'Ь�[.\ބ���/����*����R���I��4@ �����ZL��H4l�[ٟ�����T�B��1����W�\U�3�1/$�% �w1�>�+<��������ZlC��� � 9��Wc��'���� #�=�}��>�E�3���}L�b�t<�a'!~vz�H�Ϧ�>"���c�H*p�s/@f���.HO�ߙ)fBk��=K��}� 6�����
Crzԫ��>O"��W��|��n`l�6=�i�>����4D��UJy��آ���|C=q=�m�jµ���1�͵�#Rҹ�׊���˂��k��jԾ��8$�$�[�=� <*}e����d����U�(ں�O弹�ޏ����o^���?�:�rt�Le̳Ow:�Q��r ����������������#�Һ<���z��9q>	�����jp�@
��1&��\���B�喲�J_��t5rm�1�����
<�\'^m���1p퓺6��\�I�;.��l$f��׼L�d��H�A����)����'�I�r�ԛ ���U�Kp��B[��m`m�c�˻|P>gɲ��evq�PI|mx;�gT�"���e�.�&(  �欘��"�;��tL��꧱���P���5g�q�#�t8ˁ�FF�jI�A�v�j�-isOF�:D� Q%9� J�Jkӱ��J���EK���~��3'�4���zr^�A�l���j
VA��!QW5e���3�LuPt�ϑYÁoK�z����n�#3��A��;�߾��] ����{��I��
�����Â `����\��{j}p0U��:�@B��ň�r8����3�e#z_�)�$S���e^g��Z��}������ۛ��	��8м84����);D1.3����0���'cs�z�ԙ�YXR��ݏ�5K�V�8(ǙI9g�Ι5������u�_�ʙ�d,}Z�p����=h�h�q�M_�S&� @ت� 1��l2cr����2�y��c	��oȒ�:�r/X/��	���tA3�ͫ���%`��������46!6�u{���j+h�"�)@*� ��,`��T���� 菻�������X��͇�H�)��r�+d����WZ�K�\Z���=�x4pk�˕w���`ˊ`�\+/  ��IDAT���Pb��6A�g�  �#��Sag���%3��d��#g\Q	}a�� H� 8�3�8 k�쾤�bi�㵱}A���9��V|��yFC��U�c�% ѿ3���9�܂�^��t f ��ql������?^2�e|V
��r6=����|^04�A@�w�z AJ�;Rm!dC�y_w��4�kh�"eH��}��Q��c!֢��0�,�S�|��/��|79��u���������:^��/ۛ~5q��R��� +�=궢���K�?Y3.A?-���tW��tUF{���U��!����Dy��`�æ�*��/)��d{�C��q=�=)��)/�Ԟ�Tb6��$W3��TC���E3��f����\��&�� p SY	�}�Ǎ{��ȱS7��$�Aj����i�����f;?�z{�D�}��|����a�m,��(�L�y=�꺙�%Mj��IN>	�(��C�h�A^��ڸ�$��5�b��D�W�-��>!���4���j�>�3i[��S��� �r^lZ$�����
[�䛏��������_�'��_�ξ�N�����9��1�(G9�QR�7 �����㟿�ū���(��Ic�5V)ܜL�d\t>3%�(�TɒhpXԨ����Y+n#h+˖����ubXLd	���Z���b'�8�Z.�:]��͔,R
N��V ���x��8��G&}D�/i�&H6���L��>^O���,�M�ht?�߯bP4��Z�1��(O,2\S�c12�� �;6�J#� #�R�i�d.b�.ǔ���k)��׆���(�3��a���s��a�y�  ��A��`2O �h��#��`#T�R�7�L�@�e=o�w��ܵ�(ףz�p�z+�d�x��p]c��\d����X\2�5��x�1�j��i%�69�U:F8o螲y?`���ECΉ�N������K����y�˙y�y�휜�`��ӉjZ ��L��ԙ�M�d�L�Y`#�����BB�T8��:'��8�(� �D� ȹ͚5�����0�Ozz~Mw+�J��D�|��p���\�8��/0?_���O�GY�M��y�~�C��{vQ@��Za�b��L�9 ��S�GBS}I�]�\�{��q�~�[�WQ*hrb��c #�Ȉ�@�knĎql��Z�t_�u��ਓ����O�U�%p������q�R)hmpʵmt3�a�>W��!mZ7��v���F|�l�SV5�\�=�_0�1�W*�5���w�����}WR�*e�G5�þ�]�  ��/e�;�h��i3��1  Y�*6ݓ����sdÖbۦ�=�8c���=  ih�f�R���Q��u�8���/��MEc�,����Y���t���Â�s(��6��ǫv"�W�bݝ5�n-��ɥV�<�`��욃��uqL��`؆�"",v�����e�VN3�)P̓���2ԛ=.�w?.����/�y��������]F��˘��]r�����]yg�s7� ,�Ϛ�Z����.gĚ����%��>�a�z���.��Ƹq���g���?c�&�c<�
�r�ۨn�]��݇`�t���=�7���7���bD�s|��]ڭ~�1�m�;�j׌�j[�˷��h�����'��ko�z$%d�����H:���a��	�0!��o���w(�>��$F/�5^9�/�E�؎�?��xN~�b��Ǌ.��%�^�CL0���c@�H>��_`H��- �O�����Nz�p-�q"eM�K]+t;�@�)���u�h�[U��h�I��p�g�jԾ���������={������y��?�ӱy"��Q�r�OG� �����ya&uUMjWg���eA;]uH�a��4����k�?�|kU�ӧ�g��2����y䨓QJ|Bz�_����Z�^[*��i��Yr`�:.��E��8% 2ɲ`�"z������恾X~ʦ��U�����G�����kF�_
����C�h�-a��64z%��o�E�F�VI�@s ����/Je�N�bC4����8 ��� pv�w
F��J�ubH�����%��ngWJ���lz8G��O�%o�ar�4�w�a�c��{�W������{5�Z�(2�����I����ē�!8��<�/��t�c�K�xB�*�sʶh6�7�Эr0pfi	���O�Q�� #W���D�����3d]S{������E�d���L������������pJ  8��X�Q������`��Ir�/ĩ�z�O�Z����A������N�r����6�Ef��v4.7����_W6�y��cƯíX�|߇��t8�VW���F�"�p�j�S�z��n(����R|�Gj��ՃĎgre��j}w�+�b�)8��uh��c2��C�������B�8�CKL$XW�/�~��}V0��	tTӯp�+��.ǫM��̓׵���7S����X���ɸL�U>a&'Қ�eq'Yhv��κ���������T�T��g
j�s�n����Tظ7�����4�93d��s���i�[�$x�����ϙ6�䱝K�n!�H��>��X+<�� �l�IX���D�8�}2a��`o.�V�3�t���C�Ć/�T���W���)gM������/H�����r�,h%�ծ�:2
H�x��5��b�VR�.mΧ\� ?x&0!D��� ��օm$�����O�?�������r�^xmvW��>��E���aFlb` �@6 �U��6�@rf9ZHi3�;��^����`<��XYުpJ�p�CA��sկ0Ny�B�X��":x���(�P���_���c"��FOiV;t��ht�P�k`��x*�]�c`���]b��,6 '���y#0�	������jui��K:��aqn��q	B��!����Љ?A��}~��/�:{�@@#Z��������{߃^iYsݖ��<�ϥ!kd[>����7����v��,� T��[�\N8T
|�n���mO����\7�\�ɾF؛�&u.w���t��<�s��{��>���:#J��N�E9�B�3����`�>��X�ex���T��̹QQ�&g����'��|4�L��u}����C  ������W��_|�}Y7�8�e�6V��<e�kr|���Ք���1Xo�/�'���"�)@d躔^��X�����{XӦ�qJ[�LP�z�.c�i��R\#yX��=���,c)��<��V�n��
���)��Y.`L `�$@گ}M��Ӧ�1t�O��[/�so�X��x`	�gM���L�Ͼ�ڮ9�\K����2:��X��6��o��*#F�$��1͍�6��{v��������ƾ�b[�l�^��8{�6�Ȝ>u�	s~��稟�?3���n��T�l�Uo�Ƹ;�x�qu��I!�'�h���� �&����ų��% �AƉ8,וW�H�1��h&�:���a�b|����?�M��r�"["|�j3{nkp���ռ�  `k��xĵ2)[ΙB(3�y�h��dz�GHj�3x )�f��3Ko�Yu�É�l?�cʞ1&����~?��Pu�u�r։�[�ڕ��\b�j��1�7�	�K�8	�y3)]�5��Ƴ4sy���sϘY�e=`�� T��{�˔R9]���Qv ���j���;��e��΅�
��-X�n�r�
���TK.%m��f��o?�#{��v!XB��ok3��&�>�F�\q�koD?ϴJ�ɐ�X�2c�l�Z2~�W�$�����{��j�	�U9�a3쁀�݇���.��`��{'��yEǵ��������ee���u-�wk�G#b㡺�'9=c&�^e�X�x�E�Y�j��zFz`6>O�	7�*3��i���	�[I xgA�ǈe@ �T�LX�׬e�����v��궃���8��w]�9�ϛf/���G96I&��J�_u�Շ�'�ԯ��ʥ6����-*O |�K�5:�¦��i_{��2��re6�q��կ�t�*��S1��],3"����j����'9|\��>���g6��o2���~�k�.��Qv"���o�����d�������!��H̤��	���X�jlyF�j�^}g�J&��`�C���k��Z3 �yZ~a����oM2u�� �*M���Y��n;)��K��Ŏ��PU�}��9�����^�?��+G#��G����(��  ��\�^�K�v����߻}W۲��T۰�Ԅ��:*Ь��������P��D���(`��c�k`�)�,��k	��Z�ܣP��E#��i}\,�[c��F�&\���tu�5ȩ>T
E�|]��3��?ݮS/�f���b���E�M�L���>�����U$B`,���7]��b�5�����%~����8�6E�B;���t��s�����6޴�ܭ<��U������s6�ȶ�K�lQ��%�<g���.(3���,G�S��ay���1�=�����x�' �V�5��24䇎���]��=wMkӄ:��@������0N)+�b�iȀ�i�S�I�O�{�j�s�:�1:3   �;��!֤*� �џ��<��S禀�4�Rӷ�8�1����{tm�z?J�c��JhG�X�	�m&5r���\���� �����j�a{[*�|n9`�MO5^��W���:Ӵsi �]Rz�(��룇��G�
h� ���4��Cv'nV	8�$[wE��?��� B�P`x���Mm�QE��SS{W�T��K~���L�ֵ# �=˥tQbo�^{'���}����QK�0�,�[��y3F%ےK�c��ޅ�۴�Di�f,�sG�ͤ�+P�Y�y.(WɨN��q���K����~�|�I�W�F~����j!���h �u��X5�#��8��s7u!��}���G:��;�}���,����x�������N|46�x-ҭͿ�e���:��E��`� ��nZ��5/��+�-s�?���PГ�d���C[0�G9�3�m�H?��<x�/�*5�b5F�q�Rg�.14�uj@=�Oq퐼����4��(`�	���=�9�$�|i3Ǌ������|���R뒄K>F3��3��c���O���k�2BB�� ���&\g��������v>����u1M^�Q�r���ʾ dg���/����˟���?���?���d��NŴ�'�����dק��he�k����5��㣂�}P��9�qb�k!�At} I[�J����.8��������@'�ɢ'v qꢓ@���9�~v�N篰�5���͆��{n������)�f��&#����mhkgP= ��I��rm�Ԗ�3Iz�����~3����y:I｢�N67zl)Eԩ"�t���'tS�N�x��l�4����Y�U�v��u�d���f�����7�J@?:_dB�I�M<�ѷp��s8z� ��l������C%����! \6�2���p���-�4�jU�?V�8���纡L}�_�����,��pWT�q���&8��0l �"s�����Ts<)�h\�<��"��s���K�@	E.���g�J;�{�b��Jh*w��j�S7?��g3�V�m�j;�O��)����aЏ#���P��Tb��6=�S��B@]K� �(}��)�e��%�P��D�:��+>�tJv����x�w,��LΊAu����23R:g �ZB�N�R�0�V?쨵W�
X��H� ���;�(�s	Գ��ucf���1�^�^km繟�ҵo��d������O�����:��XO@=��������`�z���N0'���A���2�J�}�ˑUk�΅�C6e�뉲�,Kpq�o6Oi7Ps.����=E�RU��;*�eB���K6�]���v��_�_������8�н���.��l�r�u�̇-	���(�#�2�P���L�g���C��M#L�RQ���\����M@�ie��rc�}f{#�a�ǍNXw![���Q�Mާ���}ZIi���	د�v`�����{���4oV
ש�rz`���:L| �A�����v��}�=/���_�1�~�2�^^}Y��+�AK�n�}�e�h}��M�&%� ��4���!�B[K�Ӧρ�`Mc5֝�[�!ە�Y]0����Q?|�*���N�-�;o� �^L׳����2�J �H!�EG�H	�k���,����{�%��hh3�{��\i�c򮘩�2�D,�������-}�;s�2<ȡ3b _cWh#��%�m�z��{|b3`�Y+�A����tƜ�����,������ϼ���fqz
 ��4��r��<9@����������?��~�����?���wYE�opB9� �L��l/0	E�gZ+%����]T�M4������և���%õ����"d��������^�X9
Bو3B�B�����i�Q���$��&�)@�f}�}`	�[�->�1K~������Y�17k��l�{��'���6�?v�M�q�E���L4�*3�����6��Lj~3�{�8�ầw7�t�u�Dm�{W�8g#h���,�*�2xRު3��I�R�e�lڙ:�uCu\+r4��K�'�Q&j��Q4�{^:kZ)��	�D�N��vn�n*zp`W pmB���T�l�s��	'"��oTBEi�S �sQ������-�P �����9F�99n�r3�+h㵖�E�Z��@��{�s�hPG����+T�]�h�tm���>���J�����I�X�����c���AX�S_^1��{ ��e��ׅOUR�Z����}EzkS �AY0lس���(<'v�3��I� V�E-g��1��|�38l�*����J����c�j��?T�>bm��[�c9� 	�!C����A�'{Y�wv]rT�X�԰���g�!��R�/��e �<��kx�J����n�*̤i;�:�l�b�D�5��Y������5e�#�ՋMVq @��%�b�i �K����H���D?�Dv�'��k���+һMߢ� ����I�</�8���UoVu�>_->u���Y�,D3^ϯy�vvť� Z�d�hVs�t�L�@6���5�8R7c�K�v3�:r�7�X*�W?]�~P��3�6: }{~��^��?!��mN��'�Q���X��T�R*�`L&�����kV�zះ]+�0��嫑�~="��>+�Hu=د�Tb�\�@
*���yi�06D�?il��!�ƅ�}ْ�L���5;|�%ؓ5��#��������C)ʉgP�������<	���K��G�H���c�WL"[%�[،��&��̯uB��1�9�uR����_>(�B>��
L03r���?�I�A{��Yߎ�xkZ��_b�$�f�ɛ�H��+�&&z�,,�~\a���/O^���_��oOG���]}<7�� p���A�+  5H��qY.2�}�8��P��y>�|��sSY��D����o��r	��U�_�+��:���*�Z{�1S�$��ulXPlpZP���'��c�������Z4��G.NN�:�ۋ������N�nl֬o��("f�'��^p@;���Ԃ�St{j,��8h߶��g����ohK�	��G�M�e�
��¾��?mQc��'6m�h�>�s��8�Sl)����t#g䃬pl��>.���X��@cc�imxl|�i��9f�%�,�5�x�Bs7�.Ц_��s����,�X��ɋM}E��#F�K�b8��������_1��R��-d�|���~X��
�����Ld�1�:>�_���/ȉH�o|��'5d���c�	��(7՗�1�j���M�l߲s��*,���8�J��|�㵪j��g9+�%�c�^�n��uN: �K����䃓���S]KTOl�` ��S�[ԛn���n3��sǓ��H}��T*�E�ߨsw<�?��ac��O�� �{�}�#�,�  u/yͥuCt��Zľ4G	N-�A@n?�6zI�;� ���.� ǭ�rV�!�ЫDA�!�Vq�?��������l�fL����v��|V �O�Y����-&���Ɨ�x]��!���!�|9�B������<��t�\Ȥ>��� ��
�����,۱!F��+d[��_p�(����Y��[�u>Ւ�>�������Q����nvv�Qp�\p�ҝH�*Ƿ���a�i���$v?~�.��-�VX� T��v� ʪ �-w��xRK�e�+��]�ļ5=�7BP���3Gk��ua^���/0nG1��"�$���&�㷙����e� F��9�( �����4�y�kh��%��Ǝ���4�	T�X��}��+�?Dg]��~�>	І������̂��rQ��z
It�V:^�6�_�}]�� ������g�3�E��^~56/�7{�%�)��&�z�w�n1��	 )��R��0N���{^�1������j�[7f��U`�ّ<�
���x�׈��3��L����8k0ْuf��!��mo>�uṶ�({���[ ��t���aiyN�4���|$hj9e���z*��u�P�7���1��y}����F�e\Ė��h9ga~��Άk�\5�V��G!dc�j�W[A=6�S�����=/�cEJ�n��i�6��������͝{����1R+�(G9�Q��! �����t����v��Oʐ�7$���X���V~�W��\\�_�H���Pނ>S$�������B_�ޡF/����@�.XT��n'���@\O����	��cۨh��椲��o�2'��b��x�*kO�V��Y��Ĵ@-6�П��@�.�d7u)Jp��G�W���ߪ=�����=�2w|٭��x6�'�7�`ӆ���og�h�s�X����\��
�U�4��~�R�9������w0�SN��C�?�p������L�K3o~�䫟�<I���<�l�6��ϻ������AY}5!玓 �	�51�d�l�^�i�U�f�����X�ysKcin�}׌��]�n����9݅2�N83�58��}?���x8�D40j�ad˃2N���f�[�v#}O�-�{xa5�)�G����dB����t��M0�+�=�L:^�8��gB����uAΥ�/F4v���o��N{�6����l��:�%Kw�~L���L����Z"��3^�ԛ��nn��R�.�zJC���l$ԿEstN�򂦸��{ڲ��|k:ض���<㭱�0�@���P�?��ѓͺ{w������EA�f^7�Y��z"-�y��n)�����:��ڮD�{���Be` �)�
�7�� б��fG����-��N�ı3���>|@o���	�R%� n�v|�͔�3��kA���?ܑ(�sK�Ԕ����:��h�����6�}�n��\��*���ިA3�H�s �����KU���)x$��i� Ǔ���R�gXO`��}(��
�!�	Moh�d�T�"�e&K� ��|g�@�}��'04L��-���ۑ��V�E�,e���������G���"�_���G�/�_#@%*W����ȁ�v����D�kl,y���7�k�}.o�v���c��S_��}����N|��z��Nǫ�|t�C||W��ֳ�_����-���M�����o��|��Z���i�،��˗Eӯ�f�*����l������;8 ���ho��f}��i3^p%A�,}Hz(F��㵤s�_	��k�D�UA���+��^}��Z�8h�k���{ɠ�n�o#�4��3	�����/�������!�U���Z���Vt{'�j��}���w�ۭ�K �yC~	���/��}����������$刔�{�l��Ǜ>�@�|���}�|�į��ݶ����{<�놠��&[�oվ�!��o�r��H�/஺�GH���1�z��C ��׸��i������5+�>�Q�a�|�d(�!i�?�s�.�ㄠ�@A�3~ԾN�6<;]��7�m��v�D*5�r�w��׮6w���͚ƒ��{_,�Z�(G9ʏW ���4���������vT[�%�N
Rh���;�����@e ��Հ��M�����=y�P��(ް3�=��C�#��\��>�Z�:^�o�<��:F�]&܋o�t1�I�2x�`��?���)�j'*�?� /+����^�k���6�Bm���9���\�(�C\iM���S�}�i���3r2#��}�3�2�y���ّcO���Yb��mpj����83o����N �AMn^��h</@5��Ӓ�Lӻ��|O �q�Ps�,�2��P���{� �L{qS�&�U��D[ ��I�����9�I�
�"�NSɬx��)��͢ywЗx�pS0f��r���=ӱ2��3O�+�w4ɥ~hF�$ wd�9�X R��
悩:�������DB<��9i���)g�!����Y��S�_�L/�BL�\ງv{F��d#��Q������C5��~����MI=�ad� :�Up8�G�i�\۞?Z�~u��o$K�$���_������0'G t��mA6�hl�yJ���a$��ϰ_7��:l�<�r����W���~!�FC�F��f�ш��9/�:���Bl�<e�I��@"�����=.h]cL3�@�O��N�g��AdG�R4`��X�K	N HN������l� �� \���c�e(c5f;�(�
D���lͦ%�=��و��b�^4kHa��"��-� a�_B@g�3)@��S���/�}��(d�j}r.w{�ӻ���,��!�z��w���S�Y�c�8��p�
��?�Ɏ�� ���Z�į�>	|���U-���8to�ۈ�   ���#K]t*5IY���AjUPU`4�Q?|pŔ�1�ְ�Qy�k�rԿ���{/e�*f"+�n��;����Lu����9���sM ٧=� �? !a�E��ش�7��}  x�XK��8��1^/�Qc[�: Χڟa�#��-|/�d  ��4^�_��=Ԫ���ɶ���6_�@��)�J��,��9�c�1���'��`{q+�Z _��X+ ����1SfݘM�a��:L�CNd��:�?9���JR�4V����V}��dݶ�0���}���pɏ�	���8�v-���i�z$@����K�����55�bB)��1�� �|gmԝ�L�8��$�Ѷ����`���
CPil�]����gU�yu��G7�}U�T��d��1�#�Q�r�d�  �)���bq�w�����������lz���"WVU�Vkȴ��I)�g�W!������L)Su�
��kE��M\�R����5X�f�k0;]��@�H1���b��JQnܞ4�n$+)��Lb�V qq���o�J��2��Y�{U&��n��q-d`� v�ke���1��Ԧ��]˪vls���m��='��1T��?�p�!h�{�=k"���e���2�����.ݍ,Lx�^��UB�97���@-Ԓd�f��
��&?�̃���aSe�! ��NT��x�iv�<��o��pA���@�Mj%�f���������x�?���a@� �V�
X����|G�
����	8��~%QT2�b%t�p`���.+��lN�d�&sf|ƙ/�����K�e�W|�E�Х���$���g���3�Ԛ,�3z�ɑq��3�zg�T��BS�'8�u.�䜧����ľ'�ؾrܡ} C�ծd��H�U=8�5ȂXG��yP�߄rsʖ�;��2^xȠ��4	V ��PCy�k� h�X��<w�~��CpzA1�1���
��܉g�\ ��P�?�7���s�\C�?���u�j%������̟O9�H匙22�Lp�<j��f��M&��.�W46 `���/�	��MI� q��Daܬ��˺/M�L��n�=>��S��������'[��+�C3��:�i��� ��Cۺ*B�O4�T���^I3a�4����@�A�wь�+)�5>i�^S��PQళz���	�
���f�lC  gH'S9a%(d391�YY*�6��@��IЋ�ht5��qԯo8[��D ?(�z��{�ѹ�Z��p������X3[ʾ!^�t_a�`�|��xc��6k���m�lo��j��&�����\�x� $���Q}WSI>����wjS9g7�t}NAH gNϥY3�*-'�D T�c�w���{�-�YAe���~p��xe�z-w��� ���[Xs��;PA��s�x�VO�?���$�V8�i�H���� �����7Zwn���Rb��kE����o�_�@�b��_�v�@  ���:�)��{?��������Z�{w� �'f��w��XC0�0�0��9�(MEelx�P`�����v(�Bw(h���L
)o���1}��s���H��_`wf[�B�Gېdܷ@�!j%jj����d�!�_��Q�/@nO�M�F~�3^��}�C�$1~���/@4��Wf�v�d���ʄo��h�"��RI�tY�fԬ5S�q�7�����������������W�{+M7��(G9�Q9��������?x}�M��Lu�hw[;ͣQ�����g����ﱜ�"��)��.(���@�"�"R��>�����.^�_+A���b#kYL��MF��l.����>k-658��*��#�O����݌�v���Qcہ���v��ԓ�����:���¿�9~�f����������)۸~ �������L5�-�sl�Q2V�fxA����6@��:�w�H�'�TI6�B����GMDP�՞�S�!T'�c�Lr�S�L"�T���	5I��p�M0�eߕ��y�=o�f���{8F��Ux����2��:NHh�J'�C���]=�8���'� �*�U2�=�#1������$8��y�:Eh#�D���NP��Ӹ��p&�Μ_;rx��&'�~��Y�&��+��v`� <撠5?9Eɉ� '���N���
�&��ƿ\G���+Ե(Հl��,P�fl���K�o�A�p�ӟh�(j[<$�"���{�\� �7䀧z�wL��X�Ϟ��k�qV62TK��ǅ� 
�r+Ϡ�[�����K�TmC��d��JʂE#3
A_�>-�l'�Y��M ��鱥:� ?�npX��!��[�Z�JW'߇Lw�#�pB#s@�U u/�B5IY[��r�93-�m$�¾�\{����|b[�A�����E6-2�f��=7���0����E���d%���\[z��~���N��'�a��u�mﯫnM[�agF��5���ڼ�3е���=(|��ڋ�x�&V ���m�9�Q A�P�M��H��u3_2�k��:��ظ'��e BE�6���o�x	R��
d��. �J�T����\�/�'4��8���No�#l]��g!V�;�f��Y6����{v9��e.x����σ>�����{�ğ�dJ���	���:�X�EN`\��� 2�ZpN�t�(+:�<N$Z��P�}`�7�����*sbS��2  K i ߑK0#�S	���cfn��z�� �({g}v���=��r��+�c L*�w����J��x��b<&4c�q� ��EKe � �};>u᝛dO�O���~�Y�K�nQvi��kI㗲�-�	�I$lP_̣	��\�Z�������x� ���a����c�6�a�؇�]I~���(m� ��r���d:m�e��>�Uɬ��K��tط,�o��R�������nw�N����ö�%���u�?���e���m6�6��'�x$�/�4q��f�����@%1"9Oc:����k��8uh�ϥ}��q����<B�P�$�l��3K��r��N�{�����z�C�틿��/�.���v�k��k'ggg3� ���(G�} ����������kW�/�����]e$9X%�xIir�����"�D����f�+�KP�!η���+�Z�BV�-ZY����j�7V�2��n����0p��Y���ְ��&n*���yƾ��2���=&�N�� ���q����1�I�s���a؆�[鍥۞���=E��(o<�;����@��~Al�u#�X��3ǎ3�'GmvL�X�w�.k�e�m5�	N!sv�ϥ�:�'�]�`j��xP����3��.�J�
�n�&?�f���g@ Gl��w3�s��Xqvg3r���J6޽�?x�I Y9O�Di�>--���D=ŷ�.(X��!�ȬX�m�I���>@��35Q6 4�T�A鉋5�)�����H��@�2 L��ݖ�Q@cv��ly�JF�+����<9�8����DN��h��r4�L^wK[���ʧ������<6���3f.�R�_8Ig��)ARG��WL,�Id��f�f����Ï�W��K� ^w�����q1Ul�[�W���{����`��9ٟ\����
��8�\��n���u����HlT���]Ha�"�8�����sr�d�8���S��+��RbgO�ĩŜ>��}�K�R���ﾙ��>%Z� I;�g��-���R�~a/��fu�y��a�<����@yX9���#s�6�9�E�	�YYܛ=�/�9Ѕ�� .��II(�1����.�~b��m?� 0�c<�c��a��h̟9�,5m@�(����>3�%�Ǔ����@3t�5�9p-���>���W]#
�R�����Y�xc��� �2s�ؒȨ��� ���-�<Ô���>�.c"̢�y���X�pb�:��}x��O��ʿN�sj�ަz�v~�	U��S죚}�\�{x����"�G��a|R���H��r���oa�3a.Q���:�n��Z�@���w�x����e�A]
��1c��1Ʈ^�����J1e�z����i�I�����=�:D�]2s���� ����� ��4g]΀�bh���K��=�qHJ�����K�p�%�^ ��_�L��:����c��%���'�-,k�FOs�m��\$�S]��UǦ>�6�����N}�F��-hB��}�o1�Ags,��>]�[>�$��k�����NOc��	�����cI�a����1�����}�>�b��j���^�*x��x�XW6�z���-3_ܙ�˩��[���/~��~, 7ͱsk�m�(G(�` 0��{?��I���kWY��A�_	򫝍�R:^�)�
�䕱mE��jcU�H���(vE�v As5��_,�+'�Ũ��m�B���_NK�q@����GR�F��Σ��|�����O�md_�L�G��|{�W�_�&��`���F/��v��A��1C��M�'3P�V8ۆ��)�Dٶ�����e��P����S']Y�V&�q��:'w`�h6D-���)'���@j���������Yi.�� �'U���� /Nb ��x����-ׇGv�f�k�{q,0&��,��Kv����t��9�j&���x�:��x�3��B����4������s �Jzw7����0gW9���(�+@�zOA�ut����x���F��)$����e#�ęL+�@�����>c��d�_���������|B�
��C�dͦ�y����ѱ!�����o����0��9Aɒ*�i�z��Ϧu�t;q����;kRMYH�2*3� @�%�^fq]��.Fٮ>O	�Vm�uC�WL�[�x�1['�Ut�-��xaN/���)(xr^��_3?v��V8��<c���@����R:
��<L�./kd�>����Z>5��Z��B��G��~B��/^�PTS�2��(b�����a `��������a�^���1�8�fV���UY�K����?:, 0 �EcoV��}=�I�����Z�a�.��` �Q�}@�*"z�I`rr��NA�b̠��`��(�F`�g���M%G�Q:�jn�3@#dgCw{ u˛��Ϧ�ИT�����1>���ڪ��Ƴk
6͈)��6��uE�:�riRs9	2�%���g�q�_��}��t��\�`�J�=��n4��&�,8	@*a1�a��$��T�i;���S�%�� �>g6+��$�u�����,����S���*�V}ϱ�g��_<A��cYL$1#&%Ŕ������e	P@�@�J���@�J>5��G#�g�`��q�ߎ�y&9���W�c������蠨���z�D�<�|��j��p=?a�{��V �
��w6Ƣb���	ڂl�%���'Ir���4�i�%|��3�0�e�M��iB��`kɪ�� �{+��˳�O���
�c��(G9�:9 ��_U�z�b��y?]T�*Ш�2�`�s���Z>]��
�.Z�!�l��%20`@��,�)W�̧��nȤ4��o�*a����Lri�f�'� v��m�e��Y��oYx`��`R����0�ƃQh��R7��G�}�����k�5-��\1�����g���R�p!�C�c�̇,��,�U��_�{���� �Sdk�c��Z���kC�q)��C���i�n�*	�k�;}RC2c4�W��(����<D�<�uلR�]��꼣M�P�¦�Uienf�A羃3�X�K3r|���k0��Jt ��%j����Gʃ�h9�Ϫ�T@��~�Z�(#���g���W&����ꬁCN����bN�~�99uC�WE��z��{%��%���^88#Y%�:�}P�E��\�,�VT3�RgL��vb=2(`��R����nA�]�����IW�V���Efش��o���ke���V��=�8���~��K�5�3b��cZe�a�ݚam���+�����ⳤ�?{��+͒���̬���}�t�����16�Z�0c�=�#[�X6�H�~�o���@~3�����4/ !? ٌ0 �Hfl���i�9�m_kWeF����U;�^{�Ωo�%/���+V��o��}��&r�cɛ�/Ƿ���幂S٫.[W�2��W�pQO�3;$:|n��5+�L��ĬF8^�pVH�z�����6�<�6B�t���|��G� -��3�ǆ��}l+�R��|����97���������-�ba��^ʍ�&)��G6���>�LF&��o� ����h���?���5֩�}k�}ɔE�l��xP�y �i�,�Í!P��MN��J�V)�Z��l�e]{�1��"	傂������x`��i�¬%^����S
q$>}���O�)��h�S����X(�A �����F�=�^RU��ܰ�kK璾��P[� ܻ$�?�>�W�4��EƤ�YR�r����G�R��#��(���M��h�|ԓ:g��ID|�T\^Gtf����*�7Z�I2���ߗ�9wu[Ú��KLu� ��3�^e��̓XR���*��T�N�S>מn���-u�r����~$aR��K��!�O����lQ�����/����7bG�4X"�=S����}K��
��w�o}�/tOpQ�F�a�@����>]���)]�������hӹ�Q�e�;.n������p��k1��r*�G&e����b!�miF�ew&m3�~�Q�7�@~���}?���ݟ���xd�A^�� @j��~�w?�˿�������r3�?�OM��2�A�'��E�JV��E�ZNM5I5�p����iV�r6Ai�Q�8����l�IL�2�j+P��4Ze��$SA���d�.O�Np�3��$�����E3�_O��>��t�t���3BF��"?,JcB{�]�A7��Z�z�=Jj��Nm�5���ҵ���T���י.������:�qW�8]���t;D�����?�x��!$YYc���G�e�p�^�V��Qq�!a!#��ڄpp!2E��D�?�J��y?���<�݇)J��dך��k	?�p"��S��0̚P#[0e :1��(D��4���:�h���Ju�hT�DTi:�d_���HV�]ȋ�5|��/��?[���$���a��
�MQ��(9�7v��`D�S�=�/}��j5]�T�/�hߑU�ʞō���S����[�t���N&
�2�G�����Y2��x)��1L�s*i]�A^����Ԓ�j�N�g�t��1�0�גXӹr�?9*mE$ש����_�FKeLz����ɫ�.q�D5�K"��S) ��2�׳���7��`Z��,�g�G�^��m|�>�Ø���ݾ/�IPxq���QF��C�;qy{�LKcM3t%�oL��E�n_Yq�mCT����M���7�m�  �C�ڟ듇7_��ғ��d,Y��R�
U��h�iv ���CH ��]�Џ�>,e>��ON|2�Y��ر]�Se:0K�*yi��=7���x�� ��]@��mi>�-|~�Q����|s+��`{�|��|�'�G\����l�m��N���X���E냂��ݩx�b3ִ|_�����w>�Rq/p'ҠU�������d��p�_�����_���)7汪�' �2�3�� _������?�}����_�o�?)�+k-�miH� Z`�F!���u��߭�����
�������W�E����J2��RP]�+l1���dZ?�>@(@�ٌ�!L�y@\l�W�fdr�L0�f�i+�SAs�u��A:�y��7�	i~�tznM��]�(h�#����ֽi��m���3��`�q��K8vY��Evզ��O�צx��9}���n�ډϝ{��&#���?��M�ϵ�xa�Ġs��&�uI���W.��fɅ�Z�Yy\L��ƶ��N;�Үbz��u��5�ɱf�Ϗo����5 g�cEN���3��O���vg*!Z�*��_x,%9X���&D��6+�̀�f���X��k2���!�I{�����Z�xu�8#�9�ұ��Ǳ˿���V,��L�e����c��Ue#l��d7U�M�A�9V���������)H��/����s ������dig˙?�����ښ+����s��?ٗRWb�i��3������c��X�TOo�Y����+�^�3k%�6�\1D{�E0�}��]�[��M@�D`SZ����%��#%B��$5������j���Aj�s���~h���B��F��,��=O(�c5;��F�����zRR�IJv$`�5f�A2 ��x���db4�ܦoH�F����/�r��d(�˳;G/�{��{�x�\�^4��3.��C�u>��¢6lYQ��O��|����j��eGB�'-à������8��QO?7^�ʦ�LW3t��4����!���t���{S�In>�A���X�c�M�� {�+�����=�(	^�#�1ȩ�JB~='y[@|-���[f���rp�3�Gx=�\���!L�j�Z��h���JF˂/`2�#Zr�6���}9���G'O
������1�hy� P�$��]��w����ۧ/O/���??9���2� �,�� �	*��,��b����?�������oW���a�����9���#ѣRǔ�1�L�8�g���ӶJ}��XOI�' z��."�Ԯo F4g�p�m�3HY
e�nGii���t�����D����zC�7�4�L��t���\��px�	)�#]`���&3.�ٻ�x�ڦ_��,tv~�ڞ��8��㯟:�O~�N�+QVp
�$rZL12]{�.Z��q#�̊ݶUQ���A���0b��t�apμ��i�|A����H�b���+(F�c��'F���5�[ջ�7 Eaa<�p~]	�8�ڌ9����-���!cD��J	Y$n���:�q��`�������V�/�0�����n*�ɻ�����kV<;H�9�C��g��un���z��5�l�e0m)�0r�^�c���9�lq\4	,!�x$)��S;w�GQ�֬p��ۜm�����;�us�Z�4�[ ���Cb��+����}l%�E�*��QVLJ��8CXVHF	=f����$��]������m4���v#��([�x�儔(褴�v��}�E��2V0�{���˾m���6�j�%v�k�׃�*1��I�]NX�M����iz��������6�]��4�e b�g?O\P��|r\mǜC�Z�o]:1�8%I ^j �Q ��'%Upp��~�)C��+����qJ���ZYf���٨������yq�������@ d�A��>2 ��z:����(����,�\>�2E� W�r�����LP��)hy��rI U������X5+$�'�hÊ��\������2�m�����5* (�\&
Q��;����kr�b��ʼ@Q��Yʶ��۠z����4�O�7�vN@�����#i qn�4cC�>�Y~�9����niQ
��ҁ�� ��j��g{1��Й� +�:~���sE�Y�"hm�)������tϏ�yǘo�f�;K��q*O���Z��fTO�$\G�/;�8�g1�P�3�G���{�1�w%�\#e�Z����g�����]0>͘Xp��l�Y���]��_3�+�^���-��Y2��ػ��������饲@77����;[?l��͊�/�j�����#�;��*ۚ���NL^*u�)kc����1f+��ߺZ�d�7�{��~��Z6`��_�B���p���/;����|�T6�n:N�DM�ԩ���!Yc�9�<����>�3~7�/l�)9Eɬ�v[ �mtٞ��k,#5�3�+�u�m�*ڝ���������.?��G~F�}��Әbp����_Z�}~}D�Lc�,�%��Ў��Mg艪�g2�����+Io���������܄�j�\�n��d��>O��-�`�J WĈ�cXTln�A�TLb�b)�\�/t��^6��fM���);!�*𙒬4���]��>������H?��EM�������6۸��� |X������i �Wrff�S|dW
/�G���~Ĺ]��6D��:"baea�<�{h� �\	�d4@�I4��%�:x��c�i�pb ̺�F��|Vq�$�t����I�DC�P�3P �p��>���u
'�Ng����[����~
�?� ���� �y6�����q���}�pU�H�W`X��a1�ʖ���>}2�$�1�k����m �yq�l|NOxM����Q��X����1��<x�t�F�2Y��t��c�	��2x&8L���=�L��������,�&C�@�~���7"M�y����i|��.��� ��W�u�2�i��E��{�>���[��]��c9�5g��uM��n�Lh	e������o�8M�/�Ԧ�:Jщ)�?}�D � P�|���tQ/�G#K���Y'��$�������`��Ō"���Q;(U��=�%�}�����_N��Ð�g>t,��R^`�I:���5Ȫ����t�X&K��-���6���r8��q���ѮK�����$��]l�תw@]B:^ŷ��F���/�Zk�d�2� ��$
���흧�s���+dK���$��$�-��Fĺ�Š�im���j���Ѧ�(�}��.�N�PN�5�5�(�ޝ��@�
�v_���!`�k���h���m�ZT�iF?q���h���R���*ڇ�2J�	��Wv��\E���>cY6v�ג�,�"�@ܯ��@��O�Dw&f&��*r����9|���+U�dГYY�(I!.M����Z*���Ul<���(�!TK�'NXkdW joR�@���YB��F`�(��^��R
�EQ��J7�w��P\�ԛ[���Ad�ge/��(F�n��7�׿��ǫ�4Ӭ�U��@��&�K3����8�a��>%]ӥ�E�Y�4"�!~/T6J�o3R�.E� (c -
eM	Iր�1Ш	24i�M&��:!��</�T�1As���c�nO��yb[�ն0x�˹�l�ȶD !K��J��JR4P�*�,��ي����g|�������E��G0�D�����>~� � P�侢Ȝ�NQ�1���;��_W9�^���+K��cD��2
`�Er�IDO*�	`���:p��8�L�3.+`(r�� �W���l�cQ7ȱ� ������)��D�{i���w`�/Ψ�T�^"��]1/:�5Ѧd�=��o�A�4[��.�f%�eA�]��Ih;�����&����g���^ܿ�_�r�<��:�{��� Ws��&D�O�����R �k0/y�
��e5�3 ���V/���?���D�?&d�������%
�m�6� /ER :*�y�?�~~��x	��� ��� K|v��J3���{[���$���c!z?I�}�%bY稷#��p1����\l�Wá5��n�s9�A���L>L#�ҽ��?����A#�c��p��շF�Az�g��d�A6�� <������_�������?}�M/0y	���t���%��Mg:Y��5"ћ����N <�ئ�A�G���,f �e|U��{�Z181d���^S�C�`L`�@�Zq:i�?=?�$E��81�GYc#�}��DH@+j�M	��xڟ�"�bI�6Y"�&��+l+4�][t�t� �,Q�L���4`�I�\H�X����_�~_�C�4�y�W�}��&�Ե�ǒǟ�FA`~���>��§o���)}�>V����M
��ep~i��M���]p�O6��}�_�(�	 Ӊ���{���"Y3��L��;�3$dD,�9+�eg�y�V���՝�!��u��n噇i�]����˼�f�7���b�>6YD��ʱ��|߮r��S�1^�'�۲Kv�"�]K˚Z��]���%�̸��z��Z�6�N������f��)��|�*������H�-�x/�����arW������H~�������x��`��L�|��鞏�� �tl��R/
����qL��f�-��܋��C��*����0s����37�D0>�ɭ?�J�I�4/�yX��o�97+}M��=�]y�ȳ���ۺy�6���nm���^��;E=���<ּv�$���� �r��铀Ii�0�e�������&�?�%�#~qā(������PF9��>a�k��(�@ �c;���*��
���� �R3������������������l6����R V� �2ˮ3 �J˦����~��?S��猪�����F� c�I �N� h`d����iX���J�Q����if��p6�F�i�&##�i�������´�Z�m��u"�Bᦦ�&��Y�+�'�<I�,�E�Q����.�=����:i��F��	?�dih��MiǶ�A�j��8K��8�K������/�~��X��������
�����`�U�e�mu�:�ܟ=U�p[R���)ܾ����&�0��ǿ�/�g"�1������7��:��ˌ"s�f%0����O�2	����>�lZuF� �ᮄ�n�)������sYɅ����lr����˖(�cѵ������������mx\2��=�ֆ¦���}�;�߶��[.�+� �Nߖ��0hz����������I�@�h\�1j[I �/����l���~!9�M�q��$
8	Z�rH:f�<���lcR�����di�[N���k��5��Gr�ya��/�$ҧ�ƀV�ҹ���MÆ�SV��yV���)�͘�_�3�����o9T�3�4Q�p.�d�!(���$ >YrM>4:�� ��>!���	s��m�^���0�}b�Z���#JI� I��I�%.���aW̢jL�����]����w���w~��/~�����d�A�>J �w7�����^L]xW��2
_&�S%�F��	��3@��|���c��s�M���mH�kɀ=���F���1�u⋕��;�m�	@�<Ovq�ldB�|%���N����9-�PSR�'ޔ Е�-<A´��]�QM��*o�O0��|<�n�����$�Z�-`��f4�M�rN%��^MǶ(��%�n�׈j�5.>����Θ� ����"�o%����nJ��p���h�
�1����E����+��uVQ�`�:�ίs�>a�O7
"�&�{�5@�<x>$�Ŭ޶����c_W�q*2�1 ��w�5��� �J���>�
d�Ad��M��w��S_�3XA�z��{�
dMG4��^/N�^�pU��'o�5����آr p_�9����ž�eL@�p�?�����P��^K���h��D�?��%G���;X���^��\������^@�Tv�0[��K�m/{�xT�@~(���' ��v�����S��i��p#8P���=y>�嚡Ym�T���$1$�'��1��RgD<�b<�)����א�S|K%�] /,��ϒ�Z��LD%m2�}�a�#��:Sf�j2�֝����������NOO�2 �2�R��G��;&?���'S/���ްp�2d� �$��In�9Ѱ��	r������"��	����Ag�+��	�ϲ< k�fLH��׉�ۡ�҂��4��s��m�P[�	2�5��Nj�9������m�^��iOG�E$G4����<.Mbޅ���@f��۲t��c /�',$*�2��Y�[�we|.j����0�8�2m`>�{\X���%h
l6F�W\�B��F��%��Jf��j����`п�䐺`ܫ�������o�O���O������wF{��;38���#x����GB@Qp]N�>l_�8;Ϡ|S��\�+( F�p*��8��sN<�nOf�鲄�'9乫_����z8b���_�����ض�����iV����\H��F-�*����ί�������{��n6+}��p/�GzJ�[��Kzλ�]'_�Pw�y����s��u�o&������e��<��n��n�o4�i��?9���u����W�w��^�G��Cr �I���A�aJY�<�S���m,/�:(�d?Hv9Y�������]�lx�Cp����UL�[Xz���-�>�ܺ\�}�Khc�,y��V/���NRHl��}��՟�����]W�x]�M�d{�����6�ߝ`,����ÿ8!�?|+ݿFʻ��CK>+8!����uǑm�	Q���%���&�	�7��2$8���Kii�2�����Ӛ��Z�ڝ�$�v�{-I-A��o�S��쩜���T��E��`	nk:2� �4d ���gf�z���O��ɬ^�����x�I$���aL�����3H��Q����F�8+cNF�;���@�B�l-��&֠qIľ�IF�ͨ�@����ۑ��]	'��'�LS��q�4�.D�ܛ��URo3$��Y�l����#a���)i�},e�i�-u���LrO��{��7ɷ�	��4����c�0�^���H](��D�o3��1J ;��Wk�64��:7ܰͭ���L�=�ߔ�#	 ���ޜ۽��l�3& ����|9�2 㓌�{��BP_d�J�^d�	 ����0�8��ACK���yx������>~3��IN����Řu����+/�)0���:ck��%+��"�2Ȗ�s�E�ӵ�K�Rބ�Q��f]��!l�K�`��h�'�sg{�����x)��s�/\�W�]g9�I���6�
`O��,e �h��Y�}o�Ģ�H��/��|�P�i���â�5ߟ�czXP�l�3�3�&��k��v ��c�d-g���e
N��p.�Q��۲L#���X�A����x<� ��&���}���d�v )��+�k�s:G�@f�r�I�a��6N�0��;%'Ի�
���p�r2�W�̟�����}������ �2� �d� T@�O}�{��ֿ����/~�/}���=VW'�Rc�-b��M"��[	6��g���01�
�J���� ����0;@� u �� �Zo&.:5C@�u��0a�ŉ�����%�ͤ< w�0� �������8����v���9�ԴI��<EܦY�#�������D�����p�O\�L�I���x�!V��A��%Ȣkj/l�&�Zc�E2�k��Q�z����Wۼ��IZ�(CՀ�3Us�i7�KN��aJ)������g��ig\~Q���
��2��K��7b @������~��ʩ#Gf����҅�e	ƧOL"87prn���3	�;����2� �T�ؐ��D�5�u�d�E�����#Z6I�^���o ��Ї`���F��D
�*0��0"�	�=��3�aRFܖ֔U�Q���W��m $��$��z�H�>O���.��Wv�^����#����`K�4o��� ��[��4c��4 ��0�m�^�7���wĝ�r� >� �@;�+M�	����?��6��8���s���S���6�zI��Ї���6�jp��a{�3�����}�T�+�u?\��T����~�o�<�`g�N�e�2� �4e� d �\����=����O�����������˴3�JՃ>l
��m��:k ٢���P]�Z��$S�_�X!����|��.��P�J9��b�)c�[�,�pnauI=e��u1w���/���A@s���1�9�~0��$`�>o��|��3�\�Еda��]d�5�K������v��mq�6�}a.Ӄ�y���0��l�%��n������e���e��%a��.�B�h!�W���l��#2ԑXVs:���
n�����X��m��
*���Z�����\���p�� `~#��39��esY�:9˩T��w>U�xW��}�i>��Q�<�!9���7�9���Jt$�;�B\z��#6p ��0��$�mҔ��Bo*�.!�z^��x��s�V�l��g�f����X��Y����ߍ�/��,���k�q��}ӵ�K��Ud{���9_<�������t��}��:|�{�����:�~�1��K��=�f�C�7�\�'�XG_L����� ���Em˃?�� X" ���&O�f�w�� �
�� 7f����Rf ���	��ҕ �[�Y�������+~E��ɫw�����҃��®h^|�ӛ�W9�֥5qd�:�����Ȳ�ل�hZj�����ͫ%Gڢ��`)�xLH���} ��ɾܻ�~}h����zK	%j�,����� \2:�B�2 @d=�+��02��lϔQ�1�{-Q�Fg� I���O��=Iil��\�+�ף}m�q]k)��1��f��Rɶ�l�`�5L�>�\f�Ǒ�w��� x���Ad�� ~:�>�"��������_�����T�Ui\�3���t����� c4��6V�N��@p!]�%P9�}�i����nk�<9}f�(�Yp�Y�= EkӰ.Z �5U�`/M���M>	��&$!L��h�!=�Q�do{V|�F����yyER�Y�H����>�q��'�BX�	�E�o
)�`�W(:�|�W�t\�������񰮐},.:Ѧa_R��O�3L�9g;��-(�gF����@��:��С�8D������/��0���	��aF���A�]��� 	a�P���p���x>n�!g�5B{�~�Ay�"�w�$i�A�Wx�<-���pF>%��҇AY.���đ��} !#�z�C�1p��	3�Q9 ���o��;�`�GW�Z�sY�bĠ?J `V]���`��n�����!����K�v�d���(ޛ�L��!n�l�"撮��)
9�@nH�`��
D��|.�81��`�i�q@�3�L�s4>\�Q�_~���M���[�6g|�+qR� b;F����1�o���6y3e���
���<;����?��>�E�����iòt�AyF�A ���.���O��ڳC%)i��xL:c�Il�$�<��e���\k�����;��J��~��m��z0q4�[���vr�~�����թ,4Z��g�х��jRS�:2�e<��k�ٔކ�A'�fք����[�@�~�ǋSv�KSݤ�i�n �vLO��i�����k���l��cJ���������
�9%H!��It}	7����)e x��(%�u��5��?�,(����\b4���y�JO�K�n:%AN��N��7���D�pS� �`Q�Ϙx��Hx�J��d���.?  S`.rș��M��m��wOR䵋i�}]O�q\���:<�,�X+��F��>�^�Z���ז���ЁA�](�N��^"�O�8�U���V��������&I�7���%:�\_�?�d��ś�I ����'�>��	 �x����lG���J��A�/�kv/,�ix����&�K����)(��fo���læ�E4O����8�	`o+q��@E_��T.8vT�^1!�!�)�Fy!�u�d n��� @�i�69l�Z�,���]~m
��󁖞Y
�p�f��m�#�{�� ���՛��~����:�-|1���d�Az�^ y�g�����k�쇟~2z�� ��LS�$����K�a}��>NQ9�bmN\�s��$ �qB+<��1��I8 ��4��}J�/��4�A2)�o�}&@��+��=2�P�A&"�'Lw�v�
������I[��W��6�������h ���=V��Ӟ eP+b�����Z��U�}�%����"�(�>�'�������-j���ޫ��P���g�(O�����5����:a6�0�+)��7O���'zO��K7w�q���s���_��ͷǔ	`t�1��s*N��s������	���eWo
"`	����n��%I ����{9�c��PF�<�:`�iV������u���ا�y���� +��c�=薝�Kj���|Q�l�ƾ`�`����4��	��W&����7|�Q̂�[�M�e������"�!^Z��>:���-o�Q$��
q+=�?O~���Y�<e	�y�!2�^SP6�e��a�V�����ne����s��ؓ�������c����|��~�,�����������̕�䠡�z�D��® -�b�k�dF@����C�[��k�f3jBp����#��}ڷ��}��@��Ri%C'�f���� ��9$\Z@��ؑ��2���6�z~�c|'�'�T�Y�M�}�%����j�?�1�����?��ǳI5�w�=x�b�2� �,�� ��$EQ������|�w~��}wz5:{�;k\���*>��L�� R����:.Q5Kj`�MR��b� �,�� �r���Ӛ�heRh�%i�LZ����.m�ʟ��$�l��##|�$��d~1K&�fj�t�i�c �&�D��U��^�F(�����d̉�8�]��[��a�:����q���� /J���',+&L���X���n?N���)�|���-F�W�.oE�tʝp�� �=��/Fpz�׿�᮵;}k�+nf	����igW9\��zOE��Svܥ������6�ݔ0~������Y�ؓ�P�s��d�=��b����t�AV���ն�����,>���v;|�u�I���{��xrj�%ʈ�<b�����'7_�s9��[\;<����7��u���8�����5�
ò����>G�_|^�35�}��|6�3�X��/�'���x~���<Z���iG�G��j ���V�%(f��E�ْ���FхP `چ���k��-^ޛ����	���]8�	�I��)a��f�N�Y���]��'u�F,�p )5P��̜���7�_�[�v����\����x<΁æ:r�2� ���#�}Wޟ������������*�0Ƴ�� ����C����i�8JT���7��EFkݔ��0�hkcC�g� \�M
[�B��^,|c��l#N��Uj���$W�SZI��Rd��5�S�7J'�8QtI��N�SC�5���D��(1�&>�Z ̪��pP�p�,�-�h$ΠCۼ�,�Vik�[V>�:���;���w�Ų���oŶ�J����}�Q����)L�f0},��fz������3�����/Fp!�5��Ɛ���]��VM��}��8�3}��z̨�g�aB"�3��}3�T�Xr`|���e���I'#Ә2ht�1����iR�W� /Z^��=�IvO�Ŝ}��%e����C��G H���{�:1�%���~1�QK�*�t��D���_�
�E`V0'n#��X.�(��DR �*�$�>r`���Gb���#�����`Upo>��x�X۵LL|����l�1]�31~�Ñ��!ۺ�>>�u�5�&>�+&ɴ�|ۈƇ\F�)�ll���@G���rT�>��^�|̔ڤ�s��F2�"MV������L
�����@?rFe�`2z=
�$��x<%p4�i�g�s�O�)�eH�� ��)h�H �Zoa��������姳�������,O���Ѫ �2�B�5�4�/���Ǜ����ʱ���1E��Yކ��r�oc�y���!ʞ2�[�����E-�)f������ �I�+������k�!]���x_��ڑ������B O2r�tzn��^����S��*����`���3h��	�S���Hpp�y�F� �����u'��1-�}�� �~���m[ș��C�Բ���6���3r��oA�����v��dC�?���������n����ӌR�# ?�G� �����or������uq�S��h$�y� �O��y���8t�!����a:Ap���[&P)����X.�fS��yv>��Q��YY��?3)E�>2'�����s<+���\�O�٪ݾ�+���Ԯ��+�)��9��%�k����]j����~��.ْ|F��T��{?��9ײy��L1���C��-�g�b�����vz"����	���z�Q� 3�!����� �L x<���P����B��2�U�t|��� f3���v�;�U�h��q���°4M_��x�������{�~���N�ƟNIt��	� }%\�&����� ��99�j�4�7f�χ�1�`'��4�~�㐃�u�J�/ӣ��	I�O��3(������idZ��	�@� t��7L��m�bl+�?M����x.�i��^C�L,;MmN7����M�^K&h?*�b�����,�x��T��=]���y�����_}��	`�#�2� �,��d ��&����y��ϡrH�6�4��Dyp�L�y��<�,��E9��T�2PB�*1Bi�H��9�~G��|O�D��|�y���cv ���|��@� �c
���L����u�~)sM��::���y��K�	(LD��z"Cp�\��4W����_:����dB�P#�e�Y�|z^zk~����[�
�ۼ]ـV�@3���DK�5�B	N��C��%񫔼〢�1���O�D �ș�0G@��ϯs����_#*pvU���r��
Y���Ղ���/���]��>�UN�'un?�(��䱤�Jh� 0�ۊ�SS8����͌ �ۋ��cKǶ����b���dEg2[�d����ǿ�_�(1���\_l�۬����y�D���e�v����������׾�r[}r����=�a_y��������t�խ���1�߇�o{/�KHϰF/,��p�9�nE7vq}�rW�����Pr�Y1j�V<Y���; �ؠkZ����iP_��%r��r ��#P��A�!t�٢r 3��3p�c��8��c�s�i�B���dR���uE��kۆx�0N���Y��^RZ�_p<O�!��~}��y�}�6��#����tX�����mݬu��e�̶�䃠��f��m�{,� � ��^@�#��^��aF[cC�=(�c�qF;�=��Z�K�#A�
$q��8	v�H�����W ]�4��Q�%��6|�� ��bIh`������J��0K��f:uӋ�Ώ.�?���z�,�m��"d�A^��  ����?�3��0�K�Mf�.f�&eX�r2���BI��cD=+t^�3��I�eZ���D&<R��:��e4QŔ5NR��	����)�����N�k&�I.�Ӿ��4�е����P��$| �~K�v/�`��^�+:!~V�@k~���E5�@�nB�H��ȲS���7�kv�L��&%��u�q��w���^����f�b��6�9H���V}���|�U�ՒV�,�f��*��� p�	S�W���}��uL����_�(��e�%�*����mI��:�-���3v�]�)���n?���`?�T�J����6��J"/ܾ���y���1�@���ĸ]�������2v�k�e��싅|��`hu}?�j�Cym�T��[8O��L����a.1B���_���d=�� ;�9�ƟUD	,
��v�a��ATV��N�u�.t�"�V�#��+v�7��d��1�@� ��Q���$ �<�����3�v���o��5��ri4-	������5�nffs%goS2�Fmܕ�\t������s�AV�}��ZrLd���>�y��� ��q<l��IP!�� ɚiL3 ��`x�y�p)�G s�?�1���S��m4%�22�Fұ(�?���W�%����F�B�\ g�,E옼��+t2*�A�-v�#N�w�Y�m��L|LŖ��@����S�<����T�����Err����AY,�  �����+�߾y�O?��`kU��@j���@1^Yfё�%o'Ǔ�I�#�>L��^�d,/Y���ni�{v2�l>Q�ay����&�����7���@^P6;q�k6M�r�T�N��l@����׹	b}�8Y�E�@��3(_��e���q ����洎N��Cs�N� �(4a?���������8�gg�����������x�L�{j�H�ZQ[�)� JL���?���0�O�L���}*)�;}?�*t�'�/r����\�����u�W9��Δ��"S��#o�`pp~U���
�?U0��YNk#y�����X�� K<ܔ����
XN��̲S/�9�&��1�a���ZX$=/�`��nD*�z-�p����������:��>ܿ(��Vxw���9�l �Գ[�8� �hE�{E�����I�*N]��6��>�k��8�ҲV�s�i��W���9i���_�� (�5�+�#0�~�ف(* �}��T��ɡ#�0�s� �,�� �����(@U���{�v����z�ᶴ�������y.Y�*`��k=�[C��3S��k���p�Unɖ�8g�.�?���f���]�}����Hrrv!��߈P�-�W�/���ϟkɾ���ng��>���O�������R���M���/_p�O�8�hL\w��:���`
����6(�Yq��df�>ڛ��k b�]#�cl�/2�GAx,���?jVI��19 U0�&CĆd\6mm�P<E�H_]�	I�s�����n��\��?�o�Jyy�դ>���� �2H�� @��g�\M��?�o��?������>|���z��tf���Qa��%8/��U�ߘZ%F�'��K/5a,�#
���I&���%���)�����N�8T����5zN��$@�p-���)f��~k�\j3�_A����olG$>��Dr�\�4tO�=^k�4ϵL|@Ϥ�: Me�=w�]/h��/6p����ͫ�ѱ�\P,#s�o�CL�f��*�$�$#Tpx�{rh�A�����z����#G����c	��%9��(�>��N�r8�b �.�0���HtPG�̢�(F1���>#'_a��<���#x��(����;�`:�(��!�I ���j}�O28��2��r��	@w^�#w)�T�=Nv=��{-b�n�ԯ��f�]���(�Č����a=���wW�#z̻��iǗ�a.�9��G��l���7=yO�k����� �Ь\ϊ:�ұ����mח�v�|BQ������̩�l['�?���1A��Ys;��|�\G����_��A|��4��K�ߡ�:��b��?�Č��ǰ��r ����k��@�Pt��r ���-�'0���S�?��Ƶ�R@~�����^�YT/���p����f�J�% �Bk�s@���w��)=���I	l�-��+�xA���9R��7��5y�KR��l���h#D;*d4�����:��϶]���=�[I�c-��w�ϩ�瘢m㳵��g؅����*F*��j�=e[�R.�3��	�A{J�`�diV���KoC����1
��R@�37��LT�"vA��}�4.�s� M�%�?�D]�i� �A�D0p0r|u���������]��}Y�h-�d�Aڲ� Yv~�{�����;��O���?����۪V�Y�*�oFʎU�ΊVsT��@Q!f07Ѷ�J[_E��J���M<>�*W=�^D�:�+���uf
me2��Y4ee�I��#B�|�B�=�Y������%�H{���.f>h·�e�����k�'��ڔ�v ���:�4d�cn�fkk�9�[�lv����'F@n���ʑS��j(����VB5�/�Nx�I��!+�Z��>Z6�,���-�����侂��wF�#����ś���_}1�ߏ��"��}砦�|�m*�$�����<�����L+x�erf'�t��s�J`F�����:F%T�{�f�g�:4g�������ӎ�J��Ya\>��M��u\�Ԑ���ޔ��S��fiρ�#x�.6�}FAK]��P^�����K��9�z�0�4bb>�7�H6�5<�䘎�#�1��o����܌�vڼ^��K�z�_�����G⹚ƪ��e`b
HK�gN��xD��>+���q�4��C�H�� =��I�Ʊ�X���/�]��N�2�+�0�wL���Ƶ�����Q�d�ڭh�g�K?��M���3��٢�l��,��l��!K������9q�F9�zN��&d+�$��9�&��%fhgH��>�T1��ik����s��a/�07��M�^W�f�,�q����N��Uu�ډHz��E��^�n_�k���=Ɠ�/,�C<��9=��6�8��Gbs��Ff+���DiƧfT�LD�q GC�d3�D?�H�Z�J-����)�m���z�}���	GH �=�K�J@����%�5�I{, ߛs�ji����;=���0'+��	�zτ�K�lx2���׬�gP�i�%���t'x�,�c�eCJO�	8fr�f�2oo/NNoF#{wzz��!� ��TvJ �$��ʲ�Y[|���g>�������o��*pO�5���Ye��=�A'��}��M��͡�jCL���E	�`;a��SF'I
����%G�c�w�6�\G��E�&��}aχʺf
�(��'7�:Ygr�`�ֹ��	F�uz�f��(&t hD~����-^7�-Қ:Rb���$V_ې��������֓y�ņ�Xd���������a@������_�,�st*����rΨ*�p���4���7�:x�+���>}=��S��{��9���dp�vo�=�����-���)�>����Q���R:�H����[N/3��'t����m�a�TrP�$*���{7���j�K89�ȡ{rn��':v+r��}����cI
4�v���
ﵮ+4"�V:���7t�mI���6�@e+�Hڑ��L�̬%����iM]��'6��#mڒ�"�?�pNm(���6�����X�)�MpV���'=���?�]�����Ç?�vz�ա_ג��� gK�=j$��Փ�t�I�G268�a��L�b��Z8�{�������أlO?n~�#��W�bSƥ؞��ǏB�J�v�5��c�v�	d�e��D����ֶ*Y�H�� �[�1�<�	���ԆQc��[ܿ���}�>���=�c�K���Ӭ��޵��w�gox&$ k��߹"��GJc�1@:�k���1�[̀�b�ǩS?����b��M�)�q�c�4ީW�aۢ�4�ap)�>@;�[)�橿٧eN$ϵq��~Fψ_K���%�,�%�:�ɏ8�܁�'���u����Ye=��~��|̴�\�f_ZRc�c�'��b�����^Ȁ�[���ܹ��$q�Fߟ��[F�|��d�!ٚ��|��4��{9�<j �T�e��i�&��z�F�g�d�d�i6*L�/����$m��]r$���د��jbAiR�%Ul���Ԅ����Q�s*8�O����>�>��=2)^��e�A٣�# *iWY�t;yx����������=�(��9�I�Z-��deLi�wL��c�z�'I������%�~miZ��&��" �A>�(��#���ZfZ�E�C��)P�P�gi��$F5p|�X�h�P���:2:��3��,�"8�_]*&��
��Dz̴����s���ߚk$�ol����֔a��\L�~�A�(�!0����4���#{�2����ֆ'��wq%�m	9�o�䥶�yN��	nNg�gNL�B�:lV/r5��㻧�5�����5RJ����rM�����jo��z����u&]I]�����I��R}�Y��d0��p���:Y�T���Y0�:,��4�ܾ/��E	��}^�ׁ[*`����(�$�s`Yw��	8UB��S����'����3;G�H�_�,:��~��oW8@ٸ7|�w����}�F�IV�^����7��g	l���h氄Ȃ���ڄĎ�s�;C�[鹹�b�l��%�$(�#!*�hĎ$�r��z�ٟ��W��_�SPS�x����,١���F�n����e�k�:�Kjkz�
,{�`[��U�W
+8IĐ���kf:	�����K{��`�%�Ka�7�F���v<��;�Kˑ��7�� �efΦ�q�sG=�GF�<��T�钸P��-��.��rM�ِ@���H�E�F�)�i;zw�����\I�k�5�O����ئ�����`%���4��%@z�T�B�g��_\`rτbǌ�h��ǡb���9p�0l��'�9+Ɩ�93�F���=k�Ӿ��g�d|�P:#q�t�y�j7u0q?��T��{�h�!��4i��Ev��'Z�_�ʕ�Cs��e���kM�������7�{*�
�a{V�>'[��}ҁl��e�ɖ�O��џ]�쾸���Vb�.�]}FXe��@"M�LЀ�7��8�k���dr�#���h�x�����F�}��L=�s+Ǯ���P�Y�������ؚ 	�ki'�\H�I
��������O���zW���>��Y2� /S�B (jqOw����Wo������ei�"��D����H�}�L�W�*)쩐Y3^��+��@�A#U~�W[mטʋ>@��r��\�V��f§
]���<�����´6I(�����U�������JI	�8ss|s������)� �+i�Q�&1��C�E,M���w�f�ɇ�v[^۔K��5����09�_�����Ae��)m�Y���3\��#d,�v"☝>az�Z'dN���������љ�W�rR��EF�5����,���f	PCU:0���{x�sD ��0����+���~Ŕ��u���p��Q�w��9�p�)ASl���W�}�N�U7�E�_gp�E7<=p��r67����� ��d��7x"F
�qF'������ܾޖM��	�%�x}�O��~6+^ ���>P>�SRS�۸�ӹ��vR1�V��'�6=Y��cic4��K���V�O�Q]`H����F��3��PO��Q4&��R2�1-�d�MT�{�s�ނ�^̢�sU���lT��YFz˟�Ӈz�顒�>�d���y7�t�K߫)��� ph[�u.�W$��Nq>1D�r�$��� �y��4��|�Qg?3Ũ��h��c ��*8��Ĺ�����0Paөl�	�'+LG+������f>���a��.aBcE��t�ѝT*��9"��L*�s4������s|�Y�L �ؾ���ǈg�Ol?f�|�N}��6fJn ��B��/���f�My�N�0H����j��*��� ��$�?L��ɂk��3W�K�d|C}:��������ϑ 4 f/�m�,��@�oXS����`�ٕr"��}g��G�6�њ��
%k棽�[����[�}�[^A9���9���u�hľ<�tT~N���f',�P:H�lS����`��R�]�m���ԡj�')1��W;[�C�}]:Ȟd�"hc1�m�� ������5A����ߩ <r��(р����:-4� ���厓��ͅڝ.`�݊#y�hb�#gH�P�/PM�2[�����IU��F%�"��W�V�����?{�3+g�q&Mk�f4<��2��S�gd�L�����Ϳ��������]=�*�����)����>�F��V���Hq��Of�4�
�|Q�����v�z?ft��f���*�/����!������o���<�Q���]���a  ��r<�cf����h�f[�"��zH&��w=�-	�'\$K���\^��'\z̐� ��^��
��mgWX����#��l���({�*E�u��R�>:�	,��Z�N�97%�&�i�ڐ����m���gZ�1F�c���o�q+�}T�~�D���U�:�z �'W�O7f��b�͔@&�ۤ���h�.��c�K?�yH�����t<(�e�^+F������W�kE�#��l���`�u��l|f�쒝�E��#y��X��<^�6���ۂ�|w�*"5�u�}���8˩\E�yr�c?��ݰ�ȈAV�{�sd�%�Iu�`3���ı��.�s� ݼ�W�� 0�9L(E��I
�?(��D��%z�M�ZY�����;�	`8��:�.����~��c�lE�@�>�T���ٓ$����o����~�H�5���p�%�3�G'j�{#D�#�8��H��qzI�5��h?L��Z������]�-��@ơ74�^\�`��������a������`2�	�F&D����$0�K��O���]�:mD���.py���f.��f4}�4G�e�*+
	@{��czk�s�Y=��3I��}���J��a�����\��cxBRM�l��q{H���mF���	j�������<D�@���!8��\���]:����N9P��֧�26L�0����w���U���qp�������w�U:O����Ǣ�X���m��d���w� B��f"���o�4f�F���c�;�Y�*�/�`'����%��,����zh�{���u�Z����Dq	�Kا�9=gN���
J�!mĊ,g�"�X�TBE);�k��0..R�����I3�⨑�؛ͨ���X��3�hf�Ay��"�~SLD�˯KTgx8�%��h�=0�6�q�ɘ�c��Z�ob�~z6���3��M�߆kpN3:�kO�-+���ۥ�� ����>K1�s-f=�p��<�6�:�1+J	3���(���7����+��չ==�D-ke�A�)�� `�i5�����������jg��th�cb0�2�4��oND1"�[��b�I��*k���Ƀ�������&�NimmW��|����� [���10l2Q��.��K ~���a$�9�3_o&�G�ϱ�sX��	ܧ�կ�jȤ�>:)[�k{�h��.�6�1�6��EZ�e����$�8%`7����I@Y�آ�m6����(r��h�cЧ�[g�v�Xk8 ���(����^��~�#�St���պhFNS���e���HZJ��٫��J�@y����9g�rI�\h��hLl���Gb��mI��%���(҉�c�}�Q��g� ��>�b^�nYd���}��cb4���D���*��Wp��������%�Q@����o��,(��F��d�8�N+�J�����\��dB�:$��)�I��N�Þ�+�CQT9�d"�s�uEQ������i���!2�s`k���T����m�a���_�}�����D �?��r�ňJ� �]��>���G:��*|�ة�5��ٹP䌴�3�vU+:1��<_����)�W����@:��	Wu�^���u��{� J(ˊ�V<1�{9��5��c���Vn��p�Ө�^���$Z+�`j|�W��h̢�-Ny.|��R�gJI����?ΟT�y�QT+��8�V�Ն�O�r�k�9�7l��-�Ϥ1��p�����%��X�Jd����.G� u��Mm��z��q���ki=Q{7��HzB�����6��wd���{�Y��H��2�$�dR�B+�i#��@9���z�¬`����Wط������ 4��2��##2,ڕ�'��u�az�<Ș� �茢�3B��N���s������u�&j��ǒ�e����7�m��<8�y�X�	i8��̊�(�Cʮ��vA9 ���~�z*u��o��zq�i����n�J�����MAJY�����K\�]��||��K3�.��*���?f��F!��a��X���F��	��S`�(g��h}~I�WA��}�)fH�[���Z"�#��o�W8�kƣ8p���?�<����Ze��gb�F�~%&��T�[q�5L���z|"m�`��g�n����}��ڬ�������s�� �>}��'�Ǳ��6=W\�v�A�G���C>c:����f�`d�銤�֊�t�7�6�D�ۈkH�<�m4���4E��@I���X:�'�e���xQ��>��R��ٮ�ʣ�j�_�2��O�l����o��+�}�����r�|1����o1� ��)�  ؇2��޿-M������S����z/M��Dv� "��γ� z���q"�ʉ���h��0tR�m��&9�������,���E&�`�j�~���s��"�J�PpBp�[�"�p���M�M��7ИSǃ�mZj:eŨ�6q \k�_'�itOF� "��Mh������#@L�Wޯl\����Q~��>�n*f�߶u��	C�GZ���$T��ub�M���������d�?�B�u�/�Q�E�vD�SZ���ȩ�h)�� ���X�>��-FV�r�`?c:s�bT���7�&���$d��r�#At��*�y�c,[謽F��ζ��<#���>fY�t|'�n��t���D��ݧ��`��X�5�<���p__í���&̺P9�"j��J y�T�f�㵰1��v�` .n��ny��}	���g�F6{�.ޢ91�8r���c�.5�t��b�@'�ߘP;�O�c��ީ'6�S��0�H��xF݀v��cI����LtہA*��6�z�����g�z��d��Z��W:8�t+"!i]l+@�%��eE�u�h<#�w�_3��0���䀞M+��9��B�%��$����� ��?#�Z��J�U@kl|��k,�`��4F���~ŉj��s��]I��U��O���v��ԯx!h7�^Lʬ�U%�����ͷ
�"@}��3^�TbFD�ᜯ;��|i-=�ֱ�0�O$7~�zF����vz%��G%������)��Vr^g���d#x���cx�Ո�3g��q��������H�IkX��W8/M�g��s�s���6�]�Ϡ��A`$��M6c{�`*����� ؿ�w�O0
:D�6�37���
�a֮������s.��%�4p`iӖ�������\�<�LR�t(�� ����V���G.W�0���<���9��D _�6�$]�8!S;�M,����w/I��A��lrlw�kZ�N0B~I�8��L� #Z��|Q63�⼀2��r;)ڛʑd��-�s$a���LA���:���h4�@0S	=\�v-�?�#�, ��v��`���o��
��{\S^KƗ.�bs�BI�=u-=c��8��8OP��%xɊ8�oy!�ϒ�LM ��H5B�:��uC�M2�}8v�g�G-��P,k�kƏVK����Iy��3Xm)(�yݾq����V��B�ݥ�g���N�m�-�f4־���ɶ�%��M<ǧ�_G�ؓ���h6���y���7_���{���i��c��� �2��5�\��>�<>��7#�}������ZqV���JMM I��@�]��S�h��D�h_�Ӻ-��7)]-=��b�)c�D׀,F@A�0��鼶 �E��7L,(��<�����7��qF�US�g/tki�����$2�~Kg�����Wz�����t�Lc�oNҚ�'z���{�@�	tП���C��^*���b�*G�9�o��Jb����E:ա�bđ������3��sJ!�J������D��D��)G{��WA)�HBA���ͬ�bpWmB����ZKL+[q��G����,��u�/�9��1E�b��HT ���N�M��(���S_�0�~���Cw����0#G-�MSJ��Q?�u��c�N��]D�dE�n�|q���N�3(������ًot�M���Dq9�:pm������U�a;�&�N.dc��;�@��0��Q�s@S�ԱIY0�u�X�,��6�Ӥ��2g ��4���ᴮg�H �.Wi� ��@{*��I���ܼ�ct|3�T^����z���>���;!ǧm�Ѫ%��OFa���b�b ����pqW�}w~�c���'�+�k;�_z�C�~"�+,C�*.,݋�ֵw�X�k��u����J|�y�R�f��#q9�����D����g�?$t�Ӡ�_����q�"���PRI�O����S����o�-{�Z�s�Č�(��Z?3�p�.3�VFm!��)������3��tT �Yv0�s���;��g�l2*�T��mB��%�ge�=���-� J���{ ��
�$ <^<_Ȃ��K�Q̃e[��v�T��U�fz��+8VH4c��5-7D��({*k�r���gp���<�c;�ep=�������M��z��fE��7I6�-�5��QJ�[Ȗ����3$  i���G��V�	�3&�k'h�l�k�V&\s1IHH�C4h���G���HF+^���_ �>�{�����&�%�0��4@�{���L䤒�M�5Xa�[�T��fW�������`�{���;cx�՘t��Tu�g����*&7kfL$��2����7?W� /@"�4������>��~Ӳ�mH!��%X ��$cQMa���	@0��;�(ٙ�����i�-��o���7��sB&�R&� ��Wh��uR`���C�q;RR�:R�;/��r�U}�|�Z�Jں�z�)g��R��Ӈ���ߏ�}-9� ��-��  �쇿��w� ø�\7b,e6�^	S�O��Q?��+͞KҼ(�ތH7��"�4��"@�4M�M��l�i���QgV���4b�'0��xʒ�0a� ��f[�t�iݜ�]kV��:���OK��л��������o�E�s��e?�;�ct�QM���=�҆u��n��`���0���ҟ�cW�Kjt8E����C�HҒaI�ҽZcpF+���0�;�����it� ����"�TEg�Lu��P�2 �N�__/�/�f#:r���������j��.�J)��LR�j"��b=�sr<��˺�}�Q^���U�"��q�Z[�6'�czO��<�����˒�9����@�R�/��`�Z)+���l];�'��t��$�S�^f�x��9���q�8Nq�>�p�Y$2p���W�s:�N�1
��Up�q#Q��I}*ݶ�Ը <�l��/f����#��+�R���z��c��g��q|[�q|H!�[����ͩ���Fcǵ�%�����&���(>ԧ��j�1;e��f3.�r�nZ������;w�ǃҔ�.Ȩ�λNJ�<���f�A��:�hW���v�"�䚂�#�.���/�6$bD5&X����k8@d^9���h�1��9�ѳ��	�A�ُN%+��ì�a�����
��#螳��Z�����Wf�v�Ǚ�vA_�C��kq]"Yu���|�ɴ~=���T� � ������a83��>c��'�ѳL�c\
��lR����H�#Bb�"����E��N��6�	�Q!��q�'<?e�*9{��$0������jvf���5&������~@�W�,�n;�2�N]�k���I�:4  ���6ϙ|�6﷾{B���'D�u��xn��E����� ���}����/x-��
���;H�*��$H?�q#��+0���ZB��y$e��=���������U��u/��b����1�~���]�H�$;�<��`؎AB#�Qh'Pv��Ǖ]J�܎J�����=�B�m��@�K@�
��Oj}�]�X۳H�B�m$c�f���B�Mm{=�nR�8�uC>���#���AY�]��skjk���	�EBYN3��k�c��{���~>b�ftm�{6je��>�_:IHh��,HR�50�ef���=p�ᥭ�]���~څ��5� ψΆ������3m57���>��𹩀3*�s���"D1=g�q�5ȃ��$�l���F���&�j)j�b�9��T�&�PL�&�.D�F2B�y��1L	��N�A�J(�-/D�:�Ϝ���vT������ ��KvM  �������7?����|*NƾV��#�y�&x,z�����4��#O�2�t�  l �c~9���&&����4���.4
 �d�ϱ�-=����1��h�'���\#��� p�dמ�9������NV!��K���}�Ob;�Y���n~��w���<��zkɡ��cs�m*jw8���\��oψ�����/t���Y-�0i�����O�Mc)c[k
r}6+�E��GG>�D ����T�ck�k��ޝwbDb_?=r9҉	�����{��±�*�9ۈ�w�gB�Sԏ1ص�6LP���Y����8b��([�?.�1�hSi�$ɚ��=Q�"������Q蜡�J����z��B�J���\p��D�Spf�T���1�,�:g�\6�)l>g��F!	 �=$�h��!��L������u�����t��"Ϩ�:����:���="�R9��H6h���j�q�a�qN;�`JW�RF]�N���3�V}���3�T=��x�N9�VKj�f.�RƄu2J0ö�t5+� ~�i��9B2�t���.�
�7���	 D���%<��ױ������Ƙz��(��٩�չ��O���%g��x�9ʴ�6��&�(9�P�J}I����.o��=�2�9�8��Y��EQֲ�i��U7D���6R��r�>�� >֯[���;^��ȮH�y�l�x�K}Z?	�:k��=��/~����㔃J��t����.��d0,eT� ��P/���:u.��`s���]��&�A�� �kU?�J�sA��Vg�6����N���}l�t�RK.`*�k��g F�"Ȋ�C�Y�$�� �M������1�4�yPU�̼׽�}9߹���qs3&��� aP.2�DD��I��o���EVD'��HAH!��� XV�������;߷����^f��^��U=�3=3=3=�u��ޙ�����V�g]��B�������^^N��!^I%|�@m� @O��rw�%-����3�~� `��X��A@u��a�B����?����@��=����'0_���x�Y
���� 1����a����u�882ó�D(�e��G�^�?x��'��'� ��?: ��Y�*��CI�@���@�>�.�e6���/dV �_���dM�6>�|43���+����Lf.�#�΋{'%k��7�_�|f�^���^�pJ߅�~u������e2F���߲=_g����q�!:���]x�������Ϙ��$Qm�}����=���*+t�
G�=�*`)����D�{��7���M�`#��ƈ��k8V�ئ1��s��A�]���.oBo�pɺZN�S<z�����g������nR����W�L��F�� P������g~k�շ>����}_,|	J�ĳ�4x��d��U����hb�UE�W����!�^��b����>1:z�r%� ��b���B	<��F!�"aE����8I�+CPB�G�Ϫ�������M�����j�]	X�f't��6q�H�����N;�ǆ�g�SA�q�B�r��p�����ѣ������o��0�H�����z�Еg{#X,Gȝ��@C�' ���ذ�~67o�OvJ��^���D���/��s~*3�
G �bb��Az�)�T �c�D�*"υb���F]g�˜A�F �S�ɛ/���j׃C������ o��ד�95�+����O����	)�Ps�@�����*�W>5\
x���V^�W6&�1���ѾW/&�	�qH�����,d�xĺ��6&��㜨葌�G�H+* X�U2V4��m�a����A~���w���R2�!��NWhDG x��̄������9�!���n��yd�r�X���!�r��|��)���26o]��K�G���#9!����I�'>��(< �a@��Ҽ����
f����ٳ��Rכ��:yr���Ʋ����r��g0���nf�h����ҪcV���bi�{J}<��pW�g��.8���3p���T�S�6e�� �Ez�Ϣ~�ix���Z��*w�������9��2�SfW6��@2�.�%�&qώ��FG�`J��־�����]P�B
���_߅�~�f�e� �W ��N	�Xơ�� �,GܖL^��j"���D��<��z��k$�8:��9�AưW_93��2ô�W7��4�ҋ�q�e���SZI?"�Y�j~Z� ݆����� )��J�x��J�?,�s�@�}�uJS�Ȋ��{�	�p8��.d�Gx樿���ݧ�'Љ��#�K��b���k���w��
Y8.��!������z{V��F��-�\��$��	��J: �� ^�x�����	�ZQ�-�h���C�zU���<���z~�0� ���&3�%z��2J���������_^p�AW�:X�$Ҟ���m����匳^�h(h���-���$���޷U��L���y��hݳ�A4�#C[�kB�|b���4�OJV[[s�g�����Ip��P��`�Q��$%���'�A���tPU�K�(��:'��J3JGC�
 �R��	w��^��R�->�/(�f���e�S��'���˷��ﮮ��&; dʔi���fFhV��/Ϟ}����������_��������+h([.�L�n�B�2p/Zd6	c�6
� �)K�*�b� �:J�B&�D��Y+� ȏ�Av��7�I��{ˠ?�^�e9��7\���J�,cǃP��)�jAp)!�9�KS�(ak�s�c1��P�UiS�+��p,�2'Ov�B*/#Qj[h����lb��W����C�^�k�K�EzF�~i̢ެ��(0 }�i�s��!�Ɋ�z��i	���w�d�6��3��w=����AU�� 5|�zQ}��1�9Fb��B#���n�!���;18t �T��!z��� �Z�6�lI)�Ĉ�¸B���
Q;����θv���\�QjК�m�ް��>F0=�\3\ �ܿsh�X4J1��&�xc�*`(z��'Hc��gS����a���#�W�@�c9�+�zG
��#w*�6��K��2�_O�}���w���`�쇶`އ��f}4(:3����+x����"ԁׂ�JX�:F����i|�	�s���[`�m������8�]��SF�!�1l�_���"A.��۷s4���)�~|�)�
��Q"� �,�S�#�,���x���\���I��
X�����:! ���U�<��]�A�-Q�G!|=��G ������!S �� �)�|�O)�s��Q�}.،����=��z,����a��X��L ��'f��5:´�-�5�- �òL�����k �/�P� y��k����ec��%���%�����~B 8�<�Y��� �{�el���!!�} R�'��c����������e�L]ljpf+b�,|YF�� �T��_|�ܼ���_��C��+�|[u�ɫ�<�/}� |v$@><{	�q���b����m� H�ŹG�nّ`ۗԧ�@���i�_��8�T�u��\�"�����"���z��&�AvAp�[P���WS̪@��L��Io<�%F��u�Q�yx�!� ��ռ �XI�Z���@bK�#R��>���Rk�86p�xx�@��k�	`�����/w�L����/��E�`>!�2�|���G?pan^S�)�|&m{�͆]7��~�|��(cT�����0o��G�N��`��Kr��Yg}(���*����.���=yƼ��ػG�S�t|�u���e���O�o9�US����$�~%�>� ����zx�@�Q�!*߈Á�}�h�S�2��*� �_�����? 3�������#��@ߐ��[a8tOmA��I���������&��EQ�s�3 dʔi-"�|||p��w�.���_|��O>-�&�&�AmϠ:���{Ź�Ә>�7�F�3�G{c�gc$��0vK��W�E�D�� ��;N�A�IQpvvrP�{�L�O�
��r*���9j��0�����[E�R��Y#ړ-G���T���A�wlی��2�#�<���R#���N3�^�}�"H��u����a�g�J(J�	�d� Ԃ7[	�	��{W҆�7��C�g�ڃ�##�k�p�9�,ÿ�gb���?�����8*�r��bg)G�I�'Z2:���R!��9I �y��3��3�.�����|���I>�� �9e C��Ϧ��gTO�r��-s���j�����2N>�ԣ:ͲE@��3�B�ݻ7�����߾��q�˾��^+N�Z��rlC*�&��36�IM�����H/��$�hj��z��	i��o�6=�3I������)f<�	��Z�щ�ec��S ��'�v~ד�g�fT�c�Ȣ��Pzg6���D���h�j\�%�����)�#XVRO�D����q/S,2��.�hc�k�`*o1������{���^����K�P������ �;�d�%�v,�!�֤�{w�� �
�� L���Fݬ`g�	� �:��\�=b�����IC�k�)}�"죤���N��o}x�P�Y�0����r���5�z�!
�b ΗgX����c�����K�|l�;d6;���}�%���g�U��}?{YP� ���K���gn�#�����T�E�3h����c��[ys
r�)��6m����5�)F�VhA%*0+��6r���-�A��R6�"�lL�!��W=fpp��+f[�1����|��oB�mF�����Ӣ'`I��	��@����t�0o��赵�@٪�;�y���[���������^���K(m�������]l��u|�7X�R4+�����?7/j> e@G�6�h�Y��I��<IE_�J�� �_�K�#��IrE;�w0�Kb���DI���
P]>��v.f��xE.-��'c_�)�`=���e�����&�(��C̰���U��߹O��wb�ʔ�u�Q���ɰ�~�d<��^�*�_U'X�W�ϧ�z^�
�?��?~������M5� ��L�Δ)S�e:� 0RW������_��_w�ψm##�x���c?�y�[��l�f"#f7��US��@~<R�pXd
@'���w��,z��8�*C�[8ҟ�R�b���z:�dH�:�t1�~���943�95a>�a��<�:�j�?�,�B8��EO�'.��F�S ��Hv#̒8���@B׻��kr��:�.�|~Z�a3����������7��&���!���:DIB����6(:7�M�3����`1�@	P��86�7� �M)��m���f�Q,z�����_}�#����yJ�;�����x�����߳T�2D�����M�lq��71�%�#WP����<s��%����G�<���Ɍ28��an6�Qb������en^�����#�d�������^рc�pn�Eb������C��%'�M���K���qJ��|d��7�6����"�	L%�����&0�btV�q��:�3e[)�w�hft$�:UT�� �:�I�����S���R��-�'#%�ULK-)�'�
@�u�NnP�P�ǵ4�N"Y���r��k��>�/c�ل�Бτ�6˺i¹��
X�E�T� �����( (ǫ۷�A����z��� cA~�<����D~�1B�V�)g��Z��I�oQE���%+.����9��	6NFB��'�	�b�=�_�;@�&�$�Q��� �.�a[������l�9N�8��9���{�:���`��ѽkp�  > 찶�#ޓd��瀲lB��h wvK~')����3���K���W���)BICc���>H?�J}' ��+�%E�K�."p��~%k����<�n@&��:�q_�nԧ�����H�~v	^^� 2�-�c�
*t���\�Ms������%�s�φ�V�[�o� O�M*�Gnԟ��l̴	{\�BR�\:���%P*��2tj�+gֱ�+\e���l0g(��|�{�	�^�!�Nc
m�j>�Mt؃�m��/�v^���`�B �s��@�?�#��jd����^{�ҖO�	�L���4�5s�$���Cx~�	�8�B�E]�=��.��3�#�-�� ������7�*ݒ8����1�ly�����f?����W��J�p��o�,u���79�_2@���`ߐ̶��ޒpxg��-�]ӼV!G�C�!̫8-���L������^��`�j�L�N�� 0�L����~�/�ُ�Oʫ[3/J�iw��l�dZ�`��3��t�1 �E�9h�l�MV��"s�FLc��s"��C ��>̯(��M�%��u�4�F��:�)v2��[�cc��{3@@р��� �Me@�U;ȹ��/�jT�Ή�ǿ6k�GӃ��z��,J�d�cH�瀑��	0���� 9�;Rq-T����ȭ�tY������w�	2�<`��ǔ�h��c�NH���~n�X8ܾ�w�bSs}3E���P��]G��0�ș��'l���A0H5\�IE=�9��q��J.�a6q�
B�|���mf	�Ԟ��G�����<�1dC'D��X�K�B����Qy<�\��A��\)#\��K0�p��Oq�`J�daݾ�Ǆ�ȥ����qI�L�� ����9�Mp�R7�BA�nY���\���f��6��P�����}柁s�G^zW�}���&�,w�"����f2n��K�� �{8���0p�T��є��7F�L2 ��Hz�W_��0B~6{4(rk�6�r �D`
��!0��c� ���7] 4�I=ʞ��+�:�DafQV�f ���{N���a*�{�;�&bp:>����@����o;7��|n^}q����Q��Xnf�~x�:�-����m���!��>�r�H���Kg8^�# 8��~k��C��5��H�,�r�� ��_~i������Ŀ|���w��>�6�v&�~������Up��� ����!�����306 3�~j���^�Yײ�̑�C��}����	C��7(�@��)��y^^;��?C�a�3Z��(���בm���dπ2ppT���xz��X��ma�D����g3rf@ǊB�OP��P�է��*�����K-�L���m��R��9"�"4݈����H�2�%�8���6e��[�_�4ط�J"�U������q��b�(��y�_�� ���)���}���z��mU�E}��e]A�����=���~kvyˀ'ƌ-ϱ�RV��3k�}�����@I)��Y��-c�5G����ݒ\mAx_����\�.������g(��}�~�g@I��3=��`����e}y�.v��n�z��E�g���C�a��m�V�J�G����9���!���+B9a��2o(��WN\�.��g !����qGL��2^�꒢?ޛ8H���A��I��#�A���D`��.�ĳO1��V1����D���0�yL�s��ݽ���v�V�����`�{�A�L��>����tpo������_�������f�ꍡ�hT(�����c��Յ ������P1B��26DMA*~ тV(��,�3블U��2|8(��P+|%�g�m���������EB`Q��`p)A`�L[�^L=�������~\}Ma�Du}3�]!��`�>J��7����>��$,���X�>|�����L	���`���"$��8�� =Ŵ��	�hc'$\Wެ�ǹ��?�W���
���O!g x苂gq�;;�/:��󆝌g�ɯE'\X��Gp ���3 Ȼ��{��[��6 �0oqx� ���Gg������/)��3bn�0 Ķ�sP���3=����TjNc0
����I�"g�����+�=#@zF��j_{��1P�$tl�H����]�8�� "��f�i2�G�I6W������I���=��tI �?�����@��g��u����DM��Z���{������MW�ζ_�����?��* �`)oB�Q�q�,��W!e�؈FD�0g���D�O����E��m%[ �^�iYr$�DQ�R������ř�1P\�z���.�s�xRP�78��hf^�@��Zfa�b���Xw;��!~�U����%�ىe]�JA<��H5�GD�R���
z����~�R��өA{lH;Q�
�k��[���)
ֿAƁ�)�i�ap�����o��)kԗTg��`&ԕ��uL�{����yV�ɫ��p  ��g��"���T�lɱ.�L7l$+gJ(����a�����61[:��Z���,�L"HJ���Ñ��㿳����	 �@��5�*vz@¥S���˸����9�ĹS؟[e�2���qp�[��p��1�� �?4vB8�J!NLu!�����G>��4����# �kε�Af:��v���%l4yvU�̀��,�Y�_2���X�hL�Y.�1�̘�<'�Z�g~XKTS�|��d�2e:1�����A�v�e����m�GR���Z)�o^�����d�hu`�Ox�=dga\C��3	�rV�x�̠�7����C27�\����$+�v�X&n<�?\�@��e����G�:�3������?�����?���c���z�������ܰ�j�L�2�Ѿ3  ?+���7/����~u^T?X+�������Ȋ�%�����JӖ���7d\����8��,�vaT�H:~a��`��2`O�F�k��2	�-���n��n�o�����x�i'�L"�؁Al�s$��^�����N��]	nm�+��s��om���J�*�)^�4\��h���onF݃(;�O�[��!6)c��qtA��_r #n�EYjn�4F���͠x�c�ń���5՜�(J���&՚D�)�^N��ҤB�<� AE�����N��`���X70A�ɡq�*����a(�@��`�4��B)<y�l�kY��P	�C9�v��ETԡ�6D.� ��}�jjC7�{��Sr���*�,�Xj�d`�'X��,)"f�xa��(��O7]6�Z��/�*CIki�Spڴ��n�`(e �j%s䐣�H7Z���q�`�J�>�g(N����ggd�9Gz�<�yIA;�M��1�0v^�H�ZH}Iu;1pR(٘kFD�M@���bTe��ڰ�7l�uf�+sD`�AG�R;r�;�5*�0����&�� /��e-oo^���Gg����I6FL�˖�7EJ������ZŵQ�dR�[�i�D�Y,�d�c � �hIp�)+��ZM�����o�3Z^��4�|�@8X\���1g*9�r����&[�\�B��Y=�nBv�X�M�����e��3��Dӣ��e��uV
�߶g���?�f��Q�9rL�!P
�����=f�{&̎7����^��;i��AvQ��ˁ< gp,�6����;?t�?pN�=Y`�|^��%PW,�0뚳�V��1�O�c�n��jgC����RR��W��3��-b��fc�k��xfg�lwϊh?0��r�V��P����m�,YqM�>���]^M0�/l���v Ԝ۶q4�k�}�Q�yJ'�9r��jn(�
����Ԃ^~�| ����z5��>�a{R�$~�#mf���n#A�b珘��76������Ի�N�q��7�8`0 �y�L_/ǀ��Ȧ À�蟈E1�l�V"��ֽرE`S��X:��˲��L���Q��4�S1�<��,���$򥪕��f��ͭ��z�w����}n����~�֮�}����$u^�L�2:D	 ����<^-���f�S��"��a�B3��!kV�a��Ƃ����!�VD��^��A�e-b �w��1��|�a��̑�:�J ��^<������Y��k(��x�E�����Nn�0j<���dKH��t6�\��=ۺ�&8�,":��*��:G���i���~���p��!Bm���1%=�;j�O�@!�3F� ��FC�cХl��N� S�7yYo6�7�h>�:�P���(Tt�����=�ͥ�M�M�9���ԝ`��lq�M�r�ބm���f��g�]a�ѓ��@a�i��� �3v��e�ݭ�~��[��1��ry2Dd���ѧ�$Fu��	 ��y��	�H�q�!&�>��$VH�O�`tƙ��ה���R6g�$�z�>E�ˁ��
Amaxsc�&I��nkl>]��-i�fWoh�۞��9~�������:uȺ"+�h`��9��WA��Vb��0�=�dd&8ѕ� �	f�wG���p2�r��Y}��69g#��(�(�w���3��������7��p�Υ0���#��T��0�"_}F� ��O����i�s4�k�ߝ�ly�	; � �˾�' sMk�������O�KA��  �*DKbV)ph����5�I���g;]����wS��-�"����U!M���"Pk~_�����H�����R �A�턳����[���a�B��=�i�����N���ژzח=�yxT�M��3oi�����-g��~>1�=]b�� @����p������f�4��Vr3�=��<�fZ���>���Q�m�(q��"�F�z�B��2����!���$��*cf)#�'�Id�ԧ8k�+G�gS����C����q����؟�MJ\��;��x�z5I4k���^?����S�O��}�r6�,e�;��n�t����@�Z�]�x�����P9�z^1sׄ2s��E0��~j��Êݞ]���\��Ұ:��W�[�]_�OXW�(����w	�Il���� ]���u��~k�=�k� L�d)� ��1�s�	�(l���8$�H��'ѱ@xa[�cj�p��=p���7�B��/��f'K�Xx�!��*la��ks�������\�2 �2eZI�p 0�-ݢ\��\��ۊv���.��(��OA䔹6��G�ug��UI�k(��Do3b�ڳ��7A(X�]f���	8d�c4����za�Z�����	{�qVR *�b����}X��e��
�_�,��w���CC�N;��=ld �
�t�Ě:.�#�u���LK䥮}J���ɡ�ژ��PKc.<c0-$�!� �ѓ�q�W@�	�^ ��<���U�����W����L&�"���5D>L(��ڇ^ϊ`�1�O�$� �e��:� ����l3p6�ӳ���%6�L�Pd9���W�)��_ ˵����G#�`�(�`����V�g2�$� ���3�~��X�T RO��j�&�g�X�`*N��\Y�{�?]��R�� >�  N@4"�^��#{A�J�mc��3�-�~�P3w%Y��V�i�����X׫����̈́d?8LY�R^��:y��E�_�NuRb�pZ��T�g��U,k�(��;�Zt�.���<CH���,��X^���a;+��u"�0ŷ�Aή���-B�f ��=��:��,��C�+p\B��5M}��=�I6>w�'(� �#��8���w��uF�Z�)�m�}�]��
`��4�ঞ��=���;ٱ�P�a3c�	Z�bg��'V cҿ�_xtZ)�]l�[��=̪�{�����U�������8�dw�a���cf��_ʑZ��{�����<��,fw�L�9�!��e�ݠ4���H*��L�����
���S����^7�����"��"��1������Ӑ�̾,�td�	�gh��xF�E:�	������T� �;��c<	pĒ8�����t�?���D&��3��@_��f�t[��k�]�׹�4T�:GU��һż�|���}���y^��2eZM�p ��?�^�������<�Ϋ���#��֬�0p����%���i�F�#�A�r)�1�B�Kmz&"\$Ҳb�ԂǴ"�S�j�v�>H>�~'�����낤�dp(�x��f�"!P_\U���7k�hg
9&^od4��������c�.FLEY�S���烀4&Uj�Ж�FG]c:��=�Xt�m}��N�
_�u�A~�3UͰ!�v��	��*�����%�����{�i�UZ��ޝ��-(��5-�����?[1&Y�=�S~����V&D������ș�G�EѢ��r=�&	ǂN	��ã�;E��4h4�O�9�ub�]d�:�c� x.>_p!�H�o'I���y���IK;��͓�[pj{t$b@"��(�({���b$�Ï;�p���K�(��9�b ��hHD��=L�\8N;,��-�yS��\�r<���L� ��=T�$ �X����bqem|�bݪ(��%Ԛ�b�ɟ�I�p?����" �c��sK)��Dt]��z��ŋ��:�Q�M�X���鴤����U���i���Rp6���*Λ.��ҒJkG���V������93�t�+ħ�Є >�Wå�`�Nxo&�;0�9mj�ߪO?���y�9vd)8�(��_Nh^���v��G�}��%�l�J( ��~V�!E�Wc���a�WN�B,f��+u)O/ǣ��a��4
fx)�,?j|�jdX�P8GJ���gȥĳcz�����,�8=�ϰ��Ĕ%�����7�c,g|�T��C3_�v:���������\E���a���rA�7��M�p�vi�[��Wg_X��?�S�j6[�����3eʴ��� ������?�����������z�y�� {[�J|�l��X�G�3��x�6*�mj��4��9e`0Q��Y%�}k+����Q����i����>�O�1%�1��{f��B��G�;V��d
C�}��P��c7��,�����%��Q�{���
��)Aul7�!h
_���i�q�*������]'~-~���̦�^q�PŴ�3�-˝�R[Eb��#1��Ǫ��CEܫǅ�ԩoV i��;�o��v��p���3���d�3��}��Ų�bj��V��+If�X#e�x����*���A֬6��D��1��B���F�&�H�z��F��>Jk�
�+�T���C��i+�S4DO�Qp2J�pF�n�('�*�AJ�'��2�r�:% L���S���Q�Iֹ����Ȯ>0����~,��~�C�Xo*F����<sf���K���/����]�B�G�] ��q?ҙ�=� ���K��N�[��?%r�W[<�m�m��[	�YǠ�Z��M�a:�ߘVM�r�}��Q�(�,+*Kħ����U+�-�"m�[��-���G��̐����9L
Na>��U�Va�������	 �C� y���d����6�d�Rv(��h"%��f�Ib{�3�SX��E��}���Ҷ��6}wP���?���\ ��A�g���1�Hp�S�x4Y)Kl��Qhj��7AW��|�o���B6���X��Q_�D)b��D�4��_@~�X�t_��������\��T�Ջ/|q�3?��ܟO�z0fL�W3e�4F:H��iq����?���|���z�������|�	��aϩ���91��:�\���ߕ*k��g�l��%�QLЛMh�R<Sm�*x���w�c�d�hX/��"�={{2����ܸ���@<���=��b$*(�$\l���qh��d��`��o3C@Zr~W�o\:�R��� �xݖ�,ΐl�)1a)�:c/���F�7?�u�N�!w3���t�|L�?��@
��e ��Aa<��v!��Fb��"���.e)��y#��PBo���@�kܻYY'�r�	�-`^0:����j�W��U���ok@l�k��E��FG�Gq�f�N'��q7T+ͬ_���]��N���~�#ݗ���u@L��!@�S�S �ǾvW�'�i^ۜ��Z�f!l� ��@��"�2�	�r��`�1Mc�S,��N�����2}��.ˁ��a-�87�.�*���W|;$I�k+6�����@>���@��~�C�q1c�w��@�����D�'����
ME�}��F�ٵ��F�%�FwR2���ox�Y>�
)n��߯<$N	R�>U4�و�BB�����L$��<���^��~��?�c����%�?����j=m��V7�{�c�I����6�O�����Ϫy�����ͽ�&�h#�ǆ�lH�ɎQJǑС��OƝX�8R��6�2�Z�ٛ%�b���k�M^�����F��Yw�һƀ��=����20���F���߰@��1�7^����9QރӁ�N��8@5�p���0�'OA�Ql2n�:�/���_�÷�/���m�^^��!�L�2eꢃ8 Lӻss��������_�?~�Å/��*  �o��b�@�Ѳ�5��'�&~`abc#q��_ҫ���>��Y��vY�ܫ0f��}��5��T0P�金����
���;G16�k���r�07N�5Дz�FC���<��rc�mxF�\@�K>ʨD�m�껲tn1�t�]7_�jw�����}}<1�t�ONi�n��7�ŋю���>6��umD�^�J>I%��X=�r �h�'\������}��=��j����i��.^���c��5߷�����&٨� 5�S-��WҎFN��]�X�v����W,�� ��f�|w	g`0�����?}��y�6��S!�s�)�4'��?�QR�e���X���s-pM�%	�FG��xt�!c���J{M�P�K�M-у;Q�뭉я�<!�+�ϚWx}�^�7�'��6�gBz�����)��x����x�������+-{�����{�7�e���	4� ����w&�-��hO~[�o�2��j3�Z�&J�g�J �Y��t�%���S���%=ѵȣֶ���V6�1�@ �d��m�٣c�i���\��V�LKQ�|����lM�{�������83)�ιw�\� �2eZK{u �$��ʲ\�����G�^����W��ϫ;�t�l���N�)���D�	� ��km�%��U��/7��KNhׂ�[J�i�1�UQ���6�GF:�NV�x?ҧ��$�3�AgL����ʀvx<���S�.���l#��2@�mi3&ޭ,��e�V:�F(�X���mZN����LC��m�[�]K����ڑU����"�V��h4܀x(��K�	�y����C�q�ƮC��]h�k����lF�0	`��Q)nrO����}�G}Y�
l4����>�����2Z��Y� $�D�����ƴd��ޥ/` K@ ^��q���䩃ӷ���)>tt�AAy�=n�2��oc�:C�I�����!��=?i� �"|��S%� :�6��/�4t�x�w�ϕ��߄_D�Ko�7L����F��/1�u�h��1pf����y��������|�oj���l��>�}�ɳ0��u�L��]�R��d�Tppq�8G�	��`ic8�2q�T �e\D�q�8�rV�JI�/��R��wi%����Ix��`��qCON �
%
��*���l&� s�}e�e\�e=vg������/��B��O���GR�L�2e:D �YK��o�F�f��ܟ�ʹ��s���.��R�-L����VH������� �H��֊bƼ�X�����1�1�L̢�v����
��p�	g����9�2)�ܲZ�>��M���A{ä��0(.�����`�
�o�Uf��S� :�L3]�6��3e�R6�����������@�8�%�4��3vA�y�ֽ��:Zr4��a�	�k�w�xt ���a=8�8��R��I)��w!�^7�1�SX �����6�g�k΋A�i�>Ui��-M[�֦7n!��`>���ǎ@Z�t�3mL�ނ����{t�����]���˷n�E|BSы��[��C�ԥ��g��>�} �C.���@}�N׽?�_�:Tt]sh��M�t_���5�Q�b��LG%m�*8-�KYzm�I���t�1;��&d��X2VۣR˂]��)��Ŏ�8i_m-a��(p?��x�l,���� !�t�jz��Hx��#�(K�UY�ٕ�
�o��Ag ��b� �N\:A� 橔�0ފ�NA����/J{5��Ͻ�������M2eʴ�� 0�Ng�~�髟�K�������Y8�Ӕ:ER��.�+��A��o��2fIM�
'�ǚ���1$ �����Ki���X���t$pT���uq$(y�E�1�]��@�^jPR ��+ ���>x܉ �҇����2�Ga�sg�3̈�,�O�g獄���%���^HR��|G� ����8��Qc"����h�c��H-������K=�6vzB��hȪy��Cj�3k�q_���������Ĕ��P���ˌ5;��F.���P�n�����'�����i����A)ˮL��$�`A))�G�`�4}���c?���	�48?d1�y�)��+� ����8��� ����h��m���U�k%���.�3�E�G��C��n�M�
��)d<��2�4P���P@�����U���>+~�����~�噙!��0�2eʴ��� �)��};�_����_}��t�������ygm�x\U��S���_Z��RC��w���=D����a���bo1��1@$Z�=�B�>�l n�Q�	]����{b�X.!�}�Vs��&@�8 `;��AXz�,����Nl���ؐ>�}�~�̩~v�G�~Z�lҲȏ��IQ#�Jx��mV�g�����
 J^��G��Ó��ukZJeG���.}ȴO
KԲ^`2mD}�)�-$G����{��i��E��d횽x��L��>��W�J0�ɴ�u�a)�������y�B!Xu�(����0�㫠0	�{o ��R��Ү	p�GZ�)��;Ҹ�c@�(�����g8� R�0���X���*7�@)=�P< ���e��x�Xg�͛���W~�u�揼����j>3����R �ɔ)S�:D ���ӳ��_9��_0s^0�^Y܍r�bf��k����p��`^��͢���t1�,:T�O����b���B�Ǘ�~���%g �8��x菞j�$��
���I��,{�)#\L��%��kCx�zƒ��rM0/򺽷����e����]otؙ�h��W��Œ)S��)jN��D�>����`2H���>�}@�v6�d#o����s�\nFV+l�!��s>�b�s܋���ږ�>��WO��t�Ϫ~��l4݀�n�B7��>�ynW�z�-�׶) v^��<���*g�<���]Q)��B����yͮ'�G�Zn%�v�C�\��N��|�m�9�m����sz��ii^���6�����.���8�{5�n@=�a��v�޹�}텏��m�O����+L�F���1���n�K�m��f.�4r!���:��	eL@��B|8�lJ�_qy�����CN����J���$��F	� N㓬�1��yԆ�+XY�����`nʪ0�i5�+�^���|��_������̬���)S���� ���i1�>��g�~��[?���eY�^��aaA|ܷ4!Z�>0~5N�Ul��:sb1���.V���ײ� ȗE6���1��E�(�f��w� ��p�{�����w��k9�^�g�g��f4hQ0��%�}zN�>z�����L��D�%�AȜ�v�iF��hM�Y�f�A���>����T��T�ʴ�$Uj5����nY)l4�纕H�Zm�:���^�i5	/�
6.���1!2��ېKnd����X���y�<r�A�:KYA�7yɮ'��Ҝj�����Zv>��<��I���&� (�����L}H�Y�LC�5��:�?yn�Qt`3��*�+�cL��Ԙ+��z?	{&8[��Ю0�:���/b��>֬�z�-dZ"Y��5�-�8����\ne]V�����5K_�6��lO�sJ�5�J���k3? Rs��f :E�zr���M��պ��`����1Y~m@�G�+S'a�b.U��,��S]��G���l�<9F~ق�xDL�H���lҾ���P���G��~f� ��,:@3��)�3:`D~E��UV�P�8DwA ���%ߋ�'�O��a�%�#fc9X'�8v��&��������˛�ˢx<3�*; dʔi%"@M� �뷥)Mͮ"�����ʹ��������+��2����j�!����^|�I���ţL�̴��N��FKDr.(yp%� c)��P���5>k�A��R�%���l:����h}�w]�����z.������'�th�ω�!9_ĺB2i+�YIzL;�[h��|(�A
 ��:��M��nBA�S� F9���f�����P(��1��2��hX�y��#����9UxX�EFR7�6 ň3�[Ȅ�N��_u�K��<�+��O����gm��Z�+2�ڟl�����R2u��2��E�f]\�	���@��E�W�Q�w�8�6�qNE��:�hG���	����e����9���[z6��I�F��,B�k+��=%�zϷlG�*�\�8ە�O��Q���}�ڛ�z�a��a�C���:m�Y��5���ol�,�P�֐���8|$=1̭M�18��c�!�fmG[F�3J�1����CV]Ժbv�F�N�k���8��O��u 4��,v{�Z���S�5��J
��Ms�1iP��~J��9�P��� ~��4�i85��Y�&"�J����-�h`�/��ګ�Fڐ �4��.�t�J�L���ɪ���j�Żww��\�s�)S�L�i� ���>����/��鼚�VsWy�iG.��D?D���3������C�|����U�\c�oג-�y��$�_�z�lр{�Oڊ����M�o6.� ��wGé(3 �7&ؽ�s�tH�B-lcN�S�4��kA&��v��\& i*�[�nf2�,+k	�L]��@�P�]��V����t�gè�Y'����=_ǄW��=��˸|0@'�x�S�&��F���Q�\��c��I֨M�:�S\���ٜ��3�7���\J�TD�5�I�f�?��45#]�򮫹�ߍ�k5d1&�٣��	�+�H�U� ��H7+���Rr�U70&�����v�1􁶾��6x�X�͜��8d��c{fͱ6o^�[nG�W-��Ӻ�����s�I������̫M������ü���'�=�c�_٭׷�~��j�5x����}��z��w#��:�T{�/X7�c�3k��Z7���qY�����A���m�s=׫�J���S��yǱ�����A�#�(���kw]��P�w{��`�Z2K��+\R�ֵ�}����z=0��(�����K�ms���m�S����0d�[F[��R�U�wu���c�$�~7���%��{��l��;�eE�*�x>�],ˬp��9��0��L��6N"L���
N �~<߷���Bw1A'�ͤ�4n�������8����  ��IDATΔ)��� �/������G~�o�����]��cr6��-��?X��D��f�2�9-�S@�	B��JL��S��Yb���&��N�;nb���6F7�p6���0�a�51��O%��
=���x^D��.�����؟�PA)���+��B)
�4U�r�v�y��N���N90�'.�H�P��w��5�%��[Y��c�!��Αtdr�s�5&m(�'���v$���s�Y�A�F�I�?�Eܓ�C���zԢ�������f���c��ې6�4ǿ6�3b�]�6��5ƞ�d��hX�J�zM�J5�(Y]�V*��[�Q�p;s��t��w�o��\�g:�3k�UBa;�=�`���V)�m�>ɞ�\�C�(��V�6�5{t^6�y�ߵJ#�U���W{b��=��ۭ�w�]����2�nKv�-���cS�]�n�\�Z��]�o���������5��X�z�s#�*�ڥ��o���x�6�M��!����aҽ���Cư6b����w�sh�uL=��2�����~�h`����YIc۰�7On�͠7�%%���a��H0���J��t ��nCe�gp��k�x�p�o�c9GL�oL�4�0:� S��7(�?F�vEx�o̥��0�W�N ���],>�����?�o��:��/����\�)S�L�� �z2�����}뷾����W��/��g�Z6�O ��4��\}YqꞴ^}��"�H�jl`���% ���C�ہs�T�W�����Iؖ��אV\��?)�\�!��z]�p��8M���Y p.8� �'� /���}r[pS��RA��v�T��Xr�s���T��"��6U����q.��_�_Ɔ�2�ˈF�`Y0'M�δ%�?�yb�6�v�9�&��yNdy㡱�gu��O�6zQ�M���αb�|n����<����C��}�]�Ym�Gy+cT�|v����h'���9�������<!���k�A���ڼwQ���<��4~p���Q�}���o��)���۪c۬7��X��\���t�>��D��^��z�:�r��o"�l����=��9����6=v�>a��:��|���t�m�ˁ��s5ś��� 8�[&W4�p{g��PKefVm[�ށ�q��f_���<M�x+�ćؑ�e�C� k(`ԳӀ����Aܦ�:�(�(�8���,Ȟ���DG�4sr\-U@%)����oY��-k�I*�Y�������ֿ�/���8�tꦟ_\\ܛ� �)S�5�W���y`Z���af�����/�ʯ�:�����=-�Z�����K�:0�"IY/���E x��Q�g9�K�D� e �_��I� �_V���3�.�m]oL�4��W���B[E��9(�1 j@�1QL�y�
cc����-��/�,,9H����16'M^�7+N(��ލ�j:�2 ^ݧz��l�}�W��� ���}:vf�)�z������y^�] Q[ɂ�k��U[ǲ��>�fZM'�X���xm��׶��hO�=��<����O�%�e�8�<���Y��c<���	�#k�>���Ic��Ƙ�xk�9ŵ3�w� ��Ԟ՞�+AA#k�S�A�>���7t�Q�	�{[ĺ6�l��Z�����`�)���q��"���m�`:ɺ�K�I�����<��t�^�������l6|��wյ���T��d��N��0	P�x��
|B.�ۣ���d}p0��t>">�K�$`)�{X�}�s���k1�?�؞0	 ߱��7%f�v1�3�Q��M�J$)��r aS�~�KҎ51�U�$��N�N��8o�miM	m�=L'�L�+3�O����p���5 �/�9-�+S�L��Cd 0�77s��O�ͮ>���������E��]	��T�"�m��L�G�<�4`�P
)_D �<z��� j3`�+�f`G�]��{'�޳�b�܉WG��t/A�ךF�m(
Ъ��eY�	�� �>���m���M��^g>�e�9ʸ��)��CLĺ���X/(�W�} /�im� ��'kN��Q��'@�1��B��UVov q�	�x��<�C��M���}�\�������/�:R���36��浙�#�AoƠO�^��vK
���pf�`wJ�U����l��Fߕ%� ���(�'�O��^���I��26Lg]vG�Z�:��P�lO�\�uKlS���L<��eeZ�<�o���H �)5b�q��$S<ϯ5-f�LHK�&N��6 :8/f��c6���-���&E�3�R�0
ǁ���#���B �s:��1F�I�G�����MU�$�7+��pE�A���UZF_�*b$2m�����$�I0���sJSnQ��ޙj�n2�̹�̍3eʴ�� P|���f�����;_��oL���u�>*i��(��++��'��	�ч߉��B��L�2�nU��eTJ������T�%��/��kqnK���� �k+� P`������ɹr�p��m�/��������(x⼚�o$������ê�Kǡd^cY�����)��9*1���)�߾H�VR�	R��PcI�*�S��&P���=K�1��&`jņ>�/Q˺é��.>έ�Q����t#��A^) ��lAA:k�4|�Z�l�_��w9dB�G�`�s�V�%j�W�k�� *�˱�� �Pa^U�+1F�nP���+�-�
^��V������@�X�L&�6݀7��O.)�u��q}��ej�Zgl�5ǔ��u��a&�=X@��^_.���E�VP�nJ5F�N�LC�ʺA75֝����,��l���N݀l1^��۶�m�m2���.k�'>�Z7�����ͼ`i�
�>�oՔ�k�6û^p���rF{ �X���x���\�/eͫn�2U��F���K؅�f{��{Uҙ?*$�@`��!:��_����
Nt�._ x�ض�Dp�ø13uE�ckf��s��J���?={����|>��f3g�*ϔ)�:��t:��>>��O�ܟ��ǳǫۢ����~�B��1�(�.�k�4�����CF�����I+�+%@�8� 0A�X��)������('���1旋҈H�����mv�����(#8���K�v����L�ӫ�~�:S]�e�x.>T�<S}n���M�GK���6��*B���E<����j�k?f;α+��.���
;(D� C��T�l����>��r���Җ~�Ek��>|Z��5�s�X��+|$�8��$\_ާe�~�-G�A��Ǜ�d��:���ǒ+�<G��_)�ts�w�>���i#;��d^��9�=�Y4��_�4��z�G��}���Ҷ����g����H��� #�j^p�����݃	�A)ҳY1T�$��<���}x�p|p��sj;��aR����Xe�F��ڕ׮��4�=j������ƲޅS*[!�f��z�D��6��e����M��
s�u;���"0�8�=��\�Vk��޲�'�,x� K�ҟ�c���=���b�G�״��ؐ�^�'��\�%��5�|v����{އ�ze�
�61Ųؐ�^��O(Y7hzc�hռ�g�w�~��^�V���  e��5��m���~�؇]K���6v����>)��V`+��&ؖ��Ut���^�b�+l�}:��c)�Yl2&��J�@i�z�����=O��=_j��	��6.��֦��C�<���W�K�B0&s��;�XX |Se �Q�eXnI$�/��}�H�'�*���,����@�����HK��_L��T��L�Rn�gև0#u��Č�(� ��빰�G�B4����XP����p�/Q�=���������?}s����>�0�X��2e:)ګ�'i����ş����W�c>�m�g��rR:�XX��b���z)���������T+��ݧ�>��&2s�`	t'a���	� �W�Y�̜2�tsaIHPf �F)e*�&�"0�(.��4�iqL�9ra[��4�/��� ��<{u�7]��L̢���t�z��*x���!��o�Je�O�n��:����j�0��� ����!�(>qm2D����a�뇽�v6��7�Z2�;u�y��56UzAt��Co����KT��`oÔF %f1&��}���0�lB~ݏ��$��� Y�<�ѱ"�y�~c�c[���|υ��RҨq�ڲT�����ECΧ���΃ �1%�z�{qT������v��ml����`I���!�x���XJ��f֊}�ڝ��!�oQ�<�O���d�D�/E��a�|���y_jYsV��,���E�B�2]�t�r��1�C{}|�+-��I��OP:��e���c��C��Ԡ��b&��!�}\�	��`��w8���꼡��m�8��Y9���
:k�Y������Mh������V��Z%R=q^�ݙ�omv籏�zA�M�*{ښ* TqrY�+^��1�V��hW8y�Zv�j�<�yl�2�v��DC��^�nC$ӁT���	�����~��2.!�t��b�=�^F�$m1 ���W��ԷWccݏ�I�~�,�FKs�%f���w:c���ކ��>6�9'Y�+2�f�,N9K��߇��>�G��,m�X�*ĥ
sW�M?+?y����x������U��ٳg�M�L�2��}g @��ͫ�����f�C[>�eY��H� �B)(5K��g(������7a�ȌQ�b��x���ܺ�4���sv�2 �
��l%/��1 C'�?����X�ŨѮ
I��_��sRMigd�@�c�HLq��+o���lx�������̂c��T�U�n�������;�[�����h�D]�5���nE�y9���ѐ�M�̸��|"�;��e�ݓ��o[�����hŜ�ƽF����٨5�Y�L�o��C$�~u=3��b�J��<>�o3�C��S �x6�<��|6� <v���za�`�V2(�>Χt����M�����/�s��o����_}��� $�Y���ٛ$�Br�Q���=?1^ ��DL��N��A�V~�r���>ޯm�౽�'a'˼ ��0���<c��̇5k9[[BY�p�v���'L��{eW�+[�Om��'�w߆�������>Q;u�s��(8�4d:}Xq�T��T�֖��c���=��Ч���k�<%�-m|֘��K{~χx��ͪ�� �O�{@$�Ky�^�7P��`B:G��p����A���E#ݝY֏-�m	��L�Q�[,]�%8%��� =f��I�?�2<E�M�F}����X*!8�V/��,7(�(���o8[@U�sD��b!��uS;����o��7o����=���G�U�! �Z��)S�'@�)p1�����ե��	��)!H��+��7ʸ��rj�p����I*��Z�*� 7����p ��T��O��/�E�U�����/�8�]D�h����0q�6+�7QZ�Q�
�J����T߶4\:c�|o�']+2N�k�㱐b'���'��^�Rv!�E<����j꫍�١g9�LyN�7yn?8ʏ|o4���������H$���):�h(��˴���)S��D�)�ħ+�)��Q�cP���3@yb7�A�l�=[�;�n9��{F����7<��<���#&@� P6{+�H	3�t���9�xD����D1�^p�Kq2���x`@O8Q!��J���crE�����M�r��XK�`��Mh��W!�/�P������ra'�M^�|9}����b�j���L�2���8 dS�B�"���[��E���0Gf�h��R�D�# �B��LR�\�R�N�Ȅ�gZ	 �e���G�*k$�~(,Ȃ"Vٍ¬�mN�� ׅ�&
	������#�CF�T��6R�<-����(��%�YB�2��V=/��
נ���=����2yѴ}�kf:
��-�25(��CSL�Ey����tB�5�(�z{�,�2==ʺn�LO�t&�F0��A�ю�f�X2�l f+� @���'���|���8���^�k����/��}D����0�f��IPq&g�<�#����;[�O<(�9Y+�2ũ�*M9�vZ��g�^����dʔ)Sڷ ���������fo���U5���ޅ�1��3Wa�1_�1V��g �IRZ���.�����R�$I�1{���{���ޘ(X
�Jy�9�p��sM���nq�&�ކ�9%)��������&V	�Pǆk��/�D(F���b����/
x�0
��p�A=�(8���|�Q���Y�'AO�^2�����Ly��$�:� �$��rܔ����Lc'����5/�L�2eʔ)S�	0A�UZS̾2��u%C��Ќ��\r�d}�#�!Ȼ ��)��1 ���e����+��;�':3q@~d�q�U�d���e���sŎ�9��X��Of)b8�P�P �R�Bt�����+�7��X����d>�N�c�\�*S�L�:D��w���������_�˿��\<�^\����XPR�I+���T���@�]�W�<G�G���19x)*Y`��P�(��K��%���}�0)0�JL��mTT��Opt�~��l-��%$=d(T�UI�3��a��nU�)��X�'z�5��f� �����$-�A��\�zةe��@s�2�rы���*iרk"�h��_V�Eh�1m�ڼ�+���xW������P}�2ٞ�����P�P�g��|��۷�}���޷�M��ל(�ަ�1��>m�N��Kǖ������x���ރ~-'��}H���}�-�����:�>>&��`�?��S�'��q�Op�:�W�I�1�~ϟ
�̿�����c���� 1U��Hvd������' ~`z}l
��@��1
����dl�a��6�1@�I��&�L@Lڳ� PIVq���H@�������X*��8�
�$���9���u�*r�L�IY��1��
����ږ����jV]=��?��w�S{�X,Lv Ȕ)�ګ � �N����?���3��7��_���~�x,�j��E-*�o�c���A�(F�� J�մ�U��]�m���h�X<xMi��r��2��E�I��v�>�����<�,�g1"�E%*D�o�0��%�-cGG���-�Ҕ�"�Rc^�T��� ����?����`�~6!CC�C�``X���6�w5�֏)�T4���:OjW4���6�R���|��X��Xi��9�|��|"c�}��vz���O�Twz���3�\�VȊ��S5n���S����ӎ��I�Gzz�U�?�0�G:�A��h�f�3��9��~�Ӿ�Nh�,�`Ɠ��ʔ)�p��sM�������oҬ��w5��־�$`��6���65��aJ.�F�.v_�� ��`��G,Be��ЈAp���ϩs1��P��r�!��\,8U*��\<
��A��L�R��$�
4F��\i��������������c�f�]]d�L�2��Cd �w��~�����������T��⻓��1C#p�)b�(l�'�&�&$# 1t���g[ �U��wH�"�fй�#��F�j�EҴ����$ ��Axaɂ0�� �;N����Q��Ӏ��Х ��mO��M�|�^;��)�
�2�U�pK�q���k�mK��e���֔jf���5�M�~>������<v�m���{��y�}j~ǲ�E]�c_kwW�vL�^��i��M�λʫ�׏�yt����Z��͗���=��3����8v�S_oCɯm�7�_���x���l4Z7��{�i�#��=g㇮�H}��}��E��b��unO�Ne>�
?5������B��9�m�{J����>m����(��0�b�7�!��S�k�_@j0���y�k ?�e��9� ;�3!�?u �v�_�$�7]"@����V�/j�T���3��� b>��Pvj��\I�<�@�R�`+��dMz�xM|�	 FWZ��N�9�������?���o�|����)�&; dʔi� ��i5�����g���gX��c�{���$zdUI�z�� 	�]�Ӫ������:*gi��,@�>Q T�n�aa`D�DP=���K���
��e8�t_�����3M���o��kp�&��*cs5��d�&P���c�\���t
�;J6^]%�o��5X~�Q���	=����Ck�[����������x���آ��g� S��V��ۗ�J�y�y������/�!�����Ɏ絏���w��U�a=����]��ljW�cן�A��6os��8�yRr�Ÿ6>����m�Mn���$�b���#��X1�>n�Wqs�a_�bG�=��|T�+��D���go;����͞�����{���#�����l�!���ƪ��1n7���A��^n���d���=�>��,n}�6u�xt�ޛ���o��6Kwl�_§�_���nrV<�����9ܔ�l�x톿�кK�>'uS�i[��3�>����y�vS���WM��3?Xz��X�v`�f�_;�[��qY��~l�2�.���͇��Z�tb�~l;D�҈�
�����s�u���g�D"&cT��D�g�:F'
�$���� ��@��r�lɊe�S�rZ){,��Q��7�����r%�Y���a�oo�����zngfVc�"3e�t�t��&s{{�+�W.�u�����w����/)!"�[�t�)�߆�R����q"ᵰ�&�k!y`��~G��-3���4�o��Rj~J�B���Q��l��3P��(���IH� �SeT;m��(�sjb�.4�6jcb-������$��/���d47�z�5�2eb�������W�LG��N3eʔ)�	�o��)S�L�2�e�A��Q����`)ПRtP�1�_1(���&��M	�P�zK��׀5��f��`��*�W�[���0.�R�A:E��RҒ���؈�p��ˆ�E���\ZUѕ@�7�ʨ���R��9a���]=�y�����~��O��ŵ3����fق�)S���W ��t~���_�����~�����-k	@\�j���Q:ې-� �_ ʁPh8��1�_)��G0; ����#c��*ѻK�sql�*�)��#ݣ���kО��טG�1;�G�O,�������t^��M��Sz΢j#M�� �� �ۆs�k)� ��ڕ���?%�x�Z胠C��m/����H�~��Ay����6����p��:S�'G�n5��My��XԵގ��4Ǵi�C�Q�?�M�8e�:8I�:kdИC�F�À)�e6��y�<���X���p�2}`�&�m��s��I���n���.n<f�1z��J���1��9��>�k�]A/ژ�:�R�?v��ώ|�����W�z�ʺ�����?��?��?��ޫ����̘���4�@�L�V�!2 �o~���_���#�/�����ۗ�2��y+�׫{�o�Eݩou:��c.2c�"�������u�	 �'ABhii������P�-�uA��.�����t���c�tz��#B���8���c�,��&?��l��M{�����7[���IۧC:>�,��⃾����&������i�,t3���Ӥ]#e���Hk�i�l�<�[�x�m��<���H-��X��f:9:��|u~������q�����3=~I�~O�mr���VϠc0���.o�a�l��s����=L�r�� �t�R�7&�M�#k�1�)@�RD��^�[	�TA��o)�� �k�'��R��l�9�p�e�IY%�4���:1T�$����q�>髪��j%X4�b�jY_31v��.~�+���/���O����_\__?֧.L�L�2uо �������~VV�/��ץ+�*WX�LR��1v��������#�c�r]Lc��|��7��w������t�;�:]��IjR���������z1, @�:�s�~`�"Y� �;#	���_�{L�Ӹ���:8�D�;=���� �D�1����Lj��8;|&j�rl9+=�ٍ̻|���S��7��*7~��ҟ�?�����Zcy�WRtXR�穏��ʯ��:��e��{�Ю`�h�c���3E#�	����sTc!���a?���~���g,qc��`=짷Lے�k���]_�"����&<&�כuЈ�D' �9���X�cT���J���+u�<E�;v�Q`9f��E�����*(#�Iĩ@�s�3 -ޗ���:K�0\Zlv���B�c+�52T���Ah�� I����g�%������P����n������\����̴�`Ȕ)S&Eq p��i��.��.k�9��y}���yv�J����e�K��@Я����=H���+c#�gf��S7����F��C�*p�!��ll�o[�[ ���Yb�|�Qђ!��\����Cy��e!�\& ʇpO0c^����+)y�دd|���\�O����5����]V�4�U�6�6�ή��	��v�=ܮ�fȝ����ǥ��cϖR=�Ce��w�e�Z���,Ӯ|w������.��tL9����h��d��˴Lc}f��	>�99�bl��[c�=%�&=��y�L��{~R�;�ǒ ��԰�f��p��Mt�Ǩ~I�T���`a@R"9d�Nc��3��ĉ!��ƨ_�܏�Ap"�%�+����0@���]A�d(K�VR�@��S�c��+Τ`#f�`
��7����Δ����?�����3�j����ُ���8�ۙ�4x_�'��fʔ�0�o ��_?�Φ�ҽw�tEAQ�Ɩ&��Gp92d������N�R��Z��7��ޘ{�̸0T�ǂP��At�%��B)^B�7���Œ$`<��!dL	���Ɂי���{�^Y��<,2�/����\f��p4r��D��H��h� ZD�D��؂����C@��,��C�=�4d6,��(�A
$%AR9 �!g�3s�ٗ���twU�+2"�R]�]}]�k�w���]���Y���_D$)(-�J8A� ��\���Q\�yc�(R�?Y�5�41h�s�:4��f\W��"1����.���;�r�Oks�����^w�K<J�<e�&�;��+���Z��M����%��En2���-	����m��l�㏭�}��������:��NYuf�v�	�@߻\������W��>i�*ݝj���j�v��\5Z-�m���ո�^����k��>�������=ߤ�zc�]��ۼ���]<A�k��~���n<�l�5�\ݯ����+�f�q���Z��jX/�~��}s�<�3O���5�w�������=�t}0ʩWշW�.���� %��7{|��P�yL�@$8�`e��lG��Z�a>F�(�B�[8`.�qx�5i�!�FŸ*֧��͞��-���Y����ѽy9������CUm�-��B �WdKl���H#g,�D�2豽8}�>��J%����k ���'ϧ��{��o}��*[w教�2�:s� ���_ͽv��|6�f~+ �;��Q���Θ�~w;窪 x��VV[�A�/����O�eϙ��w�!�(�ܓ��B0�I���Z�����Xo��$��(�l�b}�GZE��qX�t��Pc½�<�a���'R�����M�l})OE���G"q��\W�7|��p��P����ɮ���`cە�މ�!�e8����s�MK�52H.h��V��+���a�gv��{o�^a��[:�k)�'ٞ(]H�����Jj��{�+�1�����~t���e-���}^�H̏���������V�?}�x��;��??1�Wߝ>�v���x�V�Gm�������ء����Ĭ������Ͱ�q������a"��2�o��r���pr$��#�@ �ɕ���H�1'��\��� �ܑ�Z_��a �33U]��&lg����h�	A�P����t>�>``�0C8��=5c��/|����bZ��bˌ�����#@��佛������/��_�������N�����t|�ud�v��O;_��H ����D�!�X�I5"E$D=^W9��Ȏ�ð��4)<g�{��(_/L(ݿN�|����y��,�DY��k4�k��+g����?�����-�C��A��<��9'zq&6�ed<L���8f�G���ddddd< du�q(X�t��q_��v��GF�Q��2`�F���9+�sa�f�tW6!��Yڅّ�H��E\ΖB���_��x-fVh�I���Q�! ;o�kA8qfd��]���5�D&�H�| /V��v�X^��,"�������D�Q�� P~t;{��3o�O��Wu=����I�������ة � �a��x;����������?���Z����( �v���N�b���B�$T��%���B�}ⰹC�������u̖ê�c&���U}A���(QN��vV�r��*�Gpi��7�u������aO������fRd	��|#a'rO"�}itR�C�`PΩ�P>~���M8X
ϝ��}� �ʵ��B�Jz-tMDV�2O,3l�3c�ؒ`���ed��x��2�@W�]vr��]�l�~�s��k���8����WV2M�����Xy,s`���(��<������*�K���ҧ��p���a��<��I�w�[��&��<]�«�(R)��!��+�\3q�vΤs��Ĥ�
$�w�Ԟ�	��|��bt`!��$+�1�'�L����Q�U��OΤX��� ���݅�W��m?��3ӿ������b����w�# ddd,�>� @�~6,ԫ/~�/����œ��h8�E���[��^����X	P'���ʇ��N��Hu��В��E��r��[
�b#:N�d�[�����]�a��K]B�ؚ�X�����&]4��X  �qmhܥ����-'B��+q���%_�'&�S�_��?5�@�p����yQd��e�AaO�I��"�:��6�E�W/���g�[�(��5��挾��}�0���
��֯�C�Ьk�Cu��O��5�Mr���ʓh�X3�����6���w���W��c��mi3�[ĬE�&I���-0t��`i��n��m��gtݫ����d�{��Vl��+�hn";|�0�T@�kv�<���fa{�*ya#��΅�e�O�I���s����L�d���d�/���-ɔ�K�
�,�M�����j�((n�$[�KG�#���r�>F�ܶ|����7�����j=�]�}�.�ȡo�g�e�q�*U9��R7�����S��Ȃ�����$u�u�n��E}Ϫ�����	p4|;(�^��cx�ׯc:g�~.������v�x���r���I��#��n���W ����3T� 	9%�-q6�	�}��:ߗ��>�[6�N��F� 4�z�mșR���㱮N��[ox�6���/&����du���B�盆�cO��N?�����x5� �_�q����} T��w�^����f�q��*� ���z� �zQ���҉e$i�˯`���(�4d_��Ix���`MFJ)t���|x?�m,DYc �ҏ�ނQ�VbAF!hF7`9��M�^7�T�6�w��iżaD'�@*����G�B����V)^�i��TVk�_!9<l��7��>�}��1,9���6�m���b�q�cƵȏ���ֶc���j�1�>����h�U�!���0~��In���/zv���&nˣ#_���X�m��[z��a���E6����@������u[��y�yi�uߌE��{��Gk��=̺2�!"?��=���{�`��1�0ox`=y-��8In�!��λ?��@��q~V,�!��Q)����Q:k�*�L��x:O�s��;��˖�{�7i�F:-�9qFQ�ωx��F��N�dP�<_D��b\T��-�T��)\O�i���*���4S���=���x<��]������X�=�̨��l�E�[���;�]����>��$���
$�(��d���ߪV4x���ԑU[0C�)!��"��rM�����@��ʓ��I=lT�� �!�f��4��J9%s�J�M�@��	d�
��E�*:��PD�ԧ����9:�������m�k*�����#��ɴEr��2�=ƀ��9���P�Ɖ��1T��mng����,��s[��ɲ�C<W��y!3�儽?�������ʃ��3222*��ȸ�5��a=_э���0�j�n82"p^�Q!�0\?@ā I��.s(�О\���Bّ��/$���V�Y��"#GA���\K�<jx��ѥA�*N�'1���lP`\�'
��#�Uu������̊_�9�_��e9��P�����N�� ����;����������?�G_|�n/��
4�r�4��?��[�����3bE+B6��H��4k�|��֒B��*
S��[���z�wdI&!kt\��F ������
�,���$-nW�}�v�&�b�I�7�7�I�c#�P��#��Z�J��9�1�l;��M-P��F���b�V<�ot��>�t�F�|���ݝ?�i�C����!����m����tB�<]�����O8�CQ)ꓻѣ�+hv�Yბ���l]e!��������z���a%ZdZ����$!��S�E��׽T�b�!.g[όj|vׅm����<���2D��ߊAD�c�%F ����|Ôࣕ�9��m�������i�����=���+^�����t�,���{9.e����<}��G�vޙ|���ʮSo��{��k���]tn�)o��gE�G/���;�x��:�G�w�P�oo�����Mo*�����l���sͭ���GQ�8�v{������i��
(v\4��˱#"�W'� � �7q&�ƙx!��&�ƭ[o��5SQ�utÎ�q���b����J"(X��m�l�����
n��'�����/�����������C��J�	 ##��� �?�nN�ɯ�ڧ�S�Ae�3�*m�Rv���v����e�E���P�ya�C8�9H��C�({��~.�8|6��e�O�^�l�f� �ry|���r��;д������L�bAK�:� �u���
��Q���@�2%��z��N��L����	i'g5�2˰��W�fHu����j���p$+�G���*��W���y{ �\�̦��2n�_,��`�4_�f�<�:O�7eÂ:����褀b����W��^���:YMQ^L'�L��F�Ƨ��
I{/�d�m5�0�6�vpӱ:���-�@��sHrz(آLU����@���e�E����،6��8H��D�W	N�M+��-�DN��yg�ϋ8�D�V��c$�%Xf^,����7�}��x�F����1�qB �;��_2�rQ�G���qO�'�Ψ@.�C�i�0�2���QvW�r�>A��8A�/)����a'sn�R9����`���+��g������~�g/��~���2FPBFFFFvm ��c����wrus�n5��7Ss��^P�Y��O��5w�d5e}�H��J��Td�$�[�,$l�V�mo��V�Е���_2� �C��5�/�HQ�'�_�@�!�#��βB�8Tܖ�₣*�.-�*QP��Tچ�Ga�SG%��b��`�'bjz��7�Hz��A�D�q�  	��FG�����Ș��B?���[Ě�����dd<��<9��N,L�+�����m� �]���� N�
�0(�N��j8��П��SZ��.��m����#��&9{2��K��3��HQHͰ6��o땵��������BY�m���u[��n$��?�gC8������*�uUK�J�Ƞ��-�yw[���q�<h�q~9�����H�� opXQ��X����3� ��Â�F���P�y��� �=;~�<���1�Bl����/m{^�[~^�{~(�~���.���i�^�$����smс%³�K�9V�9�
����F_�E�_�x�GKN�E��	_/��!���(�*�%��Po}@	�R(g��66`gO�q�m�x"�i�ȃA�s����p��9��zrT���P+O+PϾ��_}��_���:�u��T�=�����8J�# ܕ���b8(�a����_���֝UC��=�n�^��0*�+=��I�5����Ç�}W 2���������.9:�Z���|�:"��F	ވ ˭�+"cQ;�Z��(:���9!TQ��6����!U�5������}Ԏ*���@��][������;5`|�`5���J�����{R� e��?�㕝���{x���v�����Ŭ��{~4�\���kg��$�#��������E_.��>Pj��`��D�rMH"O��~Q���o
w7�{T������C@�Y��|m��mQ�Uea6�p���WO]�7oJ��,��
.��a3y��%o��"��P�v�����h�H�?�`Y�I{���*�u-��Z�(7������T�P�h΂���;�4��i`Ln+x�����)�}=��0� ���|��w�<�0�Q$ K	�����x>����`�z�UZ׏]aY�c׼�H����y���-<n�Ŏ�����\�:�q����ܫ�D����4Gs�ʾ̭�u�"��=�`u�R��y'��*"Q0r���F��p�6�t}�OQ�D�����]��V���Y�T���?�U�`TqA!�pq�iH$zl����|aB�t�`��m? u���#�,ʪ����A��s�b#��s�D%�9�H6*SOe���<غ�ƃa1����:9Ɋ6##c9�b ���}�|�{T]Rܹ ���N��*g�Da�e�1lu}��3sQ ������й�5�����"�����A��ߟ�
��y1I�:[��3l0�1&�uw�B}���k�#=cD�E�*���5$���8t�(��3�&	��Hg�(��S��1C^��O�.Ms�Pk��56)��]�Έ~7P+߆<�M��}��!����AWn{��۔��&��#i��ȂX+�-ʷ�.$1��Il�ͫ^}k
/?�8�xr]�q��刈���4s��h�l�M�؜�����rF��o^���x��޼�:R{4�PN)����h��� ��2�ߗ�o��ұ��^W���^|xW��޾"Yǅ3�P����H�㢛��~o�hn��:�3�����^|s� p����?`$ 5�n�wr�\�bFh$�!k�8���P�q�פ3��#�򳒑�e`p��QT�"�����3ք�yc���a��(��"�s4pV�e��LwX.ӦF� F*�"��R��P�~+ ��x�:Me�!� 7,���{��p�aKi�eT0�c=W"�L'o֓'�>��)@�J�����	�*I�U5S��~׿a?��{e}� �d"##c��  ;!���{w����W~�_}�����3^I8}�6�W��NΑ�� ���áĝ~�-%rwk�Ta��V�tѢ���JH�T!��Z�fê:�#i)b�˕�ϨC�mp�P�iυ+{Y��*=��vV�z�Z�&xlK��#�(�K��>��ay'<_�N��9�ڃ�6�����9���}El��]�pg$h��mO�>q̆M� ?o�����/��:��m���`)�?6�Y�~�3p$��<�d
�|�D�\����" ���2G�s$���
FnQ+��Ũ=�+G�Wp��<�_�a�GS���AU�na��(�D��^��iš�V~U��ݦТ��I;Y�~=smД�`\�tH�;�_��\�!�D$���]���M��z��E	�>���'�a����v��h������N`���������}�w;isqj8��P�o���f���[���|d����#}~� �f�m�Ú0h��{���w1vf>��[#�px�Ot�|��8%ek�)�pE��U�B�x���I��¾v�q����������H�>T?�a7����\�u�ו��6�6`�[7˽��i�+�������q5��?��v0�TU5��W9�FF�"�#@u>8�������������W���5%n`K
ߑ�ܑj�F¢eB�i�T���4�l5i�x���@���A�Uu�,�.�H8AY���\�����Ңr�db�#�EY|�+O{����./������0 t��������k�9݊���n������e��?-u\+JO�{m�٢t+��/�Ɩ&�����_E���Ru�����ѐGȅ-��ƲR�%I���r�4�W�l+�jێ&����*��a�32[1�*Wm����AJw��r��J蕓M�Ug�����)w����]����'{��%����%���^��|��-\}2�G>Ӣz�W%y�c��љv!���v4�4�%ov��Ln�;���ˏ&��~����E��ĺtnR��k4.`8R�㝼?`�����˟Ig ��@�y����g.B�l������P�z���8�k��FY��C̫`��f�����#�?A���l�7��nK 	dD��
j�":&:��E�{fr��7�KW*�7�j��4ˉB��`����}�`�>c���ƵMvx���îӯ�<8<���ڶ�����sx����b��j�~M�{�)�#��zcƘ�����{�/ˣ���̧@��|s�y�[� 5��@%�8�q2�+��y�4G`�Q�'�Z��!�`��}���:���j� 6��F�ؘ�e�U_�"y��Jk���g��z���n?w�����'gw��
2222`� h��VY�wz6��O�ٿ��_��W�~�~�z�&��S�������C�	y"��WA�IX�p�t܁�a��Ml�x_{d�$,?���s0��p���s=yL��.5�_Eak�\�,�y�[QF���⛉�x ��OS(�Ԓ,��WMQ�PwPl� ���{P�2M�Yh�h�W4##cXB*dl��Z:���:7�����<Q�BĿ�\X��WSx�b�B�On*^H�z^c]������w�0����:��|�B��u����Vn��7�f���z��0��z�Ԗ��#�~9����uY���n��ζ�*aX��Q��*k��\$���Mf,+3#�p�����yφpzQԲ�0Pd��m�(��8#���%\�,�������mA��Ŭ�C�����b �O8���Hؤ������y
j��+#� �c��e�SGϥ;��I���\�\�"X�y>�vK+1���R	[�y��f6�X.�J��A�d�����Y��CU��2�З�p� �F�X�����lD�(�M�D9Y��"k%F��{�|����O\t��}['�[ ddd,�>" ��ӧ;�|tq��û�ٛ�ɠ�0��%Z|�� ���_:C���q�>�׋'~÷��ˤ��D׸X�t<��b�1�aY��#2:�
s!���E�T���� ���f�������ţ�:Z��@�&2A��E��c3�?���9��X^�!�[�E�
߁�mJ�+��H�~8��� `ج����j4��)#��c=c�]agr�:o�x(�j_��b7ޯ��������y��^�wץ#���_P��[��P�o�0�5�:t\������m<������[��5�:���q�I 'g�K��5n��2��=����p��<s�;k�����IN�y�OQ�3��d���NN��:yb��Z�C
��  ���Ljy�^c��mP_�ͩ�5�k�bX�����:F��fu�Fu�
��@��ه;_i��#z��B�!���Ͷβ>>����I��K�_lZ�}�!��:�w�����z��U��}�zU[}��D�Z�� �X�9ޠI�cDgYߧ�$�K�ё)L��i�%N���_c���@2�*��8���G��3R�#I�1��y�	$6j�	�D��r�S5�sJ1�#eQd�Y!8�R���q 
���a�`��l����򫢰���W��F��� h�H�|�[�ʪ��j��/,��/�~L���g=r*���� $|�X�Y� +,�1�Yq؈����T��T�v�z���D<�~��u+KvF,�,+Z���W|eU���"��Ph�k��7/���o�� �(lbm[�Iy6�.��,s�Ŧ"7j)�pā��C��C�ז�Q��"���Oخg��~��έZ����=?�ʯ�>7���հ-{�f>�^��{�FZ*��Y('�}V����T?$�]Xy�z�W7��
��)��qd��m	�[�dǽ�m��o�P ˜N�꿲N�����y�v4����<-��rӇZ�蕏� (�klw��;(��F���:�� D�)��Z�i�ZΆ�\�<]�b�� ��8Îih������@�����_&Y��轲>o�0���94*�ov����|���jВ�_��P]!V��+Beo�nߣb�[ݴ���Kɵ4��Ze��i�_��y�{:�����=G���<㞠�g�7�C$��h��t��Q�l) D�K���ȹ������H��ɸV{�"���»��F��Z���y�ކY��V �_b�Ih�xR6�р�L�9��Z��+��$�)G;Z�s�Z>/�oAE�cT��dddd,�^ �������'��W�����'o����_:}O�{�Z���@>#�E�N
��3
s�"E
In�ۯ;`E"�P���""���]5�ޥ@���)��Î�T�����*�[X^E��'+	$�E��:Ϫ��S���D�+�3'&�m��[����{��)�XV$�h���y����u���V�C#���')�`
��$�Q-�ddlQ?�gb�����+�΂��!?c���4�tW�V<-LqZ�F ���x��R �paIcI�����_���)���W��JPCF ���J20��c+��G����	$<��6(��MVh�1�剆��ͰM��Qx��d���h|���$J\�gE���ĸð�ˋ��}�|�{���l�q?�w�<��
�j�������A���5�ñG��ة�U~�32v��]����X�rP}�y/�� =8�?�z9j�q<����X��}o3p܆�h�1ͯ�lv�TP�18�K"'�`�1���<��8�߀D����t
�?�۳lĠ�k
r���i.c���ђ��-��O�!U1u�@h'�TU������'����IY��hl�����э� X����?���s��?���ߞΞ���g�RC
��$�
E���*ƈV�����ܗ�-x��'�y��+��ο*_��8�1^��a�x���,Y���8�[��R���l� ��*�@
�Ce�A��<(B�RGVi��%�z��K,�����-����h^�7T��Md*�m$[��R�Q�^�s�T�ˌ���5��b<�5��A~��gFơ�/@m��[�_��-��e������q���F��;gi�O�CQ�ɊȀ�A@��d������:#���'���2� `�Sǥ��ڀe-�ؓ<I��s�yh8��! �ddl���[�K6Ȱ�����u��cW
(��P�/?oG������ @GGg�s�9\>���|�G9�ؑç�ā"����ݿUpY��t!r7� @�\�BQ�0a�������k �����:�a���N����+0�e��&/�}��rR��b���5~k�a��;��ig������Ǔ������Ϟ�z5?{���/{@��eddl�� �_�w���_��:��Y��KUZ=��������D)�g��u���ǈ���*!]�<��N�/<I1\$�E!��\Ux�?68��g�b.uA��MG�B�h?���NԙuVb�@��_в��,��-���ʙ�-�� ���{��I�O����f��TF:��"����l�x<�9�l������R��{��f�������=im/�>ŢM��*�	�V/��ܪw۷�8��O=�7dS�J�n���� �����v�n���n֚���n$���}�T����Cm�і�G����e�G3����7|%c�"ٗ���5��{߄Vo��{���6*�1o���7��4����4,p����>@��(��Pĵ����%��xϗ�9�Q��6�֝-x�w��=�V7ܯZP��uݪؒ�z7Oo:��K�~<�-�5����p�+�#��V�����z���q_�۾���B ��;��iB�E2�F�� 0��Я�$W�����D�����f���S���ಅHgG�B��h%��g��y�c�6Č@�����ͧnDK��ɖ��k�oɕ�ZDa�3��4���`��t���?����K����_���>�O�BFFF��� �-�|���F�ﮞZm.maGh=�F���	j�F��-2�K�������Y,Ϥ�Lb�x�x ++:t�_P}\��aO�XF������|h{���ʈ���k#O|�赒�3����rŀ�eE��h�,(��Z/����I���RVHwS��9X(�A�������q�M�l=������ݿ��:,�{�Hv9���_7�f��W�~729(RyU�M��	����y@K1=���W��[�w���#7x�V�g��o����m�'ڛ�֮���%�X��iG�ǽ����^~y�|nY�O)���<Q��}m�
������m��%mX(�9��� ���
�hAӑ��f2�Xs��)�!W�яv�ۡ��;�^�aۻ���4�y����괩>?���ذ��V�S�:���%���;�ѡ=�'֮t8��Ϗ{|�	}�K�z`z�w�G}S��n]¼a=��+e=�@����5�Dۻ���S3��ȫ^�[�w�ʏ�W�c|�n������eYO�����-�%��jT��H������~#�!(t��)$Ễ��Q�:ؘ3a�S�����E���nT)s�}�]��ǐ�k�S������K�����d0���Qi�VE���&����"����vj]%��;a�C���dlEŞ �;i���~�V�r���WU�=a￳��ҙ����3�n��)��b\[o��V\���ѥr�{O�C̞���D�	�Xw,(�k ���):�OO�������O3M0��YE�y�~_�C��-��Zp�����׷�m8�\k�|�����x|��y��!�A?x��6�2������~B�t4�xmj���,�X濶|U4SB�o64;X�g-+"^���*��Z���9��t
��p(���V� �7s�-�[f�Pv����p��#E%��}u�6������scǦ�~~�������z�w�o�`�4�	��@AqTaH8��9�4�}b9�V`+�J�K�s)x��N��5͟"9��6��w|O*?Eu3x�td8 �?����(�݃�B��-�)!q=L����u�7�|0?"\I���x��g�B5 �ʪ�YQ�J|Ǘ�4P�퍐{͌���؇�}���V�}�3�?��'k�۸�b�^��Y��m�9�NS:�X���_��:I
�Ols�6�v^�drŝ�vW�{���������P�{�H�]_MF��V���� FC� �� D#pD<��J�{_сH�8�ؗ'�iX}Q���Qڦ5��Vvs�/r�O�o�D>0�E �WG[�m��J�o�h���>�����^u@�)���Yy��P�ލ��>W)6�z���)%F2z]��=վ�k�~f/5��x�>��O^�f��9�Z�u��EN�s��%��v�]V�ݿ�v�M�O��=���i�;�W�v��k���җ�����Ր84lT��</<T��(��V�7u9{���[��$�jwT(�\�y!=,��6-6�^s��8���]��5��'������`�7�8��ym��xqz�����xp��]�=���݌e��֭��Wʳ_n6��U������w���}��l�����\��]kz��ש���}�36��4��7�G|���@!�c���k�P��/�N�-x>C�Kx��n�&B�S;'Mv�$�ΐ�84�
�8���D���r��|�r��+�Zm��-��T$����[��H��-�U��Z&���z`�MU��
30'����|������6�@�eddd�b� ��z��r���}����׿�f4���TS�.N�a�-��lV�{˸���++�t�i=�-a�Eq�%���?+�H��1�҅v�?�����ؐ�~uݬu+4QJ�(�3'�4V0 �I�# o�敋�v�qG��J,(ݦ�N���ʹ!Ck�2��Ca���ӧ���Sq,�$�M��A w=+����x��}�f�坱l�/c��E�'눀��2�C���P�{T�H<������h ��G����8�پ���+�;8��=�W,���1��"7�9�71H� ��qM]%�q\-\���!T?�����JL���Q�FQ����\�NqTij �M�K/�?c&U��o�����5
O�I����}w�{�z����Yy��������K��aq����_����������_�������&�}ؖ� �2�̅`o7q�/V[bm%�>�s���k.QV FBt+�$Ao��B�(�?)3ԫ����Ȁ�r]@G��L8F"��*$!�$J���da��Q�r�0����)��Nd�0gl �C^����,���噑��܆ʛ�f�
y����H�[�m�f�w���ȸ?Ӝ9�S[���M�x� �����|�I/ �P1�1_y��0��	є=Z?:(��G/�l����\f�X��F�@D��9���?�J��h�)� ǜU*O���HѴe:���Ui�z=�]ڋ�����H��S8�B�fdd,�N ���"�rxc�����_�����7��'����QUw��]]>t�&'xg�/��O!Wb�v&ٽ�:u� �_\x�h��
�EÈ�ox���Ht^��/f�ԴS��C�y���Az]U�0�>9\��VȐ���0�W������o�p?�/�/����6���=jȈ�`�J`���W�b�#t�s������<��Y�[�ج*6��kH�����?��#�2����G6ydP-�XYie�h+�Ac��lF��;�و;�G����i�o�*���l�0�3�D�5�oO���ɖɪI�GiMU�h͞��b��>W�_�6�;���@��f��u@��˶Բ-���lI�2il�m�)?�;��ʒ!���,oGm�ټ{���'��_����`0��S� o����{� P���������z�?��)���%!E�c˩@���R$,J�O�rl=��S���=t���/�<w�x\��Xc��)Oq���]���t�v�l
�d�5��
Xg>�M���� ��q�kZ�Sx��3�0(���Zɩ|%��	���5�?�D�H*-���?jİONP�.�(�f�/�(:�D=���xc=#ʐ�;pd�l��l����?����3w�+����:h�7�~ի���w��Zc�U�8��Oh�����T�.�M��U�U���{���u_c���J���{���{�l�aw\�K���i�)�5�U2j���/q�zhȝ=��wD��e�iB�~Ū�h��g� '4jW�3/�D���$�~U��+�h�|�:��>��񗱚֒Y�c{������hp��%�9�&s��<w���[���ǚL�����n�j���J\�mڟUwf;/t>�;j����)�&��5�-0`��N���h���1��ɇτC�0�mCNu��=�m�=�5�[�'qC�\�@��e��^�GM�\�����m��Ch�����gNE�4�����l��#H
�>mT7K"��Qh�%c�<C����:+�!��JY_{�g��;���L�d6�a&�322�b ع���?�������L�mh�����	�8�?AsǝZ�	�+�D��y�FK� ^�R&�qa����A1�| o��� �	\]�:�Ix�qC�c�:Q�nl�f�
���;&������kD9����A1˧x��k^��/���X0�������!�)X�QYd,��S���8<���M���딷�y�x���C|Fs{d���/X���F>���bA3�F�~����p(��}�����K׽(�w��n��c�^��_�KFR�i���G��=��#���M�`���t!���,���:�����k���"���D�/�Ā��C$QF��X���u'�;b�f���r
���E{ۏ�=���X:h����O����C±���R��\�)�m���{�Q�p��nF�6L�+y�$_i�ƃX�I��\U8Z�8�<��sa��/� yϫP1�>BrTq3�c(�8�@�0c.�GU���uZ�%f	L���⺉4l�.�Y$�<�L<#����&��$�F c�n\\e0�]'���7�]9���bb�����؋�p8M�W���_�߿*�NKm�.P��CV:a�YjI�D3��F��aYb2�3
���ڥм��
$��
�F�'��S'�ea��Qd,�o���uآ@Qz↉v�9��S���`ń�:�$Z\�J�e��P�_%�ɧ��
�Z>�O��^3o���$��;�H��Q���_�{�|�յs�����*�.[�{�۞d����$O�m=���Kn�����[�y[GQ����������E�o%M�e֣����\��񞯊fQ����T���WzO}��3�]�f<�ݞ�o���tl����	c��
,q3���A�6dEAH&k��-U�ǀI����͕XD`��^X��꣨��31���_��Yg�	}���x.�%�q�t� 2��łóZd�IV��9�'���9�7>offi������s�\��ہ槪�D��{��l���J��V��V{Ř��a{����f9�.8Ԃ_ۻ�Cz���M�{�ϔ�����v������6��Vǋ��ջ����`.�G-<<6dh����*V����V)��{ޅcm�梸�j�b�q����齇}c�-���ݗ����Z`>�&Q�C?���=� ���c6��ۂY��Α�T�1�2'c!u�=�1z���i[�8C�O�@ADVP����)�xz�[�y$+|GpF�ۂ�E�mܫ��ef�N]�~�+_�������r|
��� K�S K����ޜ��_�;��g���_x3�<�YSh=T���a�]$ ��#/}� q���պ��뼋���z�1����=�5�ߨL �?���$�V��-*Y�Q�Ლ�(w�eC O�s�:����@�?�� Q�~�l+�򟱵��T�����-b�甤(dK�dd!(C)��!�&4��W���#��>���������6�[��N-��ӖjkCP�mTt5���	>����k��	Z����=?�rWC�v=��iBO!�<����~;�� e���?<y�x\){:6��qa���W�tW��X����߀��`�cy�zr;2h3�����F
��A�8�P�ᢨcx�a_�
Z��y�[�0���^
~�ТI	��[��ב�������`\����ᅟ^It1ު�j�Θ����0�;��:Z�W�s*�����ZЧ�g�C�<��c���c��[�Z�kZ�=�)l�k�Y�!=S�T�M��%v�~���ݰz��b;û�h���!Z�Dǋ~miw�.�V��_�����Z>ߎ� "�c.����i�2R�K��T(��1�������a�n,�@�U/��+����c�K��ɍ�s��C���[L�hݦ¥ �۞@�!XL�o���Q��r�|�[P�h��:�)�eݽK�\t��:�<k�s`U	��������}�����~��W�ѳg�f�g4��G ��ͫ�?�W����ޟ���*�&p��C�{��w�Z,� ׶�%�H{�eV^��4D�X�Q^�-Јr��qd��<�A,�X!)G�PX�*4��B����y⛉{EJ�Ճ�NQT ՝�"I��$1�M��-X�ճ\�E�'��L�_�-����YӉ��6׼H�\./�fdd�;�]dy���#2�(^~x�K�[G���1���q�&^+�����'I[C�Bd-̦�t�c�����ϱ�b��*��B��c��?�<�4Ӊq�EA��Y����w$��u��HS�w4��������K��+p�+7g��L�r ~M�1����wyʪ.��+0�qkG�['?��e�9Y�|�j����5G]�`|:p�P(�qm�	��6��eIP��'8������`H��E]�vs�P΀�{�ڵ���M4O�4��D�uV�Q!?���<�AuG��kFƾA�Ͽ�M�,���¹���yZ[����ki+e
����a�˥��i�4���Z_��>Y
���**�QAw\~��G"�)݂�""Y�(�E�89�F�_c�#u�d���ֆ�V�jR�L�Cu^=���K�~����_��?qZ����f����с] ���_��1���}V��'��6t�u'[
O��.�w����[��G�@���wM���<e��7ԁ:���鐵�D��a�����, ��}Y��[�*�`.T+*�� ���/Li�zMs���V�T��(���gZ?Zr���v�(q����|���?x�	`=�Pz ��x�%]���C��c�E�ށi���� t}�����/#㾡 ?�{ yy��U;�r��i zLT3�ٴ��d�]3� %����Mil?)��wS9b�;�~��좀�'8=+��:���Ut}=/���Ui�Q����\>�pz^����x���H`cY�O�p�d���)"�U��x�_q+Y(�-��v����$>�_p���"�y�L{��"����IY��60�;T�q���3'��Nj;� k��F��..����N.d��mp[9y��B�x|zW�[ö�<ǧ�C2,(͓����.����&��.wV?#�?C�m d�@m��34p��( ����32�F;�@~�簶H�T\}�Ϗ�b�5�Ր����Vd����� D$�������c���/�$�+p	!�q0�"�m7f�̯D���ӡ8^*�����X	��eduk�X�Q��$�A�r���E\�;e����x�D򈮱Y���
!�3EpN���9�^�R�k��H�r!�L���`:������w��O��G���N}���R�G���h�>" ���ksqvZ�f����)4ku~ޅt��[��@�ǋ&r,u⧙��Uc� ��>|���+QR����ڋ�
(8]ǝ8�K�����Z���.u���C�H�}�n&r� �鵥�+�c�.@�HE$���$| �Sb�	� ���u*Dm�ge'{l�v���X^=�\�Y�����vb��$ka�^�F��-�׽.j�>���b���}�?b�^��#�DG;�\�*|��VA��o��Kz���تշ�E�EG<����=Bg%l�/2��7��>]�)��_d�C�7r�t��=i����J[�N}��T�ƙ�_�s^�=��5���n� ���u5�p{]��-�;�Yڛ�I�Gٺ��J3p N/�n]8�=�(�|�|'�#xg\�)��8��Cb�3L�����A���C�5H>#����<�H 8%�y[��@��(T	P1���c� 4$8�@2�p��������ϻ:dqKy�����H�߼��檂�;�(Z���I��8��^P^hh�Fn�T��u$���7�����.�nN�<���n�4���ڕ�Ȱ �|,s�F����Y������������ј����g�m0�z��9ߏ��� �Uހ��������z�!���UO}>���T~}n{�{F}�?W���w�N�-�7���b3إ�ظ����]�w?�|=.���/��ӻ^�ۛ���>��rl���ɽ�S�C~�w�W����&R:~f�'@���5�Q4�#���"/s�����W���z�n���Ľ��G,�#��d<@ј9���L�s!̷�rU�G�&�B��8�sn�h�(��&�$ud<�Ԅƭh���X��a�ZX�|��R_��/Y˓�L�gdd,® �2?�C?6��o����~�����̠u7U	��;�h�� �r�ʈ:S���,$)&[)�#����,����Lұ�x�`�A<��#���]�"�B�{e�u�t�bB�Ч���A��P#YiJv��IV�}z��Wce7g�'�B:�3jo�|EA7��4�f��� �C;vŀ�cP���d�{�[F_Yor�c�ӄ�P�q�8��}�w;�?���?ֶ9�g5�
�*�������������Uo^����C��ފm@�I��)`ځ���))D&z��'�H��9��G"���[���1��]H4M{�;b�Hm�%Y=�(Gj��=�O�n��:������1J������E@򿮟1C�˕-*�^�-F �B֥𞤾7u\���b�o*��z ��OG�Π��
=������ cDmP��P�Se�����X�v����a��1E	��G���8�Nh^7>8Î�ˡ� 0��*�~S��fw����#�"\\b�{���z`�Gӧ�����>X����R��.7׭����!��Y��46�O��g{�j=a�|�3� o�x��g�Q=����b�A�=Z�c]��S^!���<�v�4�C��6�~�H��|�[0i/х���ȉ�|�ܶҖ=J�0�H���(6�yc�hPN\�8+c� �*��^�4mH����|S�E<�$�*v�c�8�V�5Sm~�g���s���h4�B�8o��� `���/��'�/�������^����@�uWV(�]Qh#SB�S�Jd{P,�=曫�uN�6)�@ģ`�,��pXT3:����9��6N[�i	�[�5�`E�k,F����Ҿ6�x���ӊ�������.�R���Ch��پ�x�2X�
k�Qm�R����#xY�Dͯ6�7������ns�Lc�o�u�0��5���Sx��n^W0�R�$@�	��H6#���8ud���}�O+G0#�;>/������8tE��*g��F�����nOyI���A/z��=�=�OΉ�GC ?O��vy�]��h�@ �"4I�����j���.g4�-Oi#�y'��$��H��G�c��h/�6���a��2����e.���ӡ#�O�N�(�����6�>�_͜����
F����._�^�v����:4��H.C-��x�" ��� ��6�H�h�!ӕ�6p 虙��&cn��3(�y�w��c��BE�Y��!_3222228º�F9U��Vg�O�(��K�	7a!�4"$���=��܁l�L�Dz���\��o8&[8�d������*ܣ��##6��RѬ3���7��������sa��|���La��A��yE@.�||R�ď�����z;�����/� ###cvj �!Hj�b2�����������_���~�|co���X8�(�zDz�ȋ����H����P���X�x�,�Ka͕e#b���M��,�g)�|P�8��:n��:~k5���V��*$l#��b͂�9�480�]��4�i�@����}�(<��u�HY�)��k��I�J�M�đpb���Y0x��$ �P��݂5��}Y���S�u_�vS���oy����C��w�L��@N����U�>n�W����^۽�[w������5[v���J,Ʈ�Vδ����{�q���h�H��	i�`�5<s+v%qD0�	��ґ�/�uWN�|S�� :NQx~��/\�v��
Gܻ( �=`\Z��j\$Bb����E@�魁��:�qĀ 0��:O4@/��'��|�8f�|q,�5�w}U�{]�dRB��3ֿ����� ��[8����\G������H�m>"����Pi;�} ���^}e?��a���k� 0M��`p� j�_������y䋱1�áv�}S�۫)��u�ꀡ�%�f1�������p!����-��'������N����멋 �F h(`hǀV9h6@��둟�:# �0���|����ˢ�y��Ȟ��>�T	�T���iž+���hB�~u�~=Vk�E������?�̘Ǯ3��h!�V�ZzԮ��j��ɚVx��w�)x��6��=�=���+Vo���d��_Do{�˰��_��iԩ�o���D_s<���,g��pi~��xO�(�r(#(��\9v�=�+O��F[p:Ks�� ��<����G)�z)�! ��G%
(�ڕo,3�J\h��Q���91p"2�>+�K?��D��Z�9==�� ##c	� &Ϟʹ���������_���Ѓ���t���9	/���׺,���`CX?�N�l!򝒪�rKB��ˌXa�d��=��9�� ��6"𢥒�#Vb�ɯ�"�C�+ '{�؃��:K���Q��&�#f�P �i: ��W'3C�BL˕:M�<W������8n��ձ!�6#��@�>\b=���&wH>���;���;GB��x�<�q�En����n����a�ygC89)��q1�@i\��[�60�7���|F��̋ ��e>�-`�d�ΟFDF������q]9�y��A����x[���$�v�����Oܾ�� �|t����ںae�:�/k	����	~��ۗ3x��^|8��ߜ��˙#ё�_\��6���ɪxF�02 H��G���ě��x
o_��kK�F
�E<Y �������n�W�XWo!`\>W/�u��?S��߂�5Z�Spz��e��n	�e��k�����˧��+�а�ae�zH�V2`�%�-�奨���!�_�C�F��W�5}㯏���3I�~%��h!�[��������@N�������!��B����o���QR��{�uu���Ha���r���M˔{���ޠBy��O���qĀX���f��䬘�_����4��_B6 ���X�� |�Q&�*o����5�C]U؝q�.�#�-�����j���BJ�bQ:�12��=�U8e�����
z���'������P,Ɨ@ľl@�q�|O��VN�E�o����I5�X��o+���1(��>�Y4�� �e���lG��jY��o��`�񬝯�(�8�Ԯ/�dl}���5����v�m��-t莣�_�>rE��󌌕��F�lŰ�8�Fr���r��?�«oM��'z	]$�u8�G��}S����t �)z�k�8��"̜�>�7�[��ϝ�x��hX@ǌ�_`���'��!�1� �b�Tp{=��]	7of�o6�ܢ��.����^"Ѭ����u�O�L��{N68p$�%��v � �yM�<���mn�6��U3t~KT�hN�E8�g'�$+4f�hH�OnK!����=�V� �9��6��+�(�\����!��
7����uY�i-o��Ǽ�}�^���@Dp˅�3�� F�8{��^P2�/��>�\�e<D���gdl��>��t�%�8�П�M��sT���p��~9��1@yZ���!@bd(\��@�!g�49kR$���Iј�휹��`�h���w�
YFG��8ZF�%B� ��$6&�L s8B@빭�F�*�3M�,#�< �j��S��B�g�O�����1S��FFF�� ��˗#(o�����?�/��[//�nc��t���: Xa	�/VRa�eT𮏈�XE�rL@+���4�J��|G�����4�@!����D8)�x�-@��_c�*Q�|=*���>8�Ѿ1���Dۨ>��~,��H���Ĳ�&�U�x~��x+Nkl}A�-D#�D����Z}j�wy�%�/�������N���fEi�'��p��y'V}^W�؜Y1�k��J�h^�M�v{�wZ�/�QH:��֯I����8<Ѣ�>����>�|���踶��)~Gr=��7�#�^���UI���#��e�X��_�nO0�?���#�����%$�p����M���[��
 !R��
�޸= ��hX0�Spw]�w�[	���=�+6H��R�u�ꑴ����I��C�OXqk���Ÿ6ү���b��E��`@]�q H��y�Q��6�K�Ww6�P�r���r�W�Tn0:!c��-��"%8�i&.���ŭ��p���=0
��EA��m�������d|���c-�BL��6ܼ�����'W��mPV<K�)��5Wݫv�����.d�s���,��e�Q^4��Jr�Ǳ�=��ońHJ����|�����R��p,z�m�1�Ϊ�gH�|{�XqM�v�K�=_��@E#J%�������O�h]>���ޖ>�ci��%tQ8n $h,<F�C��I|q ����be���=���y��d rf�o.2q�e7����V��:�'��x�����^��g�&Yw��G�?T��dR�;��'�BFD%����qة���MTY����[�����/��w�y:xg��tC�����	��IeOL��FŖ_���<[x�5�@�D��������)��%�X>�����#%�H]���v�\�������?mAP
gy&�d�@�bE�Au�N���J#�l���RҞ,�RÁ�A�i�S�����Ml��	��w�1��M��z�N���~�4�����ܺ�c�q��T�oV�8M�maك&c��P^ �:��3����\�V������6�Ǝ�um�?�rl��Wz�b���hj�[��������.�v� FcJYd�Bq��� �=���%���2�]F��SF#A�G�>��i���Z�1�sd[��86�#�+�GZ����]�����(-��-m}F��ֲEYw��������T˫f �{�
�.&��"�N��s���yF�1X�Ygޜy��=dɌo�_Ռ/܂Fk�(�w�qN�*Ս򊞣x�΅���?TP-Ǡ�N�{�t��uEb�?��2YS4{��$��B�����ϔ
Kk^�Q��`��>_!�֜�R�>�V)oY��vm��.�i�q���.:yO���!�O����&,�6��Nf�x����͏%��=���p��K^�y��4ȅh�hl��99�>g_�x��^�y�+��#?�1�#�<�����ݜ(�3�"ES���� �y�wvNM�"����Uo�P����Ks�hL�"����h=?)�ɬ6VM`:�������~y��N�x�2222` ����������^�&����'�j��lZ7
�.�+dC��4��L<����� <���gբ($@��"���F���jWuw����Y�(�i8L&�����T��'i�؇
�aF�i-�U��B��c�*�ff$�yo��e��g�K�o�QP|ʅ�QI�Z��J���^�5a;���1�1�a�Pg2���_��y6�
���Z3k�X#=�-���`�C��o��V�7Yw��"1�#R)!L���v�&���q?ɳئ���p���\p��u����>ДE4B�������c�'�Y6�au$oYL¡2z��F�y��^��CZ�f����g��#�/1l>z��^�n����#���4�7.J f�eb����j��;yw�rt�����t �u��'�����3��(�6��!�l��ٴpX&~&�W�w6�eax����=�˫��.
����G+���˶�1��u�r�����A��h^12FX�E�@(����ᴾlS�w�Ҹ	i��jJ�sXz�O�U}L;!ۈ�کnK����еAጰ�v�!Cl���m���"3��Z�Σt�ק
U@q����w^��(��[�Z�u0�s}	�6=�R��4+t��e[_DH���!�&Xԏ��5�r���P���Sc�jc�]�$�<�:kA���|e����AR�Xki�O���R���m�Ln���g�ʱ�Y��]�c����[F��/�q�i�}���?�
��˷#��L�����ܣ�>'m�N5<�!h����x��*�nS�j8��O��!��g�N�G��&N�(
_��C�q�o�1�1Y���B� &SL���ڦTݹt;k�pdM��R�;������n�j��������_����������2222`� �w�2�ڻ�Ϙ���L5;�w��cϝ�[��D�s�;����#ؤ3����/.�W�Y��C(}*G�Ϝ�=H���bc%���n��2_�n딖����=r���ǲJ[m �Ė���1ߋ�'�e����R$��H���S�x@�0t�YJ�\��?�J�6�-W����x\�].�����G���{_z�3�=�m�m�#}rY>{�����?��Ug���j���j�S�a"^�\�1P�t!,�&/��v�w��U%��u�ؠ};/�I��Tg����F�|$
m�ǲ;{x仞�n�g��)�����YiUz]��ע�
����q�B�&�y�9���w��e.���[(�j8����c�N�S��ho^�����*C(�x�#��h<�{��ɳ�ۻ}0֎(~�j�!Ö\H�_�eN�0�=�-F�� ,��@`|6p�.�</��m�r��o�gLt☘�eӺy�c='wu��I��8|0�m
���O�óO�����p^��������n�mN��V���~9��ƅ�w�*x[���c����@Q�$�E]�'�G�O����B񿞖n����&���!�Ǳs�-|�6�y �y>��Q�Y��2�C4xa9�D}M]?<��\I�����V�o&on���C4 Qp�d�����cx��x��N��P�͉ۖ���,����8��Io�����L�nD�nN��6�N��-/�.�G*;���_��2u��_E�|�D��5ӔK�g��V"��׊�d̺���b]��Y��ww����)9H곔VpCְi'�����1W@ ]ڱ��\�f�e���퓤7����А���,�m�o�%�>�����q�[m�]��.ڧ��1�m�#BW�&������T8v�T��"F�=����i���0�1�)<B!����O��0o�P�$��CDbB,�(��DX�����`��Gbn:\�S�8�6�lK-"���xP��Ve	��Sո�����_~��_<�^���TW�ʌ��G��G ����w>~�����z�T���-ޠ��G��x�=x؅N=&�	m=Iw�fE���Z�^,���-�p�D��j�� �{�Xg�f�����5�d;Bxk ���x��B��F�[+���C�\D����r��s�|.�{{��8�������y�m,�������	�G���dd�	܍�v*�Wt���o^ͭ�e����L&]��V��C�E�\�����p��q�W�V�I�!��H���KG��fS�:i��2&��4r����w�#qql�<�"�q�x���d	���i�Og ���9�c��k��ǽ�K7��w7����%���SN�S\�7{�H���Gu�����pz���ǐ�H"��\ޘƘ!��X�0�|gDT�dmL>�H�?}g�|0�����#w?(�{@������	��vHp��r�2�e������EQp[4��m ���@�9��CE ������ 	?�\ZQ��j�FP$��X���(j�!\��@r�q{�2�v�y#����h������z`��Yj��������������x/�3d ��Mm���o�@���dk��F��r�VHu[�3kS���[�z�zC-�o80� l��{�n�A��b`�m����/��cV#�.���3/�dddd�#��4�Z���@�� ��ȋ?�ƣ"�]�M��R�u6�:��t���tǥ��j4	$#j�<�e��`� ����\>6�D��ˇ9�F�Cĵ�ܲ�� ܋|o�f!�u�����leݜ	�3Lt;��e5��O���dprrrH
?##� ��- ��Օy6>/?����0��{W���MT*�:�`=�{�:@����\d�hq�q�1aNdƆ=h¤3&�5/��7���ó�?��
��>�����L����G��/��E:.�F�G��f�)�_��)(6H��i*۠ă�^P�A�7R��	(�K�|:�0&T��$���5�\g��(�ma���>�ZT^2r{d�aA�$���^�	ol�����q�^s�+��|��"���4�P����½��gx����
%��C�zsԼeޏm�m$��!�ZW��+�a9ʄ�)GQ
���;{vX"D�s�C�ӳ��,�x�3)އE���&�([S�HގN�#�ѓC��9��G���%G&��?�ރ��H`#��d6���nLoK�~3s��q���� #�C�?}>t��ϟV��v$1G�DRCٟ?��x=��Hf���\ ��u����z����z�"����R�U���t�ל;��!��3@C���I��6�?�'������E�l�DGOz4��{@�{�Kb8 �F[p�BC�s�3ܼ5p�v�� 1������0$汽.YV�7��0�Ͻ�'h�0tP8O������v��.ߥ� #18��!y�]W��bX�����i�`$�����ӣ:��3���t�[����m�k����b�Lt��u�ݩ�S���#\<�EO�诉M������y�����2��ߢ1��8Y����x�`x��p�s8��:�m�������[��k���Z�[l�^[��`��*��
����*�c�oZ�}�;
���n�vp�x(m��6d$���si.
4�U��E�w����H������eE}�$	��agA�1��=�Ys:x�V(J�t����rEO$�uyƼS�,8YF��A1r��5-qT9[��a��,_I�[�ι��<bjUQOnF�B��������"##c�ص �v�O}���~��������7��zv�mz<�eU�Շ������4�:*�TCh
�B�چ	X��%c�Y:e�=�)o�4b������S�N���XA�+H\7�5+!��׹�5>��I�(���|?�_�++�.�$���i��K���x �"X���$�џ�����< ��!PT���$c��F�/�Z��
+=0?�hҢ��9���m��֯���L/�-�m���d7J��:��䮎Ms�bͺ_􀍆���{���k�k"���
����4A��LK&�pBa�+�&`bn|F���1�hgCX5�<V�W({��?{��+Ͷ��9��{��~�}�>�>�b�(��@��(
@Rx@�	��H�H<�����`d@�H!$��';�����s��n�ڗ���o\�U}Y}�^߮�wݫ�j֬1g�����Ĵ�610o:]N=�?��DK � � ��3�m�aߏqy�i_$�sY�z�fR�Cа�ULO�/Ƽ� P�A�Y�,�j���(��sm�/BP ؈B���1��)T5��"���z�9��0���9��U^��{v, C��`o��x��mZ?�S3���Y�ٺ�PD����2��
s��0�S�x7��J�	Q�/�. '�T�8�@mV���Q�P��Ci���� �	�G���Q0 p����/�������vĬ �@���A�!�d�{�>�.�P���Ʉ^��p�Gy�rfa ��t�S
�v�È��x������7�P�����t��B�^�쇃��n8��Q�tix<3���h\|�+ȡ�㻱y��(�pv�n[8T�;Է Ʈbq��!��ū�C�/{�W�t�{����Y�ڕ�x~41!�:] D
��#��K��v�E����%��%uΘ�#ݱn��m29*�*c3�@F���m��9m|x�s揳��u��U�f��@̑ɬ�莴f�+�a��܆�HX2�%P3��Z��N�<;	�(K<�����GOc�D�P��aX��� �B��q�HD���0G�u��1�/�}�X��αǢ�����S{hri�o\��.�"~~�_�u՝_m�~�>Vkʹ�U���Y��jN]��4�p�>��RV9��zLɁ�����!�Ȃ��#��FK�`#QT�+�㫶�zA��T�U�4(�Ϊ|R� ��V��UG� �3�2�,��C�`T���lwޘ�:��?�dEV]�'��������c��FPkG��I'�,�C0 ���ÿ�+��~�w��������;�2�^��*�#�| `����,<)���z�K(W�D��)MhY8o���&#q����M��2��.EUƉ�(���G��c=�M��9bl���p�x�����O�;����"q�X ���M��^`����J��}��r�������@��y�����邏N�.�}0F�`R�5��ޟ�� #JfK��7ޜכ��Yn%�%�=�'������UC`+P
3�\�&�	���tva��uF����`qB�{�j��7�G��������z�\wGD�Q�~]8sq��#"!������@�X\���u�Js����8�	�CT_������؁��u5�D��N�������؉4�9*��t�#`^�����,0� <�{����'���'�I��e�G���A^��| �os��i	�&@Q�uY�>������pZ�0 � �@��s�Yo���H�:�`���}�:J�C�N�t�T }fxhK`z��O������Fy�ݲ�;XWп��0�/��1�y�&`�r�F"s���'�z(�X>E���ɒ��Yz�����m�o�u�(�]�#06 ��c)t6JQ_L�5����VCN� ����> ����Ҟ�������
�����\06O��8�����Nc�+8f��wyrLsc{���0nи��>�!��� �-�����5��9���f�q˳����	� �X�>=�:��6+b8�e9ga�����?��s�Gav�Uێ2Ov�W�g[u�y:D����`Y�G~��c�*�1��rɎU���B��{Svv���Tt��O�"9�{�6�.�`_���t;ٍ�A�t�ah���ۛ؋��0�x�Kk �Q���]��
��!�!J�(�靭�T¦A�ρ��0�s��XM#�1ٜ*�"5��E�o�Z�R�f6�r��{�� �J��E�G�H��qO��ԓ������u��?�瞾�|}�[�i2�<Ͱ0�t�I'Kd� �@��V���\������������P��Շ��e6��yL(���g<?�G����k��0��6�@~,/8�EoZeh��814vz��NtDMcuJ&;'H����G�ܧ͐��y��;)�����K�D�x߫�����l9Q�zoq�_l�e���ߢ+�N��oﳹ�}Vr����N�,�7Y�����r�����9J�7l��V�����c�8'5Y��>O(��Ef�r3#*4'�d|`�Q�C�u���z�(�H[��>M�݇�y�-��]i�#�R;�Q��MØJ�Zn�F�)^U���9�^���ޛ���]�L��5��0���y��$@��ۂ"&��.�u�#$��髲~F���0�*,��}d��$-�' � D����|�zB����~��җY=�玞���^��fx�	�u@�C�:�y���$�]3N�s!�'u�u��cC@O'��DN��~�	�+��̰!��}N�r8�6NLqMYu;=��ND�	���3��
rL X��!�3�pG��``�ze��q������r���s��Fu���1��z#ݙF���bJjo���U̾��>D�����Kk��B�����/��r�ܘʾzգ����}#�'��Ls�)}������� ���+�?G��q��U�%�i-�A�bA;�ű�5�C��#��c[��>��__O��cud	:ޘ�,GV��~��u[U�52b��=�6:JA�퀝��lr{�@vb��Z�Z���)�Ub��T7�����6~��*rS]r:
r����Zm�5+�9�Qi��q�Lw��[O�)��Q,&��<���|0��s�q�d�P�;F���3��e�ǂ^Xsa? G�c>�4o�f�:��:#b^����c5Mg��{Ar���ne[��礋S�N�;��'����3Z�ǉ�1o )V�# ;���~� |���kT�w��z��Փ�"B�{�B�ͷ����bψ��@�?G�DZn�nl��T����&�̯�=��-�S��\�����PM��/�S��z�����Ks918;餓NT� `���}�����7���Q���ͬ+H�X��-�wE��M;�=��øS��<�w*Ov�:X��S�6�Lj�2�*m�����gZ۳L���{i�O,��y���Ѧ_z��Nѹ���G��o�=�)�L�[M'w�lMp(H�J��u�Ε�[��X�v�p]Y(lD�h��3�¿��վ�+i��ov;���i�Q�	x�^X��$��m~�bQt��3����|�fj�������C���'� ��"3�9�B����onL�/$�71�}����c��!GQ1�t�~j��dl>~=6w�
�*yj�. a�G���]fFoY�J� K��C�N���	C��z)��#�wk=B��<�# ��N`�J��-���z����p��S�f�v�G�l���D��zB�݇�L�׸~~l:��HC����Ӏ���79EDp��B�V�H�TǺ��<��0�[�q�$���L��Q���=z����
�31u����J/)��f0̀M`6�5�zA�5N~�4ʕ�	�ԁqY��t��hS1c�0 �E��V�aLc��!���w���M�� <v�p������޸7�� MG�� -�4֣�"�i�6�j=��켠��?�gL���v�E(}KQk �
�m0���:f!
9���3Ǆ�Λ^��V"��>��3����#ܲ!�W��`dz�ⶕ��@�eoH�D�����2ƒ�p �8 G_#H}�~�=f����z�3W�sJ��q;��6�sm���nŚ��CQ��u?y��������wr�J���������#�^Lk^��W=r�)�����k�~T�����8Z����0�������OA�=r ��ZX����暫�7�y���L	jO�u��؂�0va�:��t��B����?��JQ�S�-Y�w`�zz��t�����%�R2g��W�����.��QU�Vv��\t'�>/I!m���`ž��5:�լ�����c�h�f:�ٲ�N���L��f`����5��.D�k�z�-��ꠈQ�!xLU��R�����`[LÂ҃5@�ne1t�81�����N6SIk�g�,��8�i�11������>��}]��YV=Շ�";餓g�  ��<����w~�w�?L�z���r�_�Y0��!K`��"�#�yh02xⷢ(eR0F'�F���3�R)C���$����۠bI"�}z\U�9��D��1�k,�̆|�L`
�Z�F���8��'�(f��~�O<����(l�m���sh���5�!R����{��f���ea�KO���\�N�Ju?���\�U������B�c�9tE�x��a+����������7?�O�'6� X��(���x��;5��Ǝ���� ��:��=�K��v�g��h4D��fb����y��$�~:e��c둌�d����<Xw��F��
 ��H���*@b�/RT��PG��Gl��(I��6GPJ#R�	�wR�'.lF���?�a�:i)d}0�)ʔ�:�$���O��4 �8�M��G�H�sU9�>Ay�{Y�j��k�RpYf��7�!&i��1M>�H��.)m�t̹�˲	��2��}<�A?g��>S�;�W|�@�y�K�[���°����N�2���F)�jGE*�|^�i�J#�5^���*'_��=��Gx�B�QLc�9�h�[iWXW�Oz=�PJ;<���43;p���9��!m�:LSt����<3���ځ�J;��s���W��6H�Z�=�Da��{��Q�P�N�]��m?3p�c��S�@i���q��M�n'��8&���$�|�6�ܧ)ZR .���z�[�pQ���~}}�lp�x��cZ'||7&'Af�8��.�"���/�hD�c����=� N�Z�Y��"uXm��w?Q�bR�T4�#Oq�r*D�c�
6�q���S��B���絍��H��JN��x75�����)�IpTrJ�c��:cŸ ��xV)���ܸ�5�8��&��.r$��~1G6�g^V�!Ơ���U���(~���\�V�.�Z��b�뤅�ֿ��;7/JV��nk]��l�YSH��گ��	s��ā���eZ��o����&n��U爘�`)�%��j9xn�dm�b>��ȍŨp+��g;�HW��!���u6��	:����]KqƅtO+����da��w���༺x�jR�;�I}�����t��i�A z�^�����7~������1�E���b4{t���P�1:X�8ӱ�g`������q��q��yB=��7����o����C� �w4�0%���x�	 ���682D���t�� ~�������T�\�4ʿjM�m�8I�u�T<^'�y�����ؑ�/uHH�pfc��v���.���}�����w���&��t}au@v�o���4����φ�O�ǔ�ߟ�A��z�d%���{���W�J�M��b4{���R ���>�FT��o&D��Q���K2J�-9O�Rr�;`m��� ����V������n��dJ�PTBG����_O� �~��O� �
�fG��o.��D`��+�Q�ϱ�i��x�D#�z�3�>ty'�=y~"�W�۟r��BI�rj �B7�]{)���о��o'�2nj% �/P4x�� �`�i�c  }�s��X+J�<`��KD;6Ӊ�U$�H���Lz���i�Eϗ��>��t�'3m3�� �

f?���XN�V�CH �	�;;L��㽚3撮���Q�t�����r��f��b�"�}�u������̕-�p�rMf	߬+��8a_��ǃH��} 
�o9����P���=;�{^S�g6籤�"�q���e^�{�'���^���M�c���hLF�z��ycuU����s��~�9k�Q�
瓨���G�Z�KKaDA*��Z��h���5�H�_yk-8R����H��i0�uk������T�8��u��((���,
��-M��
��У��8����)8����3r���LO���
ײ_����mi_s�	�cF^Fېc�s�k�����k���d39�=��Q]6}o313�N��@������HЦ/¾�걶�!#hN�;UE�����śU� ��3���x��*4�߇ό�X���� �C�[�A[6uHOX_�*��{��I!��[��)}f>M̏���\�-�1��)줓N���: x�主�8�������l���rz�z
��h�#]��Jw�<�{�x�#�Q��5�gv�5�6��$�o��������Ury���:�7M6Mh�iE5�	eП�l2s���s���9̆{TP�4Z�6k���]~n�A��8��߳��y���@�	w�� ���f��x�ω�_h�}�6��֯NC�|0c`����c[m�&K,?+mܞo��({���gd����v#��uU�(��OXk�u19�g����4ga�.��-1������=�,2��i���N�O�9��I�}���iJ���@�mNFh�hC�Yz��yiz}1�Z����뀁k�� �Q�P�2@��O���P��G��(�?���� S+����(�F�Lr��dq���>�?��-^2@	�x<�m���!w��8Q��gz�j=�����O�8�:�+zaf$;���/Ď���]�)G@��ĕ�s���8@�o#����|�eo^nA�R�V�5*��9Oo2~� �2��䵫ig�b��� PJ ����`G���K��p*A��c�Y����B�xq�V&i�vA����P�,�ym�pͤc�-4���q�0⬑}���m�x�x[4�V�ǧ7���y��eS�Ӯ^����Ҕ�z<9�ċ�����rI;��׋��vX5M����'���!"�ǤSe�8%!�/�d�?���	y=FW��lU�2����v����ʈG��z��48>ݕ�<�Z��V���g��.�z�'��tJ#MƎ���h���a[����BI�?h���4`��BXNA�-9֕�������UQ�Ysv��>��a֪Mm�gG�ӂw��t�\�fm���h���Z��I/W�[ɦ��*e�����Ӳh@�^�3�m�U����~?�#4���.�m�;B���wK3�uV%����:�_�d�H1�褐~�X���o�əC���Ȅ�k?+�^7W�9��4�8OS�ͧ\�x��>��9�{	l�q!��0*��z�����+�����_�������e�i-D;餓��}3 `���o���o������M~�Ӯ��\U�̗6��WJ�����D��1�����8:C�ql�	Ax�Tɠ�:zM/@u
��Q��N3���^� 1�8��)%�2hy!�?�)b�tq20�i7ћJ%קz7"��g�z�͖�+uh^o�Aˎ�)�Np_h���@'�r��n�NA���E=�	��
:Tl���>eG3��8~J�:c
E=s'���:����# �D����IQ��?9j}��0eLG��9_	�qM���ν�: �g�C}�i)&O �$Z�8M=VB�c�n�����=q�:Ϛgi0���ωh1{L�=B��{G5Y��0�źb��h�k���B��.�����ҾD)�Y?���;ܮm���z�[1ϐj T���_;�H��iy�K���/�A`�>��)XK��g�A�����T51�1���Atq%N!3�6z�Vq�c�G�)e:�R�8����:!���}��8�a��,�5�#x᳤V=I)�X"iF=\��E��'����2��J��,�mpĂ3 Rz�Z$�	�0�<Q�Kj�CFثMC�$<+�NG$�q�����x�`h-��6�zk���2�F�����	,AԶS8��}�D��-�Oϩ�Ѵ�˒S���ȶb��N:餓}KL�q��[����.��~���_����6-�<E�2�Z��.�)8X4�/3���v�W,2O��w}�O�&%9ث��a�\���������℥1YG�T��s���2Yѣ5Gu6��ɗ������e��W��??����W%�D��:餓S�C� pv��M��(muY/��jR�Vz��]���\�k�>6RD�(����	՜d�w�� �E��ߓ�*�AOd�H�}H'��S�z�5��Dc.H�4U�� ��0�ʥ	Mӻ���S��IL�KF�㿵 �s��y̓�� 8����q^Rƅ��:���1=@<щ0YPȄl�7O�<O������d�{[�_U/��)��s���}j��9?��nfB�Z�y�A�m(�y:��e
��X�i͹|3ze��(쭋���ٓw*��F�`��}��L��
����Ҭ���AIK�������N�P�x��� �o�u}z�r� J@�?�ᅜi�������ԁ�v��qa�zI�4G.�+���5beOϙ���Z�ó���	J[������aj���4�z_�� 2�&��d66�(���l�����k������v������im
��1(q�w�a�nm�%�"4��>`g�ʓt�K:";6Hz�z�7��sJk�5��c��E��Iاh}�u��Y��,���Xs���	'�F�N4�d�>p̈��*{
C���:�����g(R�sk	���hm(�m����1�/�٭(����$��Ef#(�R���b���8��1�7+;��'r[Kc�l^�l�>�'�b��z��餓!1 ��yi�mp��M��\=��~�R��ߵh�^����Y�W	&��1�Ȋ"�[kx)3F����$)�t'mց��ƻ��N�54���$kl�ehT�Q�a�V0ʦ\�ʓ�U�F�Q}�	b�
sI�D.�};\\]䃋a�����I'�t2W�� ��ȍ�����z���$Py8'eb������xu�&Q�E� Ol� ڜ�b>���y�|�h�D�d�D����A9��'�b�)��F#y�y6�Ǩ/'�3r��P1�� m�1A�*�$*�l�ǙL����N�l�n��`'������3�I���sL��o<>��:i��������r�F��-;BP:Y]ھ@���$N�
@ ���Й���X/8�
�}����`���?r�^�7}s��g�/33��?gt,��t�{�%*�Tֳfp^��:�u����̌3��SGē0�[�����e]�˺�W���8t�;�RB�U��u� ]'�^����ú���m�RS������8Z�������=���+퓽Z�=�f�S�:�I��.k'U��}��"�۷g�^�)���-�1��I�ٖ۝�&��m�:77_��۾9�u�~J��ɚ��O<
���!:N�k�\�z��h �sD�qR��Z�W�@��I�!�eY�ũ �v�9qh&v4�r�񑆞k�xƴ���d��z!g�D�
�Zq�~n�wV�g0����׵.�0�.�x �·�T�c�*>����x�P}��8�����݊�%b;�m�u9����D�-��^r�O�I��}AS�`M�ꋁy��Ά��ڶ��{Z�;ۣ��}��B�r�`�)�5���f_1ED��|�GA��k=0&�z�~ݧ����i������m��Q�d��y�������z�u���s����k�� ��#��K�����L�/)H,,;{4�$�d�vĚo,�Qz�^}����Z�H]U���#�O<�x~@�O���5k�LmaS󾳩�$9!g�N:�d=Im�q�fĺ��ǥ�)�@�G����8h([Ăcނ�( ^ ?��R�_1��Z�o{��Ɔ�����6#�s���!�e��r�/�(Ӛ�1I fZa<@��u�&����|�V�<P9W������(7���!=����;餓��o ���}��ݿ����_?}3z�xW���\hu �&�K��Lu6'�4r�q����f�#�j�br1�ߙ�.૪��z^�8�������+����	!�	(&1�8@�$�2
$s�N�ޫ�C���	C�@4@���^�kMs��z�n�i��)�+��Q����E�$��ٶ�Izc�On�ٶp�k������ml_�U�;Ku�|��K2/G��������^�s�Vy�;��UZ�5����I�b?��U��	���UfʲGFj��@�y�9���E_[��^F��͛�y���y����倌�0k�0���6�r�ٻ'5����uO��3��t��jI��˲::E-��4�@�+����g���ȹz���Z�XߚG ��/ ���� %豘����h5P:�GV"�R�(`�G�C����߭u�E��)���8���Z����U�Wq����#�&_�k�[���!EX��c�$ \_�z���3�՟8����M��}Jg,t��~�H`p�ym��u����Cd�|�^Ak��}it?S	t�4Z4lI��Ӭ��	��"��iάк�wAc|-�'p=}�Џ�M�*}�����=�D
1|Q�zf���%IWh#� �#������\/�{�c�/[��Z�ޘbN�����|�K��r���6ŉ�3KUB߲�YN9��(��^7d���&�:s����3uig�����W���ﯾ�7C8�"[P�M�=A�ֵ��s.6��X˪�]�W�c2�8v�aõ�g��*�����8S�!�
z�r@:��eǬEc�6k.���S�)kV��5h���
)(��l�����'��Ê���'���M�n����/��V�~]�e�5X��cK���o���I}D����ZC�䒚���E
$<�)SL�q�	�d��)����R��z^���z]��9�@klK���M���x���s��,��j�>��e����,T�*5�'�R@���h̓*ue��v���)�2��n\X�����9����fm����6۱^�����4�oJ�O�˽�����ڄ@p�A�Z�97��/��zXZ���������*��dO���2;��z�	��$j?���eYK/�a�{��~�lh�S��&�&�������t������I'�,��; ԯ����Ϗ���������g��*;--�������V2?wz��2��9��x[��UdC�w��qR��]� �M��b�[��e�T�&���ƈg��a��~I;����V�~S�w��P7͉c�z��1-AJ7��$ߌ�O'��MS�ϼ0D�V2u��@�C�ϮCN8QT�b`��9�F6^쯴�6f�RVYܭz�E��5�=�����}PV��t�����t�����u��g�������,2���ݗ�K�L2��	�u'��⊣� Z�&�0'�50���R�q~���&8K@��0��>��]z2\>�s��br$t$,/�C�9aDU����Q��t�2ʔ��;��t�R7�l�?;w�|���$7E�76�՞Q>��HY��[��lp�x�U߼�	�i�K�j+Plų��1 ��;@�sCu�QN�N(�{g��'#����WlV�Pf�`@ ���2Є��-�,����;��(s�sU��7l�ƭp����DYq�g������3G�J� ����}���ᅧq��;ʟ�X�g��g�Tn}�T<�(Ҵ�Q� I8�z!2���zB��/H����+d�J�����PA�B����g[�W<�h�����|���`EW9�)�cL�H:�x�41�h%���\n��qt�s��"���
�y��K,:�SM��o�A��D���,tb؛��('f�3Gso��	�`6@�Dnx�^��{�s5�d��z�����`P�w�9�����FŨ�.\�a˾�N ��[f 0���_NYa�3��
�ȿ~�������-+������N¤��~�M0�;y~�����z�U}�8,�i�R�q�*� /���J�[WX�^���h$��d�Ye3�J�p;an����Z_}�%;O�y�Z��t8�ڵ�֒9�B�:���O��H�k-#N�۱(���#ɮp�Ue�f;�s�D�ݶrL�ž�բr��!v���ުXO�q�Ik�O1�i��<6������E*F�aW1"�b!�^����Zv�t�H���.�1�}��#��: ��8�&'u�s�W���z��iz ��EQ���mQ����	�e�#��W���������_�X��ʲ6�u�I'�,�}; @�����W��/�����������O��3�|�m�c�=��1�cѪcY~�z��O~iD�{1^V��cGt��T3lmb���<�R�4�_��2�/�g�)��	�DabA* M��) 2v&0��@��2������u�w^J�_��˱aQ�j�>U���X��s�|<��h�y�DG���@�ܜ �$�k�%���bup~Q�����r���N������S���Z�u�~��>�^k��\V'��3���m��Sy~7�\�˾V�7�R ����6���m��� �*I5g��I�J���tߑ���[6F��ZҶi���.�v4��V��.P3��c~B�����<�W�KS���0�\�Ҡ��z��a���u�����|n���DM�g�z��@:��E�UGp H��
2R�(]Af^����}�X����i��*}Ϯ���)~-�J�3����v�9�G�: �َ��� �[��vu_D��EJ^����zǝ�ܯK�n� 9GDz5	�+���'�[����)JqT9s�d�><9*�
��u�`;tݧQ��)�u,�z��P�NN�"F�:��sLF�*�j�I�K�,�г��:���d��g��ϼ�P� ��Ƹ��dobx3{��5��=M��hxq��mbe�g�)��Q�����Ʉ�g�����C�8�W�6�����`��p��� ���8�;��R���	f0�Hg�X��S�*}?1(*8���=�����u�������1��vc������\~d�,r (�|�ﱤ=C(m�b �/�!)Yr�X3R�4�h�v1��ڲކΈs;��u��]�L�$X�0���n�k-zo���1�ܼ�y��Z99{�����yEEW4���v6���+v�c���Z3RL���YK%`	�j	�«�Ɯk���3�#�L���Z�qNַ���C)��.��&�`O΁X3��u��U��%�8q$� 0 sU��Xg�lR��@z�u�.�b���v��DV�Т}��շ�ֵd�U0�?_��Ε���~�]d�kl[��e����+��%�D����;��	i�_�2���^a�3
�˱����&���^1���F,���"~d�����6�`V������B�0�:�L�LN��ע�k���Gf�gd
���(;�2 �t�a3�m�4Ale���oz�������������x_���I'�Z��  
�Z��x|f{�����?����[��z;)K3���_7�� ���t�K�4��1��p�`�O��R�v���-�,�|��K��`u��8�F�Y5��]r]o��9=���<)i��p焪�3��M�h�[ð֚�Ӽ;����M�|���悠)��fdRk�j�bq�8Xt��w�$��Q��|������3r*�K~n���P۳� E|��;sqɑT0N%�O�}k�����:?�(�3DK{!�_��}ӈF3�mO]l��C7��~=�^�hӅ�"��)�(��w{��$�Z���"�`�%=����T����4����tC��?��z�>椅Qzx��t)?�D_�Z��a�7?�S�Qʏ6�~�.,Q�C�/�\�.��/
(�u��)��Q�n�� N4�d���e��j�9z�L���UB��R��ݒC??���`�t�ӹ�X��P[ ��`� =HQH.u#��$dB/O�
 X<OW�)�p����S�3ң`�AUG%퉨�iEQ�	[ˠ89��Y����d�[#mP�i<U�_ �k�E��O��д�%m�����s�G`[1@A���XWp �~g	���bRP���Ԕ�o��X	@�����c<D� f��y{F�s>Ȉ}NK�3@}��TIۀ����]o��	댜G�éϘ�O>:{� �`�̃�NFi:��n�[ͣ��C�g1��Y������AB>�kF���o粫X���9Wm���d�G>ѹ���c��Z�D�3�M����
�W���@Wtq�^�C�k�K�(�}x]�+z��n�vF��3Z`���tL	��=>��9�(�B=���u��t_uͪüa�S��/�9}�����d?O�O�].��c���Be,�%�VfVV����c��;kE}E���%d9�=l��ڇ�}�c�E�@�I��\(h��UƠ��/%�b�XX�� �-_J0�~/V&\ٙ9Z:)��Uv��Zk]�I8�@��+�L#�U)up�R�8�����$�#����A��jc(�+���&������@��돬o��i�?������S��Ԙ���N:Y.�`  �Ii�����S�/��ǵ��,ҵ�`�1~�d�e��{�zi���G�L��	y�+��8��acA<�[���W�/΍Mf~ǄTV��G�LQ&P��)J�oc�	�[�M�F��hNs1?{�G��h�i
��uM�׉�&m�^��F�3O�5��`9��OfΣle^^����)M'/���J������S���]��u��yiLܰ�� 1$N�@�����iW�m[@s��nzm�i*�U]Α��GIU��=��q���E��>Z�L�wf0z��l���z:*���Hu��W]���D�nI�Ĥ�1{�v�t��&�s�J�%E� ��3-�����t�3�!���唀�<ްS
"a�O2ί^9��X[��It��|�L�������ܽGD� !U4���c��<?�8�^G`�'V G:��@)#^�J�G�,"U�?M�F�(T_�d@;�9�����HRH�T�ހ�X�y�	�1�<FO��R��\��U�::P��9�\�z��^"�B �.ǭ�~����X���?���dy�z�ڢO��}@y89�]�k��9�cN���R)�y(�������A�I���ژ��� ��{����s�,������4w��
J�k��1�5ܺ�eo����28��*4��Dk���.P���?�X"U���c�s�.���5��<��!�_߂�
1����Gc9���\���\��D�P�������D/i1�{��`���D��c� z��?���,�U�k�c�IlLq�C_��8��%s�(�-��(y�U�*GΖp�^x3�)鹮N�ْ�%�����.�oc�v>���	W��=Ig���E:g��� �	 �����9����i�I�M���@!N�^����$@��ωs��.�[�z���{����a��S�sr�F�J�*�e5��)e�9OW&�'�aM�o��4Ev��4�dl�.���7E}����I'�<+q �K�~��OF���|j�z75��*��^';w�Q�8)�`�R�Sd�I~+hz�5'���6J#a���w�ͤ�ߦj ��?�xl��T6:�w���t�$= M*B�����1��	��d�l��ְ�F���������ib��(���d(��Z<�Ŕ�=�;���J���D�{���y�E��Y�ZL��S��y5�T����q��$���n�o~F}i�E�P���z����� ?���#: plGFU2F�[E�Eҍ�e�!��^Ϲԇ�I[HQC���,��d7T_2HW��Ǚ��dZ">Y�l�@� � T߾�G#ϵ�o���1��S�k$:�t��v_�B%mI�a��h�xW�����|�zR�]�Ot�B =�ϯ@ ���Hcpv�@<6�ZJT2���-�� �	�s�pj�X. � l  p�h�>xq�I]��ے�Q��IX\�9�X���(�Cz���(��ڇ�l�ޢ�|b�� NR��h~������@:�z���4]�Q]8�c��e��V�_�e�O8_ ��	�ݏ&T>�M�7c�Ȯt�q�1��z�oi�˜ 輟�wH��:d:)�5f��r��=�pq�P\�~�[�a4��k{g���6c�"+����4��C:*Dۨ�
4��<��AT�.�Mj���gV�k}����ꘜ��YńI�ʵ�1}Ӊ�94hݪl\kq{�~h��͠r�9;�Z��@�5M�@UR���N���e�J�kf���/�7��:",����)�H.���(��ͯd>[#�"�|��{pه~;�I'/L�X� �2�?��ͱ�'g|�3��,(Rz}c4er��!`3u�������ŭ_q'����8��w'��6:$����;^��鱜�9Iw��
jJYV&�/#F\���9����~P���:UP'�t��R٫��7������?�������?�؟^>f�J���.*:@V�F�Ϸ�, ����$Ā{�-/�W �}p+��eP���r��M.�Q�JM�X��������G�#�iBS
/S���c�H���\�S�~<�f u��Q�<�h~���2�L'��5��V�Э���0���9�^���f���q��Ntu~*�Ze'n?��FkIj�
��t�YM>u�LfG���&msTY���j��RP�1�rN��yP�人�Q"̷f��Be���,�d�=ґN�7gl�KD����`��Ք�ԲL���0�������Ak�lmӁ����g�^�`Q��I�G�#�95��U�Nņ�:�c�:���@��Si�}�-̇�L����	�� �[pu�i�d��щHap� ��En�H[q�<ņ�Jɥ 4� W �?�O��]�i��uI@+�ʟYʽ�rALT����S �F����#���vjn?N�ç)9/P�|1��{p�o�s���)�!�%_����3q0�9��_h�
�hܬ�����85��O_O����(Q��@�.(���� J�<����rmW� '��hb�4!�)�#��L$8�h[8HPT9��P�[�=;!��GAh��qI!ڷ�pe|-���m��@Y@i>�3N3� ̵�����3�5�o�LϨW�]���YM�?욵y��=t~��xWf��}������W2��:��R�c�Ǎ��5��mX+{�z����,���;I��Z'{1�фFmfvX��e?�_`H�!E�CEά6��i�����纨���������l��Q�>�c�XV�O�HT/M��2L;���w���l��ML����ݗ��_�=	Ͽ��4��0��`<!�y-��D#�ٵ�?6��p��Z�&��xLS3�0Qg!Z���� >��bz�&��CT?�[ާ?%u�L�y"]*6b��Mu���t)Ƶ�I3�e��ܳ�SVf������������uoxf>��ye&�	�:餓N��! �����?���g0x�Sw��+�cS[�cG�{M՛��dpO8�S >����zd	X�xm�������t ��,y &���yb��eV.��'�.���2�m�j&8���6�F�Sxo����P�
t��d�|�L9(=�~H.NT�r�DG�h ��n��ҝl�6#1��+ׇ���Y7t�KNS0�$Vq0Rw��q7���j�/8f�U߾V���c��m��t�D��K�S�Ѥ��m��t�!c��M���v�n�e��1O�V��E�*s�`�!9���.g�Ňz��ϸ����S�����&�?�����eo1�s>��>�C�������x�.u���,N�0k�����$<���{���߱[�61��%G����㻉y����1E�+����%9 ��?����s0�"7g����z��<�`Uy���CQ�&Ds�e�����|�;3�b*��σ+�<���L]��[f/@���\��Ħ� �SYAÂ�� bf��D�������6nrppH_�{�i}] �w���w理+������3OOY�����^�m0d]e�����)��)�n�O��`(�#W&t��'΍���"���r���\&�<���ib>}36�����Y煖>��Ç<�*����L�~vO��e��c����,7,�K�S0�*��\�z�:m�ֲ�~��d\>�x�p��s|���?j|[c�:�J���y#�K��p�}تc��������Nо��q��)��1�
�6;�.m,/UN�^��9�t:_.;�C��lM�^��L[�6�g�*���
�@EP ��uq�]v	��� MC�$�0�4R'�8R��	��\�+�"�XwI]�*��^�8M�p�*V,�
��]��F��=E̥�������8�������ɍ���f�ǽ�?�����o����_�w.̥�_��'�I'�t�D�� @[����?8�����i5��u~X��j%e��.� Z�9h�Pr����eH�
���S���a�v�a�Y�9���nt��&&�e� �r!�A<��\����J"���U�w:���P�l�Z��&�d�u��:�d�~�X��#���%n��q|�N��Y��P2���E�j^��tr����N����~]b�n������d���k]���uʇ�u�k��1uߪ�i]�}�܇.v}C-��q=p0�ӖʼX�c��I��&��;s����D�{W����� �������|������/-rd̴o	<GY��># �6�# �d�Ə^Rʁ�>?|���i+�����Q�x�r���g����~�	

J! ����� ��Պ�E��� ����sP�g�|Z��q-|�٪���@��7D�������Oh�����\� Q'c�AI�)����a^���e㇒R/ �z�v��F��:)7�۠.튺��$�G�`��
8����ad�ւ)�m��c���T�?����pqů���^�.~v	�4�;��Ʊm��'9CT�ڀΆ�-쩏����BzxL*���Z�@v�DLƫ}/BuS�F6XCl�/Y�n������{�c����l}���D�I'�t��Q{�����$�	}v��r*1��b����7X�g��QP܇�����_��6F���x������̢7�o�To"�d��Ƅ�Fb�$�agN�I0��������F
�9W_�ǖ��z��U�]T������}����7?�7q�邏N:�+�p ��alPf�u��u9�=جD��z@˅��~W��:	(���`t;e ЭMJ����q���4��n�m���Cтϲ�gW�h ��J�ϞiJ��6�0"X�	;�3BJ�&#��Cɡ��Z6x.������IJ���פ�1�1�D���
��r����M������-��$�o�V:g��y�9�=ז;�����ֿ���]��E��kM`A�K�y��[[�7�jv�˯��o+�<j�e�:-S�_�}�����S��Ps�<ԫ�t�qv�1\�`yT�i�.�Kd��-����l)m�b��� @�x�}N���O2)h|Y�����= �<;N�R�o��=���"�ۙ+��=�Q�����e��l<bTP�����bx���j�0k���'���J��/�y�����g���k"*פ������RJ�u�u9���s@����"�'cS_�Կ��nJ@:���b���@q����Y}y�g��ޕ󍶿��� �+E�+��M#�@��,/�hX�u�N�!�c�H'P�� :�u�AI���q�6��� ��{��p��
ǎɨ$�����T%���2��*7#�q(5��=���`��I/�`u�y$4ΦVK�-��S���s��m���!��S-ݨ�����k�M��#js�t�ÿH��:.���﯂����ܶW���<Lӎj��b�\��ֽ���������D��I]���??�#����:���FNa׼c�k��?�K]��f;�-mbC^鶞���9>�ϔ�|�d�����ۄR�ރ0[r�Mu�2�X0�&�`CT�z4W��R��A�>E����4}�����@������5�ۼ�S������/�RRD7��y�*��_͛��N�
��җ��ݼ~�χ���s�!f{_�n^�N:��[#H�S��O{��ͩ�L�B�y15�˂G��l�zH�`=;`Ƒ3���ԓ*l H��Ȥ���ҥ�IQ^y%Ž��Z,�A+�M,QV��P|*+&��ra	������8A���Ĺy`m#rC��� ����'�Hd%����\'���:y��:���g��z)ҩ��Kkc9os����l�+ˋ�[�;� X�B�stّ��{�u��u�度���n�V.�eJ�P���<����x���j|܀�ȎW����Wi��8<��ꚞ�lP�\� +��\�MblJ6?��`�2qL�T�P[�g�J\[sqZ'�_A�TVf9�|a=��ʉk�p_��zk�mP���ܵu_��)*8�1R�po�S��j���� t��i7gv���m�K�ޛ����͌͘ۓ�R`l1&�ۭ����ӱ�T����y�6�ׯ♊�k���H�w6����~��mi<���/f�׽����>۝�&�����N^����ңm38��:��#��R��pns�Dx�m�@}�¬�l��b(�;;�4	���W�B�&B*g�9V���8�1\�m`$Hue��-=�g�4��}�=�tP�.<9c��{{�d��1�����N:�d��������������'W��ʻ>��4Hz89a}4|�!=Pҧ�	�5:#�qF`t)�r�b��s��Itr������Il�`~����8{�i����7ބ|2anH&5��ړVc|&��9ѫ~L�;��WS�Z����'�1�U�:��߃�N�������)w�s7)p��5���m�:YG�e�˔y��%�o��͑��cזS0n1^�Z����-��y�e����:UX[k�u*��.���������8��?+;_4kG�^�|�z���A�?�ʘ�߂�����%��)�t�L`��̙������P9%EvC&c~�{��c-�HuB��^8�?�|N��`�T�J*��,G���}���-�xT�9���0S��>տ�Ι%���K��?;��ַT�� ��~B /e9�{������S���<c��+b �Sw}G�jP���󇵮p>���۠0Ei���{�Ϩ�^��B_S]�^��G:��E��	�o�a
ֈ�����1ʄ���3����~Om�p�h�E��p�y������s�����"�;�v/Z#ly���^y����=7��c-��Z"�N�@о��_7��[��{���U�+O��UNu8L��6mul��>�߳�D'Ш��{*ݳ~$�����^`�1`�^�����[(B0d�?�&���$�A��I���Y�� I�W2o@
�IEȯ_	���\�2�:WN`����#�O}řc�TI���6J1�<U�a>��43�o��|�U��.�N'�t��� �P����>�����?�~��O�w]?��z[Р���J%R�+@]E�{ۼO4�@H9]��*��U ��`�,��iĺ��|qh@�>�|��|S��N<�;�+��)m�c�0J;`�!W�|���T�rl�AM�)�O�[s��2ړy\ĕ}t&k��DG�ye���8�\��H�<�ز�w�Vr$Xo��-�m�N���*+��l/�>�w#�Z��d�c��;X`G�N���o�����k��߬�* ��{[V��y�d���1�j�c���v�xO+u���;�c�Ƽ^��Μ_��拾?1@��M��c�������)u�պ��<@����\��Sy �q���	��Q�g��|U�@�	S��:��a���g$_���ի���O׀�T�Ŵ2����%Ң�#H/��i�}���3=>R�yu�~�3o��7_̫�(�=��S��m (��P��tP������w*����k�}���
S5�'���S���.�������#�dR�ɻ"����^�m0�6(�KJ�P�j��m��P�ի>�Šnk���r��}#����J��/����b DB�}�e�A�u|o`�~w`^�7ԗ��A�v��`k�D�n��}I�ӱ���߫�}(Y|�$p�x�8�kkYv���٣<��%��0�T�r���{\�v۹��%�Y|��뀻|\���7-,���w�l�Զm�$���m��9OV-y��x��u�1&�f���zM�e�����u[��� z�V.���i��_���s��?�@�%MQ�@=c1�o¾��O�	��C�6����
����w�f�'��9���B�U%t�i��ݳwu�n�teT߬��z�苛˛����˷�y{s����,H��I'�t�r�����/���y�������?�a.��Q��҆�&E?������E�o�3_%�u�4#��l��dbpq�0F�Q������N%t���&���a��$�O&�FƁ@IC��5�!����tL.��ID7�5NF�9@k�TC�1:��_���n������23���E@<Nu�k�m���Ǧ~;y!�5���c��	{Q�=7���|~F������ �V��d�\\�ٖ�%<p�#�y�,��V,�'f�T0��Ѽ��wD������MF���YF��q}.��OF�e�.st)0��G��Y^��ci�f�a
���˞�y��� mG@rq�9�+r6�l�I�e�GcQjƏ�,@%-����  <�	��W<_�e�\��:�Ae�E��{��(�����:���8>5�q�m��̇��9��7sU�#@{D�k����ä$� 8J��p��s� ���x�)�h�����wu�2 �EN!�pV�R;�=�� ���J�cY�0m�J�Mt"A��������3j�I8�����(R&����s�I'��l�P�=���e9b��dW�t���\ڢ-���z������NF�N.���;�*�����S��E���N%x�����4�4rL#M��`^It=���Jy�	@�9(�����g  ���zo)�����QeBԿ��Z�e��*�*��Ϊ��n�/��yV'����F_�W����+��\�z߳������ :餓gd� �A��q������3_��WO����ͽG��zn%�6�0o�df.9o�#}�g��d�rF�x�]��E�=z��[糄M �ǈ�Y��>zp�3���s8��Ɋ'-&E�78�Gͮ�c�/�z�)�O��{���w�:&�ֳ�Ez�٣Ӧc��(�}+iN̽��Y�'�9/w�I'�t�o�ĸ'I֌ϭ�^�,_EB��$ ����K��ҙ����ca��A��jx�g8�	��0�Qļ1��Ҍ�*�x;%'|wI~̆��@|���uA�N|��
)��O增`���?4 >gu]~S�;h��ssc�� �>
q`Hۄ�Ā��\��@ nނ� #J}�K��N�d��nmc$�Ő��E]_ԓ)�=���t�e��_�,Չ :E?%�ഐ�����55wS������<��{Gto �z 1
��	�?�h`(@J������d����Oe�? �uCZ	�%����-3H���,�����雛7`1葃�����pJ��	>�����t�I'�����I'�l �zTi aL��[ky�֛ޡ���G|ռ�7	�����\&��9�^�1g#��I�d�D.��h0b�\��UJ���F �O�������U� ݔ������u�^o��oo�_����y���<��C���7;餓Nʾ  �(��-�Ǐ��n����9��w �F�94/�tJӝ�"ѕ"��Q>�����xv<-�q��.�Ԭm�J)�2�r� �F�3�@tp�O�4*���P: O���Ej�k8H,���	��L��)}"eiS����eDE+,��4�@���ɐ�%�1u`��R��C����,����s��϶��V��\�I'��F�թ��qk��S�Rd��o[�������m}��o�k,���:^���Ƅ-봍��^n�,k����*{q��L�EQ�^>�9���m����$7��W� ' �& �ɑ����?N��mY��u%�D_�qu�P������(�g�.P�#��	����4�uyw'�� �X��Q��$`������c����SԿ���Ö�+"�%2u^e�3��|甴(6���.����+����Wu<�"�����g��@.z�q4�zG������h�q�%������p��W��<9V�72�y�-ʥ6��~��۠����cv�x,H��sGN#���fF�'��R��� ߸#E�"a��(��kv���A�|�����dݹ�%<�/[v�bZ]S��j��m���j���8#��ߦ+�N6���ˏ�·�ȷu��D캇�n'|h�e{lR־�����g��9���e`�7���,�Yf�X���o��|C������{>/`1��ӑR�|�3�����a����>��FS�[��oZ�m���^�m9܋����,�L�!�~/�}%�<JQVq�dU��/���qU�o�{|W�����;餓� ��r׿���/����4xȟ`o3���, ��~�ā( ��Z�:�+{ ��0h^�� ��g��7���;l5B%<�Ȩcy�МT�A=�ky�hQcP:���J��7� �*���qR��O�i��[�p'��'�8N�wF��uoÄ���v��R�8�ŉ<�(ܞ^����*:rP�0�>g�|	��勩�\N�O�i��j;AE��K���c��Wڦ������n.�t��N�iwG�I��[s]ד�K�N�
��Eox��:lY=�����;<j�r����z �G8�Dռ^���3.�}�٥3�Q������@ �-G�$N� z��O�tT��Sz0��N1V����?{ͩ �WR.�w8��O�y���S��뉹�4!`ʉ��Y��G ��uF���Z�� ��/���90�E���^�Z��S��nYm  ��IDATiD��Z��v�� B}�3k�\�v䀁{��"��W}��4���$>պ��0!g	��4	 �U�����whrа�lu~@ �/�e�����<���@�N���'4�t��%�A�\;8�8#���x����1r��E[��|���}˶5��V(�%���9����ɒ%��yҞ�m�d��?�ņr���x=� L6��#�wY<�-�em��C��Ouf�|F�udQ���?'��'5�ۓ�|�_�W���$mL�m�>d�`h�@���̅2ح����ֵ�@N�,%�?:��,Ӟ�=OoK��%X{�Y�#E��{�:bC�E���8��|ͤL�&�0�X�`Iв�JZ��M�3`��_2$���)��G�2�T<����gө�duN �t��R٫��4
�i>=�?����������O���YYU���������87;�1�'Vbщ@�c���� ��g'_fvr	�,�+%Z��6��u g��W���ꇷ*8x�������e��k�C�1�Z��o�U��FYں��	i�����3�:A���F����1#���w��oe!�.����j�k���?�z|�����������I'�t����揗*kt:�T��&D�8��5}d3�^/<�6�V:�����B�w �S�@z X\��C�t��9suӣk"���P�+�L�^�'���`vI�O���v ���e����/��(� h葚@A|r0(�}��@�G 4��z��Pγn��.��& f>`g����v� H?~���؀��9` ���M#� v�`/�m��?�]���k���
j�鸠tH+���C9��e?�
r� ��ړS��u]~��	�34� #gGl�w8e`Ϩ�ޚ���#J��Nv)k{��������3�Ȯq�%ժ���Ʊ�,��������e��ONI��T�o��,�m��Ԗ��m��fYs�`��y}��NB�����LA��	���c�8�{���7�7n�
���i!�nT ��U�̘pNp$�`���#A�!��X�>�A@�@�>�\��z��/~����˿�����O���0�W�N:餓%r ����������ٗ����mw!@\�$�]}�����Rz�<S/.�i�ɕ¢�Y<y��{B����SAnȔ������ciO��V�km���6r�h���T� ��a�jץ�����d���{�|�N'
�9�z 7h��^�h�ePO?��9uC3-C�~��T����.Y/�ց����kz#�{�U7�{�n�Β8���v{YEӳ��}�lrO�j���vw�s�W���JI�d6+阆�T����/�_o�������7�ϟ�I�ۍ��nkumrB<�M;��G�}���9�)�\�:wDi0p��#���x�	rǏ��hQyz����F��X��6�!�|i�c��#�<��y]<���)E��,��cD��
f%(��%S<b J{8�y ���G���U��n�-��[Ke��Y���@Rۯ�V��H��T�ڠ>�� ����1R��+�U]��BW����8x x�%�	nn˂ڠ2#���
�s@�Oe�! ���0�o�P7D�S��m����"s[4��>�y��������RB�ɶ�8���ʧ����������7�qJ���ٵh]����6Ӈ��Ļ�~6z��>iw�M�n]p��.�W���UW�d�<)_�m&���7�׶���'���*�[�b�7�?��#+s<��i�?�IZ��޸9ND��k�86�k�`0��j8F��zF� ����\�>�h�p����&;1�2b%�Ţ�v�#�bB���T^U�~�ҍ��OST�ޤ�3��F��������ߘ7����]ٟ�gWWWSӱ t�I'Kd� 4�����Ϟʻ7���z�:���^6�l�jDDu�Q>N�k+���{�8'��;��
c���P�}~����耞:8��P���˼b���o��eZc4�J%�¦�B�I�U���O��9��Y�*�UϏ��ĩk6)�$���Dրt���<�q��W�&Z?�P'�t�I'�t���K6�t�g�ɇ��5f&������������2� h`
�~j��R�����(�	��G%E��NN ������*�3 ��q<K�����)�'cf��1�l̀v&�
���MC�H%@�֗>�~� ��ޟv��� {(��L6ⶀ� ��hig�{"�����P�}�,# |Q���[I�H-��^�XI �������� ���0]���7.���%o����$v�N������yu�ɋ�n,褓N:��P�v|ߎ�dgv�Gt�2k����x�U��7G���G'7����iZN�/4E�1I�$x��c50�r	"���Y����q٤�O��s�XWD�a�:��L�	�$�.	B�� ��gH`��� ;���=�������_����X M'�t��9�=sg��|��z���=w��p����t�d��Q������<�pv��O=��ی��*ǃ2�Y(O��qL�dr`���9�I{,9Z�xC�7&�������J~KgQ/�S�:kM*3�O<�4�����4꿙�G��"+N�;z_�A�'��&��WdU�)-������ٙ���}_�;��N:餓�Ml���d�B��	���Ԁ�8/ج�ʊ��D��W�� DY?��ƅi���;~�N=G���eℌ�S�ǔX/+>�F#�.��aл�e�I�<J-��)a��OI +]���t�y}ċ����o�s�u�uEm��)�ʒ��e�n��+�
�?G�^u�����rf�,8t(��lx�1�6�2�L�-[jo/N�Y��܏�'����O�a:Ū�uZ�����x;���\qⲨ��8v[R]B?�h�������6?�sލ1G�$�Uw0!00F=�&�G� ��p�}H��j?�:Jy�%�k!�t� >y�J��|_�	F�e.�=�k�:�0��a������������XvVp��1��7�:��F���Tt�ͬ�_�y�����lf����N:YA� `���9��"�)h��R)䇵�����J�f^��������7�H��<�����S&���}:!H}|����ש��K���f����!��g��W:1�5� �0�N��P�R�KypZ� ��dk������F�����˷��򂚚ǫw1}�t
\��U6���a��]�Ø���c��XӢw �U+�~�u��1���^s��>Ʋ����W<���n��6���zm9l��s�Kٶ_lc�Y��v�o)� 5�nP�I���+���9[eg��	o�u����țA_%�$�T�`[)�=�I�׈#��v���<a�+�T�뤀~`0#T�a	dZ�����w�EKO�!�]�8*X+�:6�����w/I;�D�N�ZQ�_J��٨b�O$�&/ߩTzLR�4���29��v���KQ}��{NQ	��&u�Ǻ�.��r:5y^���v�ւ{�.d���9 �Nj��9���!�����1��#��~�OS� �˒�"��mD��Ď?�Lk��:�;����)�qR��hO���)[q���'��˄yXf�P�dn�ޤ=�RtYa����+(�'$A�Z#�G�a������?c8	��� �*\.r%�:X<<�D�]V^�a�Ri^\�뤓N+�p 𓧇�e~��O�{?���-�x�>��Łً5'�c���I.�P��@�p��K��cF���	���M�f3����f1�,�yXdVw��9��3w6j��.iJ��
�&hS�Y���W?��0�?ЖIK-Aa[��K�(��iq��l��]ιg����teFDfduUw�R�W��߽��\��22󋈤j�V��d"�Mixm�}�t������W�F�Z�+9�����nA�G%�r�Vm��T�˾��_�=�{�������.���4�@R�Z]�m9ђWH��8خ9�V��*OD-_��5k�t��w��`3��pk�V���v�|7صG�~)�ntxt*[<K�Q����-:�MŶ�,�8�ݢb���=�.�.�E-���͍$�]�g�=����{�����qXn�Nnx�����l}źիc��x��cV�?�K���?�´3�����]���9��P��^iAJך��k(?c��,�� �3ԡ�z����0C�p�EF���M��r���ڒ nӦ���`����#B���Ϛ�7�,n��8Q�zc�G��l����!��;���ļ�=K�+�M�vůuy��Fm\�&��5)�N?���{��w?�A���t�vӔvÊ�fn��+3�;g��(W-�﮵c���8���{�˻n�����K b]�+�\)m����ȉ����]�N���焒9F&N�(&慼����+2&�g)��:h�O�̷���,�Rڙ�2����Z����$��1��X���[�����̇�uJ���� կº��,���~P�~�O|��Ë�7e�6����`322��� \'d>���n����O��7~��'W�V?��B���BK*M';p`e�bgk���cG�����Q�(m�õ��'(�h�F����X ��hF%�&э2V(n�I�ۆU���#���䙕B�Ҍ�b�
�8e[evXo��E�Y����V|r�n�LWϻ��ń5��a�k��.꼯vt����Cy��M���y,�뾠�I�]���/@���a�,��Ca�v�Z�����xim���}�:㮞o&�2��	_G�]jH�C�$ִ l�8�F ~�J-���0l���<q��H����FgO��؍��I�tFB�GB���{�s�t���w\�L1� nV�
(�qG��1� �v#��]�g��y^�9�Ê;�!���Ȟ-3��q��5?�ɳ�l�֯�ұ�Qw튶�7���zOp��h+���2�Ҧ����/s6<��N�
yi�k&4u��I_Q�>P����q�p	9�s��\�b�fj�K�9��Y�Lst�� ���6�����o��o ��/� �sOn[jU�@�ʏ�������j����� ԭ52222�\N/�>�O��k��W�����z�Uxf��0�N�w���3J����f1
@�C�-�k&Ҭ��'	��O��(�t1W���m��ل&5bI��1�B)��L.�\��2�$UXF��arl�t_9��J�,��U��u,��̓�� M�v��pH���f)}�!+��1�eC�4)��ʩZyf��������{�F3���4���nO��0�Ҍ{��@oc�Ot+Cm|fT�������{h誵^ܖK�M�t���	�Yk��~�sǻ��w����� �rl�O��6*�[I�<l��ƌ�=o�q�f26�.�\�\��5�1\6ל���Ū�����/u��a��cEכc7J��nw̡�������=�k�����F�5czo@��l$���k0��c��4�Y�ol�+��2�Ɵ���CTf+�C68_�J� DA�7�_��r�f%�f#����Fް �C������I�=H'�� ��vͱ}�T-�;��(3�W/^����Ͽ{v6{�j�����@FF��j Pul�uf���j��_��+��K8{zn_�k=U���"�l�$��U!�\RE�l�Y��񔏼�-�kq�Z\N�E]!U���>��S^����U:Pb����AS@��D�$�[ �1�-d�O��T�w�J�y��Ћ���zT��%��q�yػL�79cT��xT�6(sE�Q�ɲ�W��X!��븺�.پƲ�|��{�I>v��1��Jj���Ưi�+��
�7�_t[�
��l÷:��E�X/�ݟ�}>�R�v�gw���o���U�T���>݁�`�8q������%s��v��vH��{~7��>8�a�F��y�81>}>�z�ciG�8����^�t7N�4��v��8����.%�C�|���%���5�@��1|fk����P��2(�a��`��( �6�C���ɚB�ߠF��{ʇ���d�`q>�l��0�xn�=1O���^�_�B#/�+��v�T>�����h��"vQ�|^ȓ��f�Ծt��ꍗ_�ZQL�2��3@�C}�222� <\����c�e����\�@�#��m=ĿZR, ��h�>+�B����Ո���a1-	+�pwכּL��^�����~Q.\cC��bנB:�����ҋ�`9J@�/R�2���e���,��Y�F@e���iF<����ضM@�^��A��W�X�����z(��4f�	���n��`_�R+���t�υm>t��mPؽ$9Zl���vt�}~32F	���3��P�m�	�vdddtCX���1��ƾ}�.峍Sw�������X�㌞��+�������������#���hE.�x}�Ώ^�6����O�1ظ�ˬG>�t!�f��q���#�c�,��]�8ܿ�)P�l�^��~����Y?e$ +��r,��渢[0��о���L�-!�322:`���+WW��������ŭ*lw2X`��z*�*���J�$��lT��5I�}G�n�Vb��W�zu��~k��8��g�a&�u=T�PD�|� mu������fw1+��G1��46b��P=Zl�vC0q[�:R��_��ԣ �2x�yߤ� 	 (��Х���>l�=0e�@~P����fd�
Խ�Ѯ��f&�HR�ud�ѣ�4->#######c��k0�@n�۴p����i�>������M2Д�J��S���mۯ0�>��$6�`Ȅ;p�����}�,Ӽ�p%ނ����6�6��IvҌ��,opA<H�NfG��u�#C���.`1-���g�=0�������X�^ ��vVz>���ܯ�ʇ����G�W��T�����rHx@z��g�h�7w�L�ǎ�Q'橯	3��RAi8��-h{P= �\��=���
���4d	�&>@�$��+���+��5GH�ף (���r_���,����#ɲ���(�A*riǃ �����V�l�{�]��Y�|�w����D�=g�;~�>0֠kU;ݸ�mw���N.k�M�L�Jc�Tqhk���xo�<�Z$������K�GFb� �)w��0�ݳ��]��j���{0ڥԆ�l�qӺ'�Ha���ă�*ٮg����wY�]@̑[�M�7�9�'�]�Y� I���[�~�m�ߜј�uQu�+~u(Ds�~$��|gH�3H��J8�{��juwt�H^�� ��h\��
��c��g"�#0�n�u<\N��dH�DV��S��c(����pa�]�6�xQ9l�td9"2��Q�yK�蘩�Vˉ�5"?�|��r��J[�h~�he��I>��CY9�	ǟ�-�u���^WO7!��R[��������o_�������~��.Nf� R�����!" �/]����������⏙�>p&^ד��#���te�Y�� D*���r*���U��*���x�%�a� ��:a����}j����OkC�-�(�]LfE~H��:��� �6"d���R��K+�a A�[cj�D�G��RÉ��ј  �?��H6b���P���5Q����H�VF'�h�2F���gS�<H96�8��#�Z�}��M�=�]d4�ezW����ާ}�>e�O9���Ԅ1֩��$�жvy"|�-��SbKy[�&����I��y�+��sH�LA7C 6����
���F�����:��q׷���t�>�}=|���ю�7���s��f��`��bqz���p����������9�b���DzK>EE��I�bz�'�xG�;�ݖ43>3�8�CD!��l,�7�#K������O =��yq{�?w��9)�3!���Ҕ����`��K��I*~�V�&^E�1�v��/e�s��7�W�p;�>o��G~����_��/�7��ܮ��  ##�} �����&77/. �(���U(�;E]�����#=��ыT*���w�i\XW������$!�l��,;t�>r��C�h�\!cgSդ��K��\����PB��	X���kn�J FH���)�>i�Ӂ��
 ���ҏ����qD��D$��G�ʀ�c�̃��`��F*�z$!	V$�rpc����T�
<���c�j��v��ȹ�۰�3�M�Z{X��n�*h�>ɝ�=�dW5N����RR+~u*c�y��fIv�T�Gꆕ�.}�i��t��'j��Bәv��h�F׹vc#���ދߓ��_ r����3>���~_���uHn�ȏ�yjS�����7�>=�#�{ޜb�������K_������V��Q�����:��\b�;�nI�^|K��;鲻<?C�lRF��uy�v��:۾؝��v]Q��Y���/Yqd�����]*#y��@�$���ׂjP<�\B��v�s���-CEy�,�)�z�O&e�����h�rX�ӥQ�E#m�ƭR>Ɇ����2i}q�C��oX◊��U�M3o
��
T���'��j�J5�����>�|�ݯ�}���½zz322�� ԓ�+}r~25�a
�O�꣼K�Xfub�ʬ8%H�;�zzH��=o#{-�bq}QD�+�ȣə��e��W@VY����7bp��Bo���~���d2��U�߬�^2�
�2H�)ԣ�� ���۾)R ���"Z��9��(��ZqL|g���Ѩ�T)ҦFc��hg{��G��Q��:<Zm�ݯ��X]��b�bUІ�����K_R�XAk��>��V��jD��=��u ��=ѭ�>L�ZXkQ{��xۆ�"׍R� ���/n<���,1@�_�d������xh��].?�^�s"��u�)�Oȃҩ�<�m1�6�!Hz&e��ǖ@�/�N���tD9�\�._�.e��^����j�غ
bAuoXU�M˩�+�|w{�;���P��_tZ"=h��jA}d� �e�V
��/�Q1�l�z�(i���i�����'��L�����1\��.ܞ��O��\���4�ʋ2�sV��+���d��o��3�J�R���W.�EY�]&'�/�|�㟚i'��i����ш! ��_}y��}���/�y�\���UVX�J;c��BR=�w<��*t�Z~_L���2�\ZEV\�e/Yc�2[P4�J�u���8ܤX�B6����8<�EVF! _S)â��+���`����T)�p��`�y��hL [��D�~�x} �݉Q�%���'BడA;a�c�A�^���CX��n�ph��ckSf�^uv����W���Q\��{ϋ���H�l�C��?�Ou�(������;���2���]�Qէ�j�Ѱ�[�ִ�09����E@+�wL_�X�M���L�t����!x��G^Å@K��AN�E����A����l_����^�eL���u~�$���ZMeҟ�'�P�5ߒ��I��@F����ލC3��C{���#C~��c��g�L D{1��<�Z�<,�y:�|�%V����.T�E\��x?n����s�(��}}����Oj�o��!gE��w�����9jh$��b�!��F��" ��!D@�ǡf��^f��s8�~��nO�.+��k㺌��cF� ����o�|�7|�{���Ͽ����,.���}�k�l�Z�EO�ZNq�s���oUO�'.��u�
�2�a1����Fܹ2\��L��q�~��V��IY���ʈ��+% �c Z��� @��ˡ��ĉq�LS�&\��u��/%�}��ȋ�1�
��1�E�1 @���@c(�UQ��=V���} ���ٮu!����M��z,iW�&�]�p0c���c� ��]F�� �Q���y�z���	~f�'���ә��3'�fէ#��#����e�|�٩�i��ԓ�8~�c[��?=qy>ߓ�"�І���?�Ҝ]p~Y�i�y���E �J?��T����t�?�E��$+͏s�N�gEu�
�(kw�����[��{0��a2�h�����`�������?��M
M�Fy�;c,`�)z��qI��qo�� ��2���[��\ �!vGt��6�	�4���T1�يc��^�퍫�jP=!JEY+d��5����R���%|��G�42��^
"���	|�ߎp��uw�sCa`��i��6e'�`$y�Bk���d��S���8m���?���BϪ�%\N.��`R~ߏ��l6���Y4ޘ����!" ����ş��������������sU�N���>$?���rJ��6.�Hk��Y�	�Уǹ��,_���1ky� z�U�3�g+.��}Ar�mIA�\٨�D��2��m� ��Iq�L��DU�H�2Y�Scxa���k��B �<ldi ��!k7���c��[�x��.��q��î�����m�sl*��SԊ�U���� ���f��.�����d���`Bk.�^��N���A���%��:��W-�{l��a)�zm��~�πj��ش^�����n\[�k��?���#����J�����ڎ��D����;�Db�Պ�]}y*���P�|4�O����N>�p{���y����)<ze
M�oG@{�
%-��ͩ7�\\��ݯn�`���\贒�E%w��=Pps�����3�@y�=p��@Y���_7,���������ʷ��o0��AO4d�����Au�V�����xc�`����5�=��r�?���c�z�����j��`u=����=���6�B�w+��%���vX��=1��e�:&�l��o�y���=y~C�V�5�ދ�������2�iB43�A��[7���X7$Ҧ(dZd��|��hEQ}��<�^$y g�1Z�;%"��Ķ��o���!�����x܂�9{J����qQ.<Q�ӅV�B"�!
���� �ͳ`�H��C��쬒1Zu�N�է�[M���-����?�O?��O}P]�����6~FFFFz5 �:8�:�����u�?��?�ƿ���>�����fng0�M�H�;p
_�S�;]J(Z��=fZ,&�����Q����U����Y.�e&H�Y���:���ŭ@|'���H�t�)�h��h ���:�C����4ԯ��,?�N��\���OҮ`�Q�� �b0�S���F�
w��.e��{s���~�IfF�;O������8�A�4z�;���._����)�s����(�g._�y�ؑ��|>A/u���ޫ��O�i� .L|��GS�~���sdv���<�]y�^���._�T�PL���h�b�1���~�� �  �ܿ�݃[��_�( �P�TT��܃(�'F���5M� �����	<py>Z���U~��_�FU��V�L��a�5��p͔M^b���8t��~#�NuI�ܥ<�aÇƘ�r�����cY����s'���<r8��H��@�X�����-�g�Dk^Cc��X	�GH��"ނ #�p�1���h�������[!�������H�F��9��<I*N�	x'4� �(?O2U�fpb_{���'��{:����Ϫ�n  ddd�� ���̼|�V������_��f������+j���gK�w�#z���++I�H��s	k�4�x��C?a�9�;&����r���&���l�f����i�Pު�}/@�}.�� ��JS�
.*Ii��k�:��C}�!�$Z�I4~j\О7����j��G�)���������n�JZ����������)��Ɖ'��.'�p��2�\ĵW�S�����|=���%̯�_�yQ}w�L.ܼ+���KU�����M��:�;{m.�Sx#���:a8��$����e���일�2�ә��\~N��f�[,�p������^���������;�x���Z���k'ް��7ނ���dddddddddd��� �S���Mȶ����r�#����r��o��( l�5���2Z�����8���2 p�DQ����^����(�#3��:_Te8����D�hv�BJ��ܖ���S0�-`��������W�|2ѳ'��đ�%��l.##c�� ���e_��W���z��Uf�"�X�I�|���eY��ƞ��=�Y�aX�Bt����;�H�a�H�h�ŏV]�}���uB?�X�h`ɻ?*�ҖTFJ�K���ˮ4OA$����]$��)���]���O�	G�ZCi$ ����,8� [�-/D=�[0n`�7�l�ﻱ]u�F���j��ת�j���yV[]�6���W;�K6�z2�̛�#5�Z��ڲ�.eu�ݓ��\���>ٗV��ʿ5_Vɠ����6-o��w��RYn���NN\<��+o���y�?{�h��:��G��Ǿ3�N�eCD�ɬ�����	̯O�B����Y	e������x�M4*p�������p&�p�T����+�7��uz�xσA3Ea G{��uR	벒�m%���	<2���xc Gο����0\H�"�Ǒ����Yu�%��W�p{�	\䀫���m=��|��S�&hT�r�����U��5��nW�{�Ӭ��
V�u��[�{�]��q�2���e���YI2gsԯ����6_����m��t*q���.ت�������Z�F�n��]��^by�]����=�����=�*�v�s��	k9�hZ��O�u;(j���Q\���j���E����M�?�0�}�ۊ���.͗q���;o���iQ ���GK\~��6P"�4F�����5��ъ�@��Q��B�D����|
ա4�[Y堜ܔ0��}R�����V3J�8###�C ��OO߽~��/������/����,�7ag�gP�?�i�dt�c�Z��<��芳���H6'�$[�I��"�)���~܃���6(5ٹc�������&��w�ߓ����h�аpF��;y� �0xM)������r+ ynɢN(�(S�?�2�*��$��mxK�q�
/�w��A���� �#�j���zx8���������^�:�����n^��.4�K���(�&>:���k�B��nl�0����t�Ճ_�q��寞�0�Ƈ��Q^?�������+���m��Y2��1޴���d�ᴺ_A�9�}�����7����f��`8O}�Ղ�rɞ�<��>w��E�ޣ���\�k7�rF.@��3�pF��8�$;��z|���AX��9�ҒAF7��;####�����&�k��{��a�tL�f�5>��V�V�Y��S͓&�_߸	����0u<��I��'WL4�V�ܩ
��m�Izv:t�1c-�����޽�G~����Q��Ǿ�f�hC�B�f@'T�eEP��sL�=!Ć̍ ��"8GN�_E�[(7S[��}�⻿�3󹚝��`
9
@FF�J�j `-������������������˩���*3�P��I�׼�Q �iY^uY����ϱ�X���^�2S!;i`�ɫ����%I���+����P(J.���Ѻˠ�b��2.*:��IY��R���A[4h�P$R�VgZ%���C�%.��hշ��X�> %�J��8�e�`|�����*ؒ,�l�b����f�7�8q����CFƱ�XރU臄.��Ӗ���٧ڳ�1~�a�#�� '8֞L0����_%r���G�	8/~Gk?��������ϧJ�p�;���0���Ly�����4=�+w�E����4��ML���0�duzV��� g�t
�~�@k�}!�����*Nh+ w��\�����xv��Q�����J�Y�pos?�/ҵ�N�C2u����CY+׽�����q�ϯ����ߡ�g��Om��+"_��U����N���׆o yv*T-c���/�ʯ=��ݗP>����q�݈߲c#qCVl��4�
iDhKupd�e� ����1J X1��1/a Q;}B���RV1��g4~`��#Wk�&`x��}�g66�$O/u'3��la����������j����?�=�{��-`9V\FFFF� ���������y�<[|�\���ō��L�;xO�����*Dؾ�
���&���n�v@�S:��H�%�~C��ŀk��y;C�4��u)��o�P�-�0�7�.�~.����dQ��Y��k/���0)���pە�^�c�fh�V`� ������%��[3F�J>�lM����C>up��v���kB���Yu:�6���]���,�}oD3z��5A�=�nE�b���=�v}���^�!��)��T��t��@���w1����j��{�MM�z�{AS�{��R!�����:>��l�ϰ�6Kh\r[}�q�,2f���S7K:�PT_N��>�x΅�w^���/Fs5��1�����������Cڻ�M���5��i��L���U�߾�s������_��Du/J26�zY���7�v�/d�ݠK�=�e���s�:9o@���k�� �"��T�{�Tr�m�qU�������3�b�gI���c���I������>�=��u���C�����c�k��øm�9��e^^#l���r�T�v.��kl�������7�	ڭ3U�gq�o�u	�14;6R��9�	�3K(t��?E:&��E���9�p��)��%LߙWs�)\�����|H��-�\��	@[)���������-�U���'|;s2w#9�HŒc	�)č��,����n٨�e�y#�J�Mf�+�2l�56~"���z��~�������~���o��o=}���-dddd�@� �+�y��ً��+Ɣ��-�f�v2	�;f���NZ	���1,}:��]_��p*Ėx�,l��������������~�
�Q\"���B�3�Qiy�H �*�RW%��~��9\�S�;�8/S/�Zۛ<��A�U�pҴ]�6�p�Zsz��@���>#oCFFFFFF��Ȋ8��[F�H�O�
NN�0���N������J��&=\$�ɤ��&��tc{��Ny�����ĩ�#坼��J^�z�he"��{������ӂ$)ب��m 
�\Ë� ����-########��,�NJ���i�^�e�����%�����g�� �,��no4̾�!ܜ����X[�R.�����Q�Eѩ����b]6K�G6,�i���8c�N�B��r"����}��q�Q�	�����;�h�Oˇ0��������|�wQ �CFFF�
 ���pr6S�ʹ�X5S3�;�x;G��� kJ�=������0i�]m4@�v.�:ui�V��bz�-ڨ���=�z�^�.,��{��E���� ��� ���g��|\߾0~Q�,KX�Ŧ���iէ�k�0+5L���r�����y�V�}` � B�@�3�m���iT�"��X�� ��oV��e��	��s�n1�r�L�:Y��Ok���ȸ3�-��2#㸐���1V&M2��U��57��d ֞�=�U ���γ%_&���Y�4r�F��cퟚdE�QN8G�*�Qƪ�Uu�|%eL�u��Q�t&,��ck�7cl�����c[BA����-��JF���/�1>Vy����/,z�"#@-��(��r���D�3x~���ޘ� 9���7
�[��0���caqf�vR��0����VsS*ܴ��e5~�э٠2���S�����0�=i͏�=�4nI�1&�P3��HΠR�#[F)x~���^�� m����E5�0q�K���f���Q�]��g�dddd�� ���>b>���?{g��\�[�$܆������ƮW\$���l uw���W.���["�1o"��Bꘙ�!�ɫ�_�"�nL��ڸ���,����{��� [:����:���꺨�pQ��R^����J۹/�[�����z���b�-t�+J0j�*�܏�1���Yq�$�SbQ-���Ѩ@�|Z�t���<�p�kpV���E>�G��B9���i׼v��dǍM��5���F�ݟ�mr�4V���z�k��b=�>�K�y�ݣ���ؑ�}�G�D�w1���V�mN��#�]�Dz����W��ܮ*��1{�m�m��^���j�W�ϭ�Us�y�:�	��|��ɰ�v��q���*�������*�!ڰ��C���1�'d=A�f��=�w-��h�,z���g�eeԐC���l�x��A�^:��N�� ��ͳ.*⎛)������p�? uY@�`��)��8�	T��zM|�agC�cT�H�K�;+��������h����q;lP���4Q�@�^e���� l(�e���|t�B��u[8����>�����G��,��\�]zFF��m �:��ճW���'������[ja?�ϋ��\(��r뭞\�EEJ��~IN�}a U>Ix}`�?ZpQء���!]�y�IP��Ggds!Q:A�p�.܍;�,��F�*�����4�%,��������+���wU�ܵe�;VIމ�@��5����>oe�ֆ&�:n��.,����=�P`]�>�o_�cy�v��jԿv�}uf[`��c��`m�En���t�?���]��n�zp�E�>��N�5���wv}���d��v듄!������d��c#Ft�5ۗ�i/[�T�L$��FR��Q��G��Ŗ��y���ZCX��uR2IcR�SlW��H��A}=ny]n�2x���[������a�yzt��|ˇ)m��}ی�b�Qk���A'���lSP_��˻v�|� �t&�ǄÖ��վ[�vů~Q/+Y�<��|�+w�m��	��*UOD^+a +9���]Df��p��\��v�O�x~�|������T�q�H;��ة��=f�(O��Y���U����l��,��C ��ˍ9��a���y�Kk�q�����Y�O=dX?]����Qqi��������y1Qӫ�bq �`gddd,c� �b�^�ԏ����_��?�ܯ�s�/����cG�Ŏ�������C��j��q�g��� �t�Y�J����a4��>���U9��]J#�n�S��ߍ�d 	qR&	�)�x���
�+��Kxt���( ե������i,���8�qdT�̯���X"n� ��X���L�z�>95�TrOX��i�ָl7��}���{z�w�6k�c�6}��?�C���X��,܃������TmpܮK��w���@���Zd�?���
HË��]�l�-�����q�P�}���c�7w���Oϕ>��<�!I{��y�>r/	��,"Թ��� ��_M�*c��Nar[x.�tZ@9/���X��O@�vv����oC����#x����qҧaI����b쨖&*M�η��:�ܰ�N �Z�sYd�@[$����.�V8nI��O拏��拏�����<p���@FF��j Pu\�ut���Z�����������ճ/»�c�;���Β�bd�o&�����^�8�"P�υ��ry�{�Ĳ��U�Z��X@e�}%�����Rx�"JA ���/�gES�dU�zfmQ7LLg/��O��L�tq���p�^���)A�5���A���L�[��#%�w�("�[�nA^���1>Qtr���	�_i� �7�4,WT|K�vEߓ�;�l�u_����3������d�%l3;N�K��E�Σ���z���a�����>�N�����Zn��9�ý�]X������c+�^���rN�v��v����7�]��v{Ϸo+{��+a���_�]�{��=�d���g/����{svAs���� `��qe����i���{���~��:RCܟ��CC�#��q�eI�C���~-��`�]p �(�9&vR}P��aR�*4ة��＀�'p�L&SX���,4m��.�����z��x�����\��X�\��X��*�Vʼˁ�F�'R�F���ARFX׆L���0_CΥ%�VNV�J:}���O��_|o��/���f�����" ���܂�wt1�ڻ_~�y��IYN���I:o"=±�ԁHWa��h���r����/�}�!+/�k0�������>5xC��:�Ҕt-����m��[0��׀T�L�����VY)��&��BCa\����������G��[�%1ϟqQ��:~���)��6�r�"D#����M��1L�B=�"XR�gܕ����1nX�%������3򳚑�����!�Z���X��"��<a{�
����~�P�}n���;�Ap/��8�l�𜎲��� ��.m�L�����o�FVb��Bl�\捘� y���W?��lXP�s>����ɂ�h+�_ޖ �"N��;!��r�S8����mq}����U��>��_U�K����X�A &�Iq�����u~���cx���(Sހ�:PE��⾫@T;D"����ӝ�
{�{�)w^c�(W�} �8O���|���,�[>�6F&���;n���6����?�}tf������W�f�:{��,Fy`탾`NF�E��G%���v*��?��§"36�{9�|�0 �� ���H�Ty���t�sGm�-̙vL��z�4}��q���	�!<{�P�6쫎�,�:��~�x��!@Z�fddddt�6N�d[���=����2Ɓu/���i���{�^��]w@�XqL����΃�����3n��#G���n��t���Uz/~�8�a������ɉ��l��7�C�UAR�J�K<	9���n��+فS����c�&�Տuz����o���|X �d��2򟖶C�� M	8B���<!��nSx�bsǟ��vdddt�P ӧ��_�����O^�ݨ�P�O,($�#��C'ik{��	og��^�ZX�yV9����H \&m	�yD7v�A�rEjhXି(  Doz^=Ɓ����[��	���t�-0��E��Y����J���!���H���e˼�e�����/!�d�^�I�`�?�@B�{Yʽ�Q@�Qd��FHw�������P����)��Z5�Gc��=6�v+s���fv�+��U��nt��z}Աb��hGt����H���ߓrO�f�����3����{CR��%��>���c���Z�n[Cw��/�̙����*s�u�!��w���5V8�����K�r����;���E����5�?o����Rz���hع�xR��{o1�=���q�{�u�F��{EX��� �s�y���\P��җK��� 9��YKd����
��)�"M�`GW�\0��j��������w|�����d6��Lr������� �z�b�8��?�[o��O<���^�b^u�����.������<�C���X�JN�k/�av�l�L>����=0J *��������&��Xp9�;�;��m-`�wVn����+�7,�� SZ����$��D�G��������Eu�^��D����8h`�k����1n]��l=���+��#c3�S�ݫfnc����6�<Pϰ��_]֌����Gv����]�k_h��l-���.�U\�娮v��uUٝ1����n8ܾ` x_��d��8�g�a�z��gg<s����8�T�X&�S�=D����墈���.�����������I�~�f�q�5np���������c�T����  �&�E�BZ@�7��9���J)�[`�4��r�9�e0F���Q.��(���#��i�K�9q�ʜ?��ү��+�g�����K�wf ��p�dJFFƞ�w �__�~��_~��O�T,JЋ�mաM�eX1QP��߿�YL1��C�h�$��"B�x�>LJ��� Xi��"]wQ*Xo9��p>`�BM�k�b�(0k��{�#���z��W�XA��so�657�<��M0"@��p
��Q9���l��D~<}gI�2��d�x�R_*�`���1av��w6Fy@�6#�sJ����a�t�q�p������I>�C����C{�/����1�5cHo�������� �̌�V��q�m;$��>���=��2:�� #�%�CJ܎OoH�DK8�k�r� �;�Oc
�9>r(eh�e>�bمs����8�y�7��#/\a�Ep�g&��H}N�N�!ڀ*�۞s���w���sq���e������4x6b1.: :��D	sH~k ���� �&F�
c�c^�;��2n�[��/`^���W_�?���W_{�'��{O//�2222V`�- ���7}v������1S��CU�s�bB]o}��4M�׺����୯��*��RQ��+ �*��!�0O�W�=����?*����c�=�O�E���V1~X&F}�F	�f��z�[�^�u��4ET�#ʘۡ�����j���(�Vo��/֗�J�?|��3222222222��@4##c-l�3�,5�]ed���$3G����8����<�C�7�	��(/2�sn�_;�A��;�n������Q����ʚ`""3cC\�6�E���r��''�XW⢢w��Al�M��F)�� y=Z(hP��Kpn���gZ�ξ��/�|�����z5,####� �-o��>�=y�tf�y���դ꺬���8/{�{E�켍����:#��gR��z
�:w��M� K-i���}�T�Bd�<ѯ=��Ũ��}����2^1	k̘�o2|��tJ��5b�o���r�(�6
2J@Z�x,=�r���}�>ĺ3���|\�*R�L�t��G��g�׎i9��m��_ԇwB�����[w�{��p?�m�2���T_7��cm�ך�.����x�U�C��K���]�wkp��W���Fkr^�-����-����ժ76��ƪԚ�ץ�j�6����=��n���b��1���X��n�or7�������_�R��gl÷�|�1��|W�N㑮�~�s��{��H��ե�W�۴5]�\�oɶ-Ҟ`����_�.t�,�>�����ڻ�R�]��{����L�҇��?�k5����.��Z�;צ>T���\���}�^�V�է�����P(����[:�k#C��EENZ&�Ad?'���#-׶Gf��x�@`����1m8�o�����h\?�J�֣��@Y�.�|bz����'ʅ�����X�� \�e>���?��G�������JX1��M� �N�u�ы���iC5�.��������+
��;a"���2���NW���
���Jkj[�q�|�d��E$�U���d��&̤����-n��i9�*�t+ f�9�B: h#���:��Jl}�Mf`E*�����}�|��C�c��b��MN�ٻ�:��R��eЂmĢ�or��X�������������fdVX��F���"��ᡭ�kc������t'���a���k��:7���4o�����{���К��RVek�Y��o����[ q1!R4��[�*�(�'P0�B�{'&�[v�DGS����*D���C˭��"+[4z���9�ک���B�������߹}���c搇�k0�@�����w�����ٍ�-eP*��<�-DOu����eܻ>%ģR�d�T4���}W|'JD8��Vt��T8_ˊ"��|-�Ֆ4P�����P4!c!!�X 녚��m`˰�fVx�����N�}Ͽ��X�um�{��ʑ������i�)R�\?C���Ae�`�CǌCC^���󘑑�yЕ����q��f���vSIe����h��
�?"���;)2�/E�FnA�Brs�$���L� p*� ��O��a����m��&���v��� �4��g�Q��&ZKgI��<�H���!9���-���ޑ�ED�,��K��ͷ~�_��j������a2222j�� ��\L.���w�[_������/�o���ũz�LU�+
M
BCl_x�GK�HK���ĸC��]��Y� m=��ҔT�����AҖ���i+�L����	�6�����ORNd���|>*!���j��#!�$����2�GK�[�I+�(k����Q��6(u#>%�}��.�oZĪ�7�k�3���S�v��������0Х���i=(��o�(v�$�3��c�Z��t����m��697�ek�WdkG��o���O�fחa�.��k��,�]�Ǉd��l��=���\ئO��������=��tC{�_�)�㳻y=F������{���~χ�K<W^�������f��`�O�������v���}�>1�\����,���]S��^'�ř�T���F�n8��ΰ�+,�r��n��[��C�H�rl`W�ܼ����=��܅�x��~�v���H���r�I$ &�k5b_B5�{!H�(�I/"1c�hC����-�����]��t����h�`De�gf�D�<;}�}6o�$?�C0�沪7ߊ�!�,9LZgL0���b1�����ӳ'EQ\U'� 222֠W��s��Ӻ��y>Q�?�s?��o����w�������Tՙ;# �1����rWa�-�p�ZZ��T����C��t������|�1��EPT"�"�>gI�(TD�MGR�����<�58�#?*T2�n~�ފ ��N�L�KE*���rcK4�u]��m�}�y�PWu�<R+��hˣ7K� Z�Ǆ���1�|�i�C��ю��yD�������w�vlPбȶ/�~�֖&�\���l�ѥ]7n��� v�0,˳?d���,�e�RU��gB$k�6�?�|�Y�+� �w�HQ�m��z1f9g��?r*r��$�� b�����h�b�Q���W�[Sy�$��h`_�@�s����G����ǎ��;GKWN8.���rI� )��@SY�JYQ/�6:���.O#���$J�(�u�a��QB�������7�+Џ'����_@�!222�`� �x��R�{}=����~�Ѕ��*za��r6]ZvȤt�b��'c/Ih�����)a���[����dT ����� k1��v��>�O�W�K�z @���	�.Q!�N_~r���qm�LIi,o���<�L�,�6m�J�׷X��3_Y��ޚ�5Aj(#####ca��������ϣ��gd��=�o�3��/RN ��D��2?������~d���q�z�ԡ/yz���'��o�UD���W�gO���C��!Va�}�dK����H��QST#z���"��W��H9�`��޺9nE�r`�+:vFC��~�M��N0�Y�&�=O���7^[(ev�Z####�� �׿��گ���}vu���ҧ����� �����&�Zg�O�":Ğ�`d=��s�!��S@�1�?Y��#�ef|��c�H{_���W*�3'�z���M���B��r]$��T�X�?^��	Xf�h��'伭�H�n����[����r��F���ѯ�G� Y�����}[3%�q7g8�{ e�~߰�md��Y�ۂ�RT�������XmRQ75�� �[�]q�V�&�K�>)�M��q!߳��I�e��ln���,�s�����>36B��D�6G�]�dz�KL���E%��b^�����^$!
��oIsC���gb��)�N�g�A�-�8��y$�c[�3�ۺ�{������(�ȉ@�nc�<I*_���_�'0�M��	<wS}�vO����&v�W�ͪ�2222֡W �+F����+�[��?���كf�.�����m�����y�P���T���I�o��2����a�6��_\�(R4����X��4�aD�c���9:���:S�Ƈ�qו�JG��W�K�uu���mX9�����Ve >��rz&�e�~��uC55�?)t+C���@�%z�G�FVEe���|98.W���B��0�P��a7i8(�'5%�ɗ��P	3��#�#T��lk���$T�V�6�sw��m*���n�t<Fc.�X��l;#1��H��,�͡:�΋��#��Z�0��gt�^� .���-l���-���Q���ю���a�h�6�O�e����<6����5��� w��q1���ܸ��W��}�����^w���@��O �Ov@�>�y��=�%�B��A��##;!?�G]�H�68�/�m��ȭ�bcX�"q�5���j� ��w9��>s&XoC���FU�#iu̖��%]�����O��_��ѹ>?�L)� ##�CD P�,�]���g?�;������c&��!�	�O1�ɡg��ly�Ä���\���n��
�p����K-�?���*(��%h+RbBٱQ���\?L��a�&!o��u�����ߊ�v$�����x"�e#�2U5ُ���O6���T��`�'UhS(�������#�4��/HWy[p;9x���k�hG���1 �:��/�4���2�Ŋ�M$#�
ٍ��x7cИ��&����e������\�<��B���r�/*���X%˵3�����_+��}q�@]6^/	�_��O'�������Yn���fW٤�Ut�q2:B��� raZ���)�QPF'4���[�^%�,�FH��9�|p����Km�8�M�IZ��/��'��E�Qv�xE��$
�)�����s0��|�'l�86�0�-� ����Y���Y�d��E�
<௯��R���ͼDX	O"˴u��x���3��_`�Dj?ec9�Ӊ�$��y�� ���v��"9C�N>Vo?%Q��6̙T4.�v��zcQo�6�V�p,���ы���{�_�������W�'��J4{���dddd�@� ~����_?}���W���u�Sc��+� ᯋ��(^ɫ)� ��{ͣ�8��3dH�hYEU"K.K�)�xK+$�5��[8K1��6�N������*�:V���)���Ν=���Tb�Һ��x��kR٤F2,<����KY�{����,ۭ-!FP�U����+e�L�k7�����{_�q!Uy�ò��j�0�����|W�A]�����iQ#���°���( �Z4d��@v�i:`�������a!Z,�,�S#O�Y-���1�w����j_�V�S].F�S��s��ǲ�ת�:\�E�N�q�➎���J"�5ڍ��C�ztG��y���e�Db�9��bj�!����ݖ�?��<�c�d���kz��*�Ʈhb_��P֒��Zq�&`?���JbB5[����޴�M���\�����7��\�8Mr��cl[>��=�)¥6a���.Ms s_�����E�z�AW.��'U���T�|v��=Gtw���4GP��zlе.m��=�z���.秼V`񸏪��Ǣ
a��scl3'oK��>|_}Ow��R����0��*��m>O خ]]������}�r�c�ej�xV	�����vl��Q��׮M!�,�@�i�5�����>�j۬����=�4��k�a��g�Y�Ͽjmª�ٖ��C�uj���# 7]9 ���&O�ebmMA�ɍ�4S=�lP������,Q��ԻY���L���Z���`��N�*l��D������Bw�1F�'^р��)+���T���\�����b^��<���o��o_�����i��E�7�����@���g����<2�r�N
(�&��
�4e5�/(y$����OC��,�8~�N�;kJAY��(.�� ��t �S%��\|� e� �-
8{[�`T��:*��.2Z�p�_��S,�;#Ӥ�L�:-Z�5��e�[�{�|�x��*OV�5�2�st�O��M�?fނ���⚌%h�T.-��&#���v�Λ�1��s���������=�q�T<���e��\�&�{�:�GU�y|�M�f'$}�JuU2���/��`%ҵ�`���A�k Q t�ؠ+�B�|^k�-�ض"��1㱁4
�儅3ƲY���y�ge_��+��`�@�B�6�X�N�S>OF��H���F�<A����:��td�B��V�)��8p`��z��U�UO���V�d0B�T0������5Ď�5DX^C����j�IY�]�y����Bp��0�%��B<��~�q���������8Ml��xl�v|�}�cggE-����	i�%΅�ak%υ�V��1W�_v[X��X��	c����.'�_������:l����q�1� �t~n\^�w�?1��1��a:+��Ƒ��᭿@��@����>Z��"�k�h	�x����'`:Z���aK��}�@PjQ�h�L��^ى33!� {������] �������k��A{9��/�U?��Q�EY+a%��,���]�^m\��#�t=�V�@��Hu�zmvM�FS�gh"O��/Tz�W5�{pw�zj���^�6&�=vi��}]H�Ԟۘ%�m���b����إݮ�ğ�T��P�Hj��ؚ<�s8l��+��l\4U��c�r�'�����}~��د���l�вڱ?�p? ék2�QX\�-c��� �s�����`pa)"H���~��]��/`yҴ@D�p���-��
i Qƺ�m�����{�u��s�er�".�>W��=�,Ӱ�#�P�ע֨�l�u�1>{��ii�@>��n�~��������׎Ew6�Y"�Aʕ��}^{�k�<��dDVzX͘��˫�������,	k%�GDG@^/�t ����p���{��ِS�!>�16���܏ �zEʐ��E��`>cpKfv\����T0�<PI u����(Ӽ���ʭ�Y@�X�l�L� F�&��k�꿉+������N����������Uo�C �o��'�o���o���wo�W���=,v�>�^�t�2�}TFQI)���s���g��<1�U�&,¨���
�$����.<H�F��P�J���XǠ�thc�`�������� MF �\q������?��^�Ҹ�.���CZ7�`xX����=\�ڼy��H��H�x�yJ��Ӫ��4^�ю��V��P߿�ez�d"�dt���"4�Q�m��� 	������=/�Z_ྰgO���GMǇ�5���@�ǎh	��uݫ*#���#��� ~V��1(?��C���������!����H����5�2�`���C5�dtBb�N�q݀�	���
�e���k�e�5�<�?�D��uԌhY7�R����N����$>$ĺ�
��b �F��^���}��(,�p�����,Ty�L�&�܈gEI+,=D�5���cL�\��5�$��lxN���^8�`Ɂ�qK��g��ه���'�����ë�bqIH錌��e�m �z+sV�]�؟���>����W�0�0ښ��\��w����Rh��?��
�n¹��P�D@[�����$E�a������vJ�D��\����a{A�S9����BT��@lw�vIA�V��n2X��m�P�e�D{	ݘ'���z���:|:�ѐA ��c����b ��M����Pې(c-���-���us����r_�%6��C��fP�OM�16��r�m�-��J��lW�&Ķ��p<�y\��zY]��w��C&	�,ߎX!WU�s�<a3��q����j��n�=V��3,ɘ,�� ���ù胕�k�٥sY�ݰf1c5l2VZ�/V�2�m�/��Wh���P���%�x� u�sҘ�o��C�eͨA�mh��h����}�B9������rM��"��;�*�M�	|�緔�5��IU���l���?���o|䃩��.//o  ddd�� �d2y���/�ԟ��/�w��?|[	�,�7r&�)����e�2ׇ%���@���&��B#��"r�����P/���d:�����,�w��?�&t��+.*�k��J-dK�B�:�0�ʦ��\��s9��2 z���������q�sR���\8_ܞ�[}��.�dDq���	)��hA��ŐXe�1�!r�ӎ��^�zkG[�j�4=���(�U��~�ޥ�ޕ����թ��N��p����B��������l���q�2���v�ʽel�H�,�����"s���������rw`�vo�}��~�M���}�m�]�륷�ܻ��~���9m=D��e�R�.n��M?rW�vX��G��'���<c?H��M�~<��?�w����\B㴘!���0���3����Q��&O��G�����m� }c�:uN���d�4x 'NW�^�_�7q��ȱ��Ȉ8~ĥ+��bn��������'���Z�gUg PBFFF�
�j Pul�uz���������O�������}�\�7UF��"���#�]�$�!#)�v�N`���<�Y���xl2��N����D�W��b�� D�1Pl��LY�s��c�M��GO��p!dЈ@E�BA�"��Kk2!��i�\Sc�vŽ<��[��h�3��+���14GM��a����58��v���m��k���K�> �gk�C�v�%B�s�Z�~���vlr��Q�y��V�����V����(|�we�`�?K;#��l�\��za��"��v!OY���L�.�b�/�����t�V�y׋�}���z`�Y��Z��s������z6x�N�x����x�w��.��}��G��o�m�^��mL���}����T~�w�ns�m��&��?#�b,�یiw���k;��]�~��~�&c����1���U�w����O�70W��sDfy��=g�'��I>~:�@c�e�}��1R�W1D�k�Ȁ	��'�}x�F���CJTH�J�DΆ���T�Ψ�f�zW�)M��;�\o�y��t���=�1�y���<�;x��C/�q{b�qu����d�?##���  ��n���<�}�������k��4J�B9�o�aN|��s�h���Cz����,�q2��H�[eI���)�ُ�!b �t=v֔n�{U��G�!c��"��K%E�ˠPE���N��-@@T~�dX9E"�W8c�� ���\���ʆ��:��O�� ���Fi���x�v�?���Uao6�&��9t߈|0v�wt���M$]�M�F���0�6��]�3�ep����6H�x��/>a�2Ԋ�C�aǢU�x_��k�G�'���{�q�0Dg��	v�ed�c���}�~�Q��K;�0F�p�uZ�1�����]߳�d=��|����z���k��z�5c#[��2��L�K�A��Rȍ���&�y<�O^ܪO8nŇ�7}��`�����L��5�#	r����`ZC-�c��.0b4 я�LS��zM-���,���!���X����=������vq{���߷�|l���������h�  �'�����������%[��v�M�ѻ�Y0�N|��I��ߖh \�������[�a��{?f�ץ�-�,͊#X���,L�c��a/i���|]8D��V�YH�+e������T�[K#J�hP!�0����E_����,VTKr�o]���82@��f�e���/�0�z�s�D�.��+I��k�}�k]��oh�i��=��y���~��yF�1#�/[!��g�og;lA,9�&#��<��!\�H�N�
�6,� �C�@&�Ƽ��H�s�a�{�� 7em8�\��2�y$�C� 0X.;��hϊ��t���H`N9'���m.���`���WO&�xz��ţ˹ֳ��0�cYu���!z5 �dNu;�=�>�����_�o�wj.n]�袰8)��^��
��Hݬ�|8J�*l 
� 0z ���
1i�z���f�Ll֏���*�՚�Vb��	�5^>���G=Z�I# *��?���`�9�+�ȶ�Jن�i(hDR_kA�B�`YΡ>
Ĉd=v��}�^�]��;�HYვgF�1�����3��/�P��4���	�=?\do��*�>�}_e���3�|����}��g�/��yS[��/�~�h���=:[rDey,�<�k��\�ޟ���5m���u	|��8B�І� ��!�D�s�_Qd5 �A��_��C1sJ�?���"9�XA[�ʹ���> Yp:���o%\��ӟ�������/�G�}ǧ������ ddd�� ���O����u��#O�������PL14K�kEE++dw$*{��d�O�r"�Yp%}�
��ZzE��R��t�'J�^��o
#p:H������6v�"-�9S�f�Ԭ� *�D.�]2�� ��B��=|�5_�_�� ��]8	�nOE+���l�섭���]4���l�!�w��f|>V.����1<�X���)2�1�g!###########c#䵢�0��z��x�i}���_&�W��ڄ/�ǩ�G��A�D��In�OP�ԣ��������6k�1�2s5
R��s2��M1υ0_�x'OE�V�1:�lo*k�l�$��\�
�oa���S�85�'��G�W����_V��<z���� 222Zѷ�v���b~�a[^�P�|Q�es��'5Ŏ��>E�H�3�,-�����넸�{� �bJ����I�~³D�BG�F!�>�\�`�eI?a g8Ph�gƁ� ��1tM��ʄ������V�k]�D�HK����i2\h�A��\z���2����u���<��ݗ����}$��T����_FG�<�i��t�����1޳��v?��~n����egddddddddddddddd����2�Pw��ݢ�ȭ��#aSU���\_U��i�_�,��AN&�pE�B�*���0O�T@D�<�B%��1�B)����Gh�������̫v)(u9�g��t��K_�ڃ7����pU��!###�CD PO�~���ͤ�M���F���ٓBF𗀧�E;O"˃�=��a��y�俴Sm
#t��o)/E�F�t$��Bq�:����h��sI�݃w��lQf��`C�ڌ쿼�A3w_ko�_�-z�7�[�B8���9�R�� ��%� ¹R�?'G. ���$JFFFFFFFFFFFFFFFFFFFFF�`P	nk瘠V���n�俼�_A^��l�T<9���L�78>��i��_iKr�4��W�9�=Җ9R*9k<Kqa��]�w�42h����S8z�1���"a�Ԥj�-.-F��/^L�%5���)����!###c5�0 �x��!����u,�DϠԦ�Đ�.
�sc��U�8T$�U��@�u�ʁ��lH�JT���-%Ϲ�ޒ̑�U����}8����������V`6�z�6�K����M(Qa%RI�К��!�vO}>צ��ܚ�B���i�v�W��M Aɱ��l���>]X�/y+t�n�B�i	2�穭}v���m�t�e���CWq�����LfB_�?c��[�뚱�审
���6�r�~b��{Kl|�{B�>ch#ͽ��]ߕ�+����7���=oE~�W#������0�pw`���k�}��,�]�]p�7�h �O_������M띾-k�w���|U=��������X@|6ɰ�p�@=��R4�ڃb(L�E�(��)/Q��裨(��nL����Y�4yړC"�ˑ�`gѦ�������ZP�d޺:x�'N���_Fl�4�g�����B `�,\���NԹ�̷|2�����} �>��ط���w|�����������7�Ӫ_�إ����@�ҨdX��,b')�� ��V	�a�ao~������.�*&x͋���m	��dF���7G�D����]���b�/ �q� {��"��~c�C����!�?�&��O��V/y�.x��d��q�h{�}��r���{8ƹV}�a�u_�!�*���M>c����Ƈ1�-�_�垏�u��^�`,��X�Q�X땑�	�s�����1zH���iF�(`���ZӖ ���������x�^��S�j6�VG���� >!� �[��O/Z�ԓ�\��=)��Up��>� rI��K��6KN&5Xj�崲��%�g�z��/�{����������kFFFF3�� `�����?�����������;W��u��?�
C�ЅFk.�׊�,z�������u�$7�|��rؗEǽ_B�}D �Q�$�I���L�� ؙ�Y�WBT��TW���ŝy��V	巊hE�m�֑���ؚ��ҠR��v���K�����mKv4��Z{�s��Wܾn�c[±#, J
rcY8(����K�
��`$DB�-cp�PDx8![��ݾ}�����{�9��U�Ys͵�\Ͻ��5��Yk�G�k�Q�c�-O��,��2���+U�T�R�J�*U�T�R�J�*U�T�R�����_���t�gVa�8�1�|-�w�:{�%l'�b4#�0� ^���@���^qpg0����8�Z��q'�(�D�0("��hB�8� �j�`1.��(���G#*�/�~���/���#/����_\�O�<y��@�J�6�Q zF�A�����������ӿ�������U�o���ZS���y�`�z�aÞ�H��g����A ��1>&���ƫ][|�Y4.�& FH�^� A�t|v��&g� �����,X}�������>����=%�ɟ�ٸ�$=G���|Y`�o�g���FL��Al�����i���O��a�V��|�zuwq�އN�&����e���񼯻���8�u��+Z�O`�Q�k�:���ۺ#�E~�9�H��
ùI�N��dW�wF��84��d���Aε�8O=��$wFeي�<':�y~�|���9��}�u��y��
Ǡ]t�C��X�;v��vaȧXnKS�Ҕ5�yz���r⾍�m�!�s���o�^�o�7�S�.#���J��(cA|�3~C[}	k�V��)��ہ��4b�h.�h]��$L�� �eM����Y�E���?GkS= �I'�?;�&GT��K���������������7�I�M���@�J�6�)" ��bq���[_~��o����z��u��Ɠ{	�'{���@����|��6͑9�����n��H�?bA�霤S2.�W�0���|�K�i����w��@tk��g�X��Y2Sih��mZ��Y�>�k�=��\�ԑ5�[���C�C�}n�)e�wM{����m^i=�2ަ�e>f�g��Ǟ�8�*U�T�R�J�*U�T�R�JwC�xB1��qn�yzMta�Ԭ �5(���l%Z;	@�����8 ��������D�b�oz_��";s�ɑ�#�1v4(`�{c ��F�GSنGKs���i�sRl���CMl.�n�2�����l����A�1�T��:�@bp.t7�?����/��t�D׸��z�=4�/�U�[�h�����#c ���#�ǿ=��h��$]/@:���ӳ���w6N�y�%��H8�x���;��X/�S�eY�B���0��#Hy�B���j�I@�l�W�G"�]��:�H�*��Ԅsj�sQc�N#�h�u���l�m�:'/�]�ˏ����9�yt�t.s{Hc����NXC�c��]Q{���֕��}��P���J�*U�T��NdAy�6�E/����C�c���`�_�o�FΌ�b
��Dc808F��̟�A��A�ےdl)e��HG�(0��W�:k�3iƈ�6\2 ��78��K�D�����9n�� 0P:�3�o��n�J�*U�H'1 h�fvss���W�y}	���;4o�x��S�������0m�yb��(L5��hɅ� �����8̀SF�!`�2��Ǽ�?�PH��}s�I3�S�����2 �� ��W��� �Q �H��{����-��/���������e���+��i�mh�����b�ұP���87�ݶ��>�òoj�%�4�yttqh(��K���m=�֎���>��ܩ/OL��c��1�uя$3Nn,�Kb�jy�����C[�ѯ%��.���4�<��T��
���2�i�s�牎2w�p���a�cw�~��*�X�|
��}�~�x徴y!u��0�����X\�J��u�&��F��#��^zz��$�X�5����Q0L�sޤQ|E�%;t:�G	�c=����~���3���FĴ��9�>n����C<*�)`=<�<���vS\
!� hAФ ��Iv�o��]���5��������߿�܏����Ţ������ �T��tT��n�gJO~����/��������lႏ>f+���=2Ht�W`?�кL��JC k!�j�<�=�lUftj P7SN��P.�<��>��`QM�	�&ˠx��T��?��*A\
����o	�����E��>�^�4�����e��	�� E�08��)����py��>=��=T]�������!�Ƕ���^��t���\�U��}�s�O�Z�J�*U�T�R�H���eǨu�۰��B{�8�N ��_��! t��>����>:��o���1���l��Μ@� ��>�e��s�8�F
gFVo*�gV\����F0�AXY��x�O��뺐��k}��~�/|n������~�����T�R��t� � ෮?|�7����=�/��nó��"st�3g�8��bf�VR���U�e�x��H{`-���3�� |��)�[\)X�aY|�4���A�6Py%C/b�\ ��{��I�����F4 �PP��3�^�]A}5���*�E�F�=P{��ʲs�/�m���c0�`ҁJ�O�0@>5��o���r��-�S�}�t�mbiJ�<���P�a��龕���xɹӹ��]�͛�V�s�:ϧS�秣�V�s�:�+U:,UU��H��� �W�9�7�u�{Й���Y�ތ���(�3�ɑ_��� Y^#��#x�o�
���<,و@0��`T�i�1���GWSٌS&c)��>�.}��+������?�C���9�/�y�[�F �*UZC�8��|�鼅�:X��3�y���q5� @�-f�� ۫@a��
'�
��	,5��%����$|??+����8a�r; M��j�	>� �s��k0�aϗC�۫C���3g���Z��*�kL��v+�W��u�$ȣ�5��L?��O�(-��wj9v�c[7�5)MHj�f�yؔw��5[����oϦN1�& �g�C��9�X`��ۗζMOMێ�sm��[w�t.]p4���q�h�r�y^�@t.]��<�r�w\��|=�� {\t.���3ǹίc�c��.��>v����h��?��8�ۡ���e�ɋ��b�b"'g<�@ygp��g�� c(C�=��96F ql��|����#c!?�F�kƫj"D>B:_�g�Κx4@�N K9�H8�+���JQ:�w���y����K�E?��3�+U�T��) ��o|���M�]��󳞛-f�#-����<{�P�8?�����b:>��g�����;?I���t�w��Z|�e�y''!� 7�EW�W�1�<�K�z���X~d�d0��F=`���P���ͯ�سeXq���)��z>禥����R�J�*U�T�R�J�*U�T�R�J�*U�t0Zg�0t�~,�^/���<�)�����/d	�/'�� "�h�����9@�p4�(�|��BR��~�.0�$
�H���T�i�!}�^��C+�4;J24�����v�^ݛ�<�$(�g�
�T�Ti-��  <���]<{����.\�=g��s�>B��G�&�T�
��⼔Pd���z@���G��##��S��<;� ��~.x��$o�Ay���dc�rH>�ECP([Ns@���x�(A��,�q3O��`X?*��MY`�B���>,�J�����T+���?R'��c���ۅ�}�ߖε\�И��{��]��X�m�|(���yn�In½�k����s�S��a���c�iJ~��N���H�*?�3�v</����cPm��:�+U�T��ٓ[qM���+���΋�#��=��>�P��_�Es�|'	a�~*Y4�?������3
ܻ1:��/��A�P٫�q��'�Jn����ыߩm��������w��>��Oy�A��$�w�q�sa��&^5ﵟy���{���m���mT�Ti�  1��GϏ���x��?����;�n^�tW�Ybq�e�>�5�����{\�]T�ϙG��@�գp��^�x �2m���	��"��EHP��d��� ��'�C���s-���< 6P �Ùg��<Fڿ�����+ߦ#�1���J;6��㠾|��4��������1�����NS�XyoM��oڎ׶������ܥ��݀���N�k�gS��:�gK�)e�P���sj���w���7_^������H繪7�Ӂ�f�Ut��b�th�ˡ���[�k���#����dϕ�<?=M/�w���c-��N�{���綥c����\�f?��i��pu�>��<l�@����[}_ǋu �ߗ�co�2��T&��̸c/��E����A�
�C��<h��SZ;r���C�̌i
��kQ�þ&� �f�ޅ %J&���a���/���?�s?{}���u۶���T�T�RI�� �͟��g��G��/����_������]w�cB��2qb�%�P�n=#���p��A��Og�$�=y�0Пs�*@8�>�})����x�=�3c�"s`˭�6
�VZ�f�Â*�ͫu��ix��8��
����F����+V�P��P������P(#p��n/�R%X�����R7��F��C��)�gjy�<�Kݏ1�i\��A�=��z?��<?z�}^i�C�?�C�c��J%�>�T�xT�W�J;R�p��J {�����5X��ȕ�����E�;��������'�9SCȻ�Ȁ��5 �¦�
�`'�!�#U�Nҗ�ѤA�9³���ҡ���i���g~�>y���O.����g�P *U����j �3��������x�[?�?������O��u|���8_@G :y�;��p"lhF0\�0��l�S߻���ouN7Z;,s�@����F���~"���BF��3��OS(�,[�-b<��Z��#VЍy�k�,����a$��6����	`!^F!��*��R۲�4�j���zU�O�n��α����q#sJ��ާ��sW���i����mꘞ��y��" f�O�J�E��k�v�tJ���n��{�J�*U�T�(��J��,9���zM��%EJ���Ʊ���
�n��}��h@݌ˀ���s�.rzx-926�(T��߀���3~bң�҈k��W���VZ��8K�PΦ�<��|���\����E�|�5����-<���J�*�N ��v������o���p�3��m�L�2���a�qu
�_�9מ������Y,!y��%�_�;�7���m�>}��]<�;`��l�EyF�)a����EE��o���?������_D;�>O }�#i`��}������ ���ގ[����_4���6o�fHؗQڔ�@�����ҝ�\��@	�ۋ�r�����ZnY�ÝJ��#���JS��﬊w��T]:�ۍ@Ώ�A��M�<?=�j�݃�E|�t��%݇���}��#m޸)7F�WF���<?�|�(��NW׼G2KJr�<:x4WkW�a���#gO��@n	>j@p"��A�(�J��|�;Ġ�I���p���G���>E��xIƣ{	xĵ�#�S�-��\;�i�q!��xV>�:8��]u�x�y��PZnT�T��(��  >�Y�¹�}�������{��:K%��6ZQ�ƈ���㠴0�B�{~�d�x���乯g��Ny�s�#��L�0M�#2�,���Q^>O���z���� *���`�S���J��/=�K����:��g�*	����6�":�$�B������ah���ް�*���IU��=}��=��}\�%N��}��+�.���(G%�x�G2��}{}�[�]ҡB
0�3����$wH�Hx��;v�N���ۻHk+���u4�\;�m��	���C=N��F�N�c��#��%{�y>���q�_YES˵�:pO��.	�y~�d���*�7���%�+U�tX:k�T�N���X���q	��2�ǟYe$d!=1������%�>���4��;��Ű:N.F
2a1���)�\9����GL��*�Q|t>?�#+F@c�.;�2n$X �Y�����@\Wt������v]\@�*U�4�Na �z���_�O��/~ϋ��O}�}2]r�Q�"8e�N9Xy���pc�f�T�0��Nd�z#�2�V����|�]2R o{ &�g���A����Q�ҿ.1���Q��fɖQ������Ͽ�)HPp��17"�c�+�5KO�od�h:�li!Xh����k�����1Uѿ?�m_M�9
�j\)�;|�Lq�y_i
�}}�?�w���P���9�<�&�s�}e�*>����I�e�!�t����/ȹ>�69=�y����y~:�<?��8%���c��w]�S��Ut�u�T�!й�J����э�/q��[뾰�~)�L~S���R����(����8�OT\���z,S~>��bƁ��θ�=�������!�BVG�>�Chk��D���Q$kj<k�i�>���M���N����K�s����>wy�����匚��J�*UZAG5 �1�+���˧�o��_��o�����gZ�UϹ�F��ߔ/����� ���
�3s�o*`l>��,�S8~@�0���t�y��( }6�"y�G�@�B @��¬Ř��(|r�H������})T�	Sc��F�I���)C!�F �b��!��<S��uEП��H�EX��wBkvN�T�I!�v�;���"�S��T�t�{�b�XWzwXﳘ���I�j��=������`�|��C��{���<%���g8�n�UV���V$|�f?�^r�tj�r�yn�/�Hk�m�nu��=�y�1��^z��N�B#۽b:w��ֶ�d����>��>3�������C�ɔ�S����M����������X�|�������<�w���uP/�1��|v��`�gV��8�/�%��a0��	�{p9��3�Aj���l98����ŒA�R|cE���^�g�ٶo6\�A�f��K�s���y�}��}���]�O����}�9��[�T�R�5t� �����'�7��Ͽvo��{��n����9-���0H�_
��}�3T��F7"�K9h`C�D�'�����Ѻ@UٺML�r
)�L
�Ҁ�M���H7�<��2������(<����C�$�00$�L%�@��c�9�,[G6L>���c�]� cT`_qZX� Eg���P�a;P�lA*U�T�R�J�*U�T�R�J�*U�T�R�J��c"�� ���������Ƹ5`�m#5���ޫ�q+�'J�J KIo�%�����G9:3d����4@�c�{�r�`C�����:	��G���N�\�Y"�GřBJ3օ�&�t��t�nv���>�ڳ��?�z����wށ�T�R�5tl�����w����-����_Ʈu�]�L�23�&���G��	�� 2�w_��gO���t�@׵��>d<_����<�sؖ�	�	�^�� F�+<��������=1����_�$=@���úp��T��P���Q=�����e��^�Ҧ_g��m�D 1�?����
 yP!U���IV���L����ܗ}�r_w������Q`���[=i`{�u��H}[�C�u��9F���n��Sϩ)�<�L��ٱ��.��%/{���Ximj�]�:W9x�o��%{䷎N݇�y��y�0���|]������ѹ��u�>�~�B�+OI��*Uz�T��'���?�p pde�������{�M�Pz�ۈ��А组�g�H�#���ẁ�z��ψ ~20�E8)�}��8�Fs@qL ;UF�7�Q��#Ep �%��؊8�}>�9�_��u�6>9O�c	�!ί���/�}�W��z�i�9��[�R�t� ��;߂'λhঽu����`�!���j9�`;���W�x�/���r>��l�&��A�xOw:Se! ��ѳA��!��w⍟(����� (0�X<[f�7{5f�,��� �=�W�Vg|�3�*m�n)���Y���P(�.}��-�P�R�J�*U�T�R�J�*U�T�R�J�*U�NQ@lޫ���oƉo�Rd���t'�C�  �EhR��|���D�6���GB����O�c��eZRX�h9w&/�.��#�����#��A�t��w��t􀖆�L=a#�"�U������ϻ�W�{����(�T�R�J%��  ^z�}��Y�ыڗ=�5s��K?��ǻ3�.3;g8�р�J�t#P�����r�9tL&�X3����H�`����x���G��G�<�p�_
i���sY89W�;��O�t F( *���DB����ah��wE9b!ۆ��0�?���cErN�]u����6	}�okבu⸒P�yǛ����pko���O�)���GhГ�0�����*ژ���6�R���1L ���{	��V6�='�2��7��h'/�S����Myn��If�㢽�늗�������	��N��P�燧:�'�Ђ��lj�=�y��Jh�1r������4�t,��O��` ��o��p����,�����;�y~:A�)�;����x�G�������7{�r\�R���(|�:$�i��4-���������	|' �A��`���5��8�b^	�A���^��9Ejh�51�Q�q)jO�dP@^��#8u*�#����8L;r.Ӄ\�M��m��,�|���?��_�^�T�R�)tl��ֺ��|���?�;_��}��ͫ�Õ��̻d%?*s��S��a���"c�3�1��Y�`V|	X��c�PXeQ8�,D 3u1,0��?d��(�l��;���pX� iF��C��Vl^��D�=��3X�Rp+��u�wI6:��5̰��$(�E�>�r��69,���s5�ݝ����z�>����So:�c0|c�a]Zw݇Ǡs��S��r��K�	�L��-kW��T��z:�<{n��]���J�����T�y�J�6Q塕Ι6�13�� � �W:�i8z �p�.�qc����C�*�6�1l~ �����K�B)S��@y\rv�%v����!�L�JN�
�k:��"�r�j�J���F'���)C�w���+���/��?�S�����[]wz�B�J�*��)" �g�g�������W���?ԅ[�G������,���#������J�k�m  ���g���J�x �=3p�|��ĸ��g#��r�6�Q�������H?��=���-߸�+h�3�<�&3.tJK��BmY0�c���g	�* |~�'!h���6�$�xU�V�8E�+hj�l[�	�K�]u���GM}_:\���R��~�l3kU&�iwM}Rr�ע~�����X����h|�.j~.r�Ҟ�vˤ�Pp�3dݳ�E\��N�����d�U��<?2ݳ�?�y~�<�|��;y^������{&o*� �����ؑ! �N�:N�͞��i�&�g��\y�1@X��������1�.f|� >�,�b6R?��d�i0�φr-���ёC��6.�RVПJS���9�j=�wG0��������;������Ͼx���o�龄gϮ� T�Ti� �g^11��mo.�Ň?�?����_���k��p�dWa�H��أ�6��z���;��b-�T�qZf�D,߂��Z�Ϛ|�~퉙�[(@�p�rF�f�)��7Fl���0̝� ��Z (�;������&����%��P�s.��"���srL=���b�B�ң҇�������䙜r�cj^˖�'���:3�=�"N���t��`���������vU��>Ϗ�''w@���}�θf���0i�6\�L:?�iޣy~��,��C���:ϧӔy~��v6�|j�[�ם�� ϗ�w.s��{,��u�I4l��P�Ut�e߅ց��F�m#��s�3*#BB���u :��0
�X��[r�3�2���^w��cpe�A5
��ر��j����7������B��O�s�Jf�G>;�4��?;9��8sr��䴜��U+�C8K�WJ��=��Ó��͗����s?O o�'��P�R�Jk� �����u���W��u/u�K���l=ꑔ1������DT�dϸ��g&4/~��/L�χA�w���k=]I�]R�<ɮ�E<��p����p�`����`�v���߇T>��ԋy�e�`����3�巇�C+�Ij��V{�C��.t��~�ʺ�V�e���sNm}Neن�-����C��P�}h�����]��]�+�R�}�z���P��9�C�����O=���9�}���Tt�y�K��������m龷c�J�6S�珂��u�����-B���l$�eC�e#�M8C���%��!�0��y�4������cW�A|��LLBc:��1�a@��C�R9�����6!����ψ�c~8�C	�0G4G:�9{�t,�Ze<�ӣ��~����.�1�s��:�q���}���� T�Ti#�� `>��޴�[��7����_,>n�k��W�v�W�zf����92�}�~�W(�7טc�E]%=�#��_��/�-ۇ����H�H:d��)�K��; ���ɶ�<�@(��(��M���=��6��b�,��uրl$Q$��v�<)���H؅,L1?�Ϡ��AcjBm��36,ޚ�5f�K���s��F�u9p�t���}sT9���8���C�ǩ���㠇������n�*U�T�l(���FX���MF �t=�����S�Ĝ
'L�`��g8�һ�&��R-��	��9:�,}�}���	_�`���q?2��b =��I>�>�EpEڋ�G
i0�"���j|����@�${�F��D�R��4��1^-��]b+���*U�4F'1 ��f�������k���������g����<Yc�Ȍ�@߆LaF�L�Z�	�"�`������)Z��0=�9\�A}:� k�s��@��g��"$P�ܳ!�)9ţe� ��z����3�Ie��/�{m-&�"�����0b�����A�݄\�e�cE��Vk[�w�չ���R��q��J��t���n������B�Q&$7^I�9�G%����;�V�ʹKޓ��&<�MFwS�.�֥��!p~<�y~NTts���u<��a;ܫM�A;��?�ir]wѷ�L���^��P��wLu��]Z��<?�
��~�y�%����v}�z�`��ĩ��]���o��v_t�;��t����ot�tM~���hϱs���.�!��D�Q`�������_��4��`L�-Π�,�\-���*k��Sd�%���'�W3h?p���c-�N��%_�b�G9�#�M��0�?97�����e|�	�N#]ШЂ|��ٹm[,�����/����Ο�7��;o_�.��B�ZW�T��
:�@Ds'�a������/}����_,^��p�����d)	M��3�#`���[�we�N��9d��9�ò� 996 sNd�ޖ�ė�g�2>�FC�w��l�EFl�����!�kF�n|�l� �������01x�`�웣
�ޛ
b�oJ]�`��/H� ,�|�K~�&
I|έ=/�R�iݞæg���n��Xk�}�r~�<6�3	�>"M�sJ�lK�^G��fp�h�}�ٷ��e��z�l��V�=��+��ZS��çIF��*U��T�y�J�*U:�$�^���=�#,���I��@� ��, ���#�mt ������tߖ-nBۧ~Eغ�fA��&�h�Wഀ"��qPf>b@�����xL�-(��9G >����qZl��BF K鹨=�_���m #Iӓ��������g���k�^|��������{�����o��ֻ���t^�J�*-ѱ# $V�|��7���o��/�����%�����g�w�?k0���c x_f�G(�������6��H"9� �|�V]�ޑa��hثD�b�	��r��	��_�*��7Nl��ג����j�Z��T�M�O:���vy���A�d���Z�j�*U�T�R�J�*U�T�R�J�*U�T�R�J+��]���� :2H�C(�iz�8����"�L?:`��䀘���bt�/ғ����ʲ7=���z&A$N�"�x�g��eC<"��'#L�� )�X���������W����f���y:{��_��o��o=��g�xo�}�*U���Nq�{�^7�x{Ջ�'��i�����z��p��6n����)�<�m����+�{�x��@��I!=	��,2�u}�	��@�}O���Y4"����=���pIr�C�|}�<��t�I����xL^ֻ?޷��mZ�}(�a��eQ�,��
�#7�&=#W�yTC!���m}#�����4��X3ĕ?��b_�}܀��߄���׵�U��q������Ne�[�m�l�5��m.r8�[͹z�l�i4�j���LqUZGǏa��ud�J��I<w(�
01�cM��M�J�Ou�o��V��y^�\����]�~8�	���ǰ��TtNe9%���Hr�<�Hx���8��Р��w�_K�?�t�/@��MD7V���-���L�$�f%d�~�Θ�!��{(�
 ,&.�Ho��&g0�T�� 2f�`Wz�@�N������8�j4��l�Y߷��OX�t��q�����Og}5 Uc�T��z:�@�u���h��8�����g����N ycC�{�o�:}s�YZ�u4&���)@�!�n�#����wM���y���h`o�@���� ��mr_��!b@�eC�5�|�?NCPm��W�7,���U�ƵeB�	߷��*�j��?�>R�Om�&�{�k�J��}�ct�˿�����3=�~~(��Bu�WږJ??�zL�:�+U�T����'�q��,nb�lo���k�Z~c���Z�cn��ޱ���uB�1ҳR\J� �c ����^��tL��2�H�.v�8�1ƈB�
�~Ŭ,f`�E�Q
N~f����N����y�߄g���yv�U�T��:�@x��~��Ͽ���ۯ�x�\����zg���L����;~G'k��L�˳]��wȐ��\=ЁB��O�^��\�"�����3] ���^�$ǲ�x�Av������~bC�dֈ`�ٿ.ܿ-ۺ�ՀB�6G�l8n_nG�̻ �.Ea '������k;l�ܾ�3��i_ ��:u�3�C�S�c�Ec�ٷ,�]��Hwj���]�p�q,��.��9x��]wY2�1:W�e�>����t��_7�븺���qӱ��:n�ݩ��J�*U�T�^Q�Vg���"��M��������/���o�{ז��Eq�n�2�0�4��[���@��+�^���>�$N�-`#��`\�*r$�F���ݒ����bFs44�S`P*�ĩ3�׻��)�4��d,���8�;�����(�u�B�E�G$�f���࢛��;����'n���/��i��~�\�R�JG7 HL��=_���?����������ʯ�W�a��x���-3z�ņJ��"Sq 0T"`� �37�̱ ���F\�������0���k�]�Λ�\.2"��B)rS�Ζn������EB����6Y����-�?���6X��C#�����/�=�.uLBQ�d��I�u��U6�������;MǪ�}����Cv1v�Ǻ�W�w
ڏc�m�'~5n��_z���<Ϸ��X�DG��^ɺѯH�6���b����:����X�:ϏHu��Ϊ0�#�i�$W��2�ϒ��ؾo�T�\�>͝�/+B��.@����p���� ��H 	��y�o����є���ǽFX�lX�ip�-�@X�S�?J7D��	g(T�<�˕��h�j@�b{GGA�f\E�&`=�1����$����g�ˢN����{Ƥ:J��&#���5dW��{s���~�����M����ٳ[ ��+U�Ti�N ���7�y����'��?�t��G��W�n�<��\�ߑ���(b��/�G9>c��aL��=��B`��g10��e��+(����,��6[{��`~�D迧_].�ox��X~i}bC�<�$G(�6*A���ZEE/Ч��e?��E�2JK7��JܷK}:�5�+�����D۶��Ѻ=��P�]���>���6��wn�%νM=���um}
�ڟwm۰��&����}�S�J��w�_+-Sձ7KF�qu^T��R�J�*U:SR���H���[�o�@
��G ��F �y�>]����|�0T4��\y�N�p�_ɛߡSgp���3�'�/Gɒ1�p�(�Pt�J�#9�nS��@B�����(g��BM�� >�A|@#��:�X�Q'�R��f�ޙ�u�3?��]�.>��}��X@��*U����j �3���7o^σ�'Mt�����|�筇[���֤/����!a����|���e�b�b�����Xe	�-^�@ ?�(��B���Nd���B�R�����#�ڲ�䲯��x�.�=�`�sH���eY�k�j��\n{\�X�Ya����EPv�so��?�zslLG���1i�v��6�D���]����m_��yp��]5oϝ�8�����حT��t��R�J�*U�T��(�q�i�����m����	��`q��� ,r�� ���b���:�`M��k~�.���D0��Q�ɰ�YD��4�B�C@�=_�Z��@�0���^ӕ���C�}JgJ��7GB�Rg/G�a��C��H\���5s%��D��x��������9|�4�K@��R�Jk� ��o���7��o\~��'�[�����eK�&�������:�F��0���i�XJ�+��똩�l�-�2'�zg��u�ߤ�_K�	%@L}鬚��jAc�m:&�g� �1���	T���c,"�xT����Ȇ�JLM{�����/e���-si��%�?���͡mr��]W�ߙ|a=��"��e���w=&6Ri�0R�Qљ�<`,G��\SC���F�ZS�a��|�ܛڎO����!��Js5�*���=�k����,���0�n�8"�r���W�ﭚ�K���)ƒ����Ҡ�a��\M&-��Z�8^&�]S��fj��*�AB�-'�ʱ�ϯ(�R�#d�)3��p</|��1�>�e1E��/��|�(�p��;��#�N���]��i\Fm.�[9F־U|���E�M�����mZE�Ԧ�.����|e��P�mo<7�cc1w�C0�~D]\����6ye���5u�����a+������~���7χ�'��!��Ϗ��>�vWc����y>���<����ڴ��g�<ϩn]�{:�7𴻛�C2���4�|�=������܆�+=]�Og�������<vYN��{�[3���c��<�����m�w8W�_��1�ssj�J6��&]m<����3ϧ��y>%��s|�u�y�ߗ�Y��Ҕ�X�O�U��|�@�ED��[��O )���hT � ���o �>]?�?Jb���ό�M��'Ϯ�����8�ͽH���a�Ep������9��`-�����sN��~.�3kf�H�����>B�dXh��v5�y�~i?-f�߹��S�}��h�9\�'�G�utP�R�J�$ ��^}�ճ����o�W�6��t�	Db�l�7[�yP���U����$PX�d@��g
�
�B�L�l��2�L�zN�O��d���җ-x^�j�^����A���8�t���g�����@)��S�5�@.uX��c�b�Xaq���С���|E�G�g��<�1�2�? t�ƢQҵ�s��1u�Ҹ>3u�e�����-M-��2�����m۷��Ӻ�<��8EǢ}���6<f�>ܷ}�}�܇yW\���>y�CqýS��}Қ*+W���ٷ}�чS�ǔ��˘��㎡�<>6|��u�C꥛��w�OMwUS�=�:�~�v�3�w��S��U�yh��t���X}~�y~�u�9��C�(����"���r/kS�۴϶rw��E�j�s)��韺S�z'菼'N�v���S����! ,nB�����o�~�޾����5���ݢ/B��}~�_;�I����Q���:����Q����C,br����f���}}!�H�>�Q��`�G/|̇]��FϦ�ӑ�M�Ѡ �=t�$��ѱ��>�p����҄� ����H �7;��S' bU�ԡ�2Ej��H�����ۢ�����>ro?y���޺��KO޵��T���Q ""���b��/�����?Z|���/n�u��1t�5
�p�@<�vWa����;���Wz�)�16]&:�Y��/���{
���ǥ�� q��'H�d�B, ��?�1��) Ƣ�B�k�h����?��1���-S��� �O��L;;�xȠ1
6O��!uR8#R9R{'�\��4�i���Q�,�zŦ�܆��"E�&�V��N*;+6�h����^���e�쫮����$:��}�~:P�k�)�+��̋}�����x]*�)T���Mxfx_^�f�9�>�=7Ρ�鶓E�}g,����-x�ػ�1��g}'?{�y��.��yf�<���.�����9����� ����lϩshM[�?���,��a���E���x��צ;�Q��yzn�����k�w��,�k��y�X��[������_��Oy~�Ϗ�N�\k�م$�Yyyj�1�W�;�G�,����4��w�9���<�G/�'�}d���N��V�<�<�ri��6I�H�P����<��ջt����cc[��Z�3�<l���8�� ����l����n���P�|U�ۇ��L[���{��[o��g��_�t-{�����/ p�����+� ����-_�}���t�p�����ql�����k��SP(~N��}bYJ6ȅ���9�ca`�M��+��t���`��(/��F*D�^��	1uK��(J����P$���o���ֿ��������~�O}�������?p��c *U���N�������������]��;!vٝ>��!_��nIrǁ ��@�>�<�J32L
��l���%O�Y��c��Vv\J	��_��ʂ�-��z>:��g��1?�1CTy)���r��T�R ~]� ��>c��1� ���Oy���~�ٯF���>�2��Xh&A�+�M�mO�ۂ���δ�W����q�rC?N�ow�|<�]�m��u{�I��S�wW.>�&{������V�}۱{8�m�d��ƭ��w�13|7�ih�&��q��tyu���S�C��]�:ܷ��ՇS��T�U�צ;QG9��s�9q8:�^����z�~i��<?V�m�cv�>5�C�}�>��|{�7�C�����~���cf5 t�<8�������G����LI�����(�v<q�;���������	���n�С��!��>�o��z�r�;*s�z�ӟ�b����x�dϜ����-FH��o>�~�,�}� #���|���Kό�s_>S�/��*��!�%����t�<��5O�r�rd��A�ބ��| -��������8�5��N������51Eՙ3�@5�y��c��/������݋w�������o�}�*U����m �9�7���yn��x���,Eh⦉�ye��9M�͕��	��&t���&��s�ų]M 
�_f[2oz-�:�5o��qT� PH�)Jf���$P<G7p��c�^��>ò����c�y�F�|d��l�|��7��&P`�8L��ؠ׿o�q��p�T�T�R�J�*U�T�R�J�*U�T�R�J��l��O�������E�n� �1�A �_܀���y�����>¸�2��8@�[���gƍ�T��s�H�|�9]2F�\��W 0>c>[2��)�:kF�8{�|7E�8�2F!�����qӶ����� W�K�L�^�x�����ߗ�m��=��맟|��U���VE�*U�Dt� 7�����]67��G�tm.z�Q;���{�c(�X��h �5%_ ��#����z�m��+���; <��1	����ϑ,�P *@�G/�Edoo�Y� ɖ`!	?���d�#�^�9�M=K!Ŵ����s�
֫@���hz[�T~*�FC��h� ��4���D�_�F���*U�T�R�J�*U�T�R�J�*U�T遐�!a1��"@6 ��Z�����8�Ő��m�K���h������y� ��D# #^BGgp��8�c��
 �9)�?�P(�>{-��9Z25��H3�H��@׵* ��ry����&�[��,���s�������Q'�%֒"��ϟ^�?���.����\���!:�R�J�Na ���~�;ߵ��ˏoCxb�%K���x�= (�{f	r֋�1�4 ˖U��W�����D��a@2�r���J@��x�K����7��*P_���ty��fș{6�L	��U���%Zi�^��{�4�o<���U �;�|�A��BA���jz�'r@av�Us蛘�u��<)E��l��[o7��{\�=7{~��yS�{6w�o�.�K����f<��٘�h?ncۧ5�e����lP�81`Y>ZB˝����V<�p~����ѸKXɐ�C����(^�Ʈ�}el���(�Q��fV���Ge9s�d��s�� z��1��L��b�ȟ��ؿqi�����ƛ�y�z� IC,)�wh�)�.��j�1��vԦ1�	�Xx��K��҇�v^�R��q�R�)���-/����?`�|���ϴ8�4���i�1T�)��|2������6�j���/�q���!����pk=�c��͘�r�p�1��u�!-
�y����H��N<��D�ڣ^�T���xy��h'��筵��7sڛw�W�l��sB�(/��9����miN�sE��?5�rkߧ25��l�h��Ϸ[S��ːM2VK^ZUS�Hn��}N��AP�<�GQ���5��۔��͋eq~?��(�~YN'�MK�V'�YNj�x3��U�[�T�ہ�*������|��ަ����1��猕J��,�
��)϶�S�c���enZMx��9�7G��}���������?�!i[�<o��mG��8�F�����ˆ�N"Gy�uLg����c�I`~�m�mD�E�3�V�\�X�{ˏ�N\+�3���# mrT,~_#`i��e��r>�@2��2��O�t�|b��yH�9~�r�ȸ3)�rq;��`Yx��,_�<�5����8^#��!?�2+oyz��g���8���Q��s��,'6�4���_�����d(��1�I�U'�+˫������(�1��IdD�m��u�5�f^�̳���'+�S�w9opl����:��C�g$Ӹo��۲$%O�����H�ըL?������p�緺���h��W�F*��'�*��(˩s>��2�o�q�� ��������;�����?]ð��Wa�U�g�y]$�幈��t>o�{�`�p�S�L�t�)�e��g�+K���5�{L?e�59?�kx�3��N�qPG~�t��\m��PhY��:k���7�K��϶�]J�c������1d����[��{ls>��l',��t�b���6虆ڌ�E����X���p�i���3��@׼ôt�0�)vlZ���o�y	���c�/R�L^F�2�q������Y��^�V�r�qE�C)Ϝ�嬮)��v<��:�f-���<��:�����/��0塃��d>l�L��}���Q�&y��,��7�?�k�r�.���+6�bP���:(�2�͖uSS�ģ� �������v^�:�?��A��y�C�g9_���ɺ@�/�yA�:����Fg�k_�:��,�x��p����~��H���A^ddZQ� �*�(�uoP=�ZG��G�.�}����]ޓ���T�B6��x�Ǯ�CG���=s�fL�9��&G@�o#�Ĵ�n��uWO��M���+x���>��x���\\��J�|�m����ej9^����_#�S���ߝD���f���>y�ayN.�;�to�^7 ;z�i9]�3_/���e2s��uj�sn0.��+q�/�m�O��H�ו�� B3�`�0c
x�c��[�z�r��ٖ)�,���/����'�4��6����|q#gS�W�T��) �;O�m������kwݤ}�;Ps0VB"ƻ1�R��� B!��V&V���m��b	餍�.��n��J�s�P�7���	x�%��O�O�"�� "@tW*�C҅�.�ݸ!Lc���8�pQ�M��`���A��5C�J��r_�%��~��"+W�~�j��v������|��>��'��3�i1��ݬ��ŵ3Tx���c,o����3)g���lH������Rz�IYq���,���q٤�H_� 즂.eg@�P7t� ���b(+m���|�����t�T�@�`��r#���n�F3����xCG�,����gR�x��?�4��*Iy9\�"ȍJR΋�~�ا��]wK��א����q��e�PP��墔>�>^���/�@����"i�!�H��?yq�KO֦��F�P�O�S:
��3��2+��S���_}�8�2a����T��(�*�҈C6�3�py."��u�-G�t�F�������4��#��u.�����삗J��L�x#�9c�%��d�`y|^�������O< :�@3�B�;����f3H�u��i ص9��	\�B4Å�1��m�ld2oZ�{?����(B8I�ps澠E~�e}H��i.{�͇�a�f���nR[y��S��M9SiR���9�VF���W��*h��q|�����'x���ܟ������Y6I������k�"	�I`p���2���3O�2�%�HD�@+Q�~�1�|<Glٲ�@F^��1��J<��h��&HZ�"=�ߠ���8�(3�c�x���φ@��Mn�̃��& �A�|I6��������@� ��"(��6�IY�b���J��*��)�gA��K'�d��/�}:�RwQx��(CQ~c�qĮ<�i��ռ�ɼ�`�K��>f���Ug�>X���Ƌ#��(Y_ܾ�)v��ȝ���x��������J΍��ƨ"��)�0:��rc��D��ö4zG#գ@�&0���@F&�O��F�,t�R2�y���a�x��|M�nc��(���&�eJ����L�~ar�:�]� �H��9�a�cb�����a]��(b9��PB���4Hl��Ei_P>K���ԇC�6K���d���_��q�X&�3h�|Ц�cZ�7���o�^%='�9���+��u�����7\â��("��c�)k$�����F��B<W�h����4?|P�:g$�U�������s_�	��u�y�tf>�Y��5a@�}H�a�-�?��v�FHe�H1�u��O�
|h�������2���`�I��$����c6<?�n����ض])��?̳��x3�R��5?����2<�E��8pXf�Lۓ�S}��Oj�ٌ�&J_$�n���&�9F��8��W�kF2�c,ד��I�� ��ѕd�H7��p~V�����?���27E����F9M�(���U�kI�FiO �y\˜*���l,����������{α.�KB�
�D�gR�%}���S�C~�<\ew����Q�<�>��`=ÀH".T�)���[�����v��iʞ���QZ��2h;��,5�>�;�?R}D�)�iS��Q�G^S��O1?7�#��2��1�G��x���e�P֋nẘ�1��h+���,���Z��cY�
y˺7�E�MI����X���y�g�A���ԙb?��>�c�Q���Б<�_���O��a9�c��9��5�k!?�}����s��G�9���>�Y�ލ�;y.��9/��s�)tJ�C�{�'���ΕB�'^���۴o�2;�_�3���m/�9<�����O��M�ל˸����e�uX/O��otF3>���~��W���.�����κ�җ��@��%C]@����n!�T�z��$���)S��&�G���y����<� r��5�Y,k���,��e����ƿy~J��O��֤�7���0�y?�.���͇.��?��ڷ��}����*U�Tұ �
���������w>�裯����}_���X!���Qg�^��b�@��w͢�\�w-Vk�!p錄�gtUE�6�͛a���
�����DyS�tS����K
����fA�u^����p�|����Y~�y&���X���K�,�l}���寬g��ic�W�r��<��ԀI�zho"|��[��i���.`vշ�E�˙�i�<�SݢW<vJ��E�lI�q�r�v��M5�8N��b�ѸC� +sQ7��^r�m����E,���y��Đƴ����b��I�,�R���vee�,�S�X^L{�8h;4&���d�Xṛ7,e3D��zT�e.E���X���7o좺�ސ񑼭�-@���x�=��xn4�����:����O�z9�ꏴh�?:Y({��h�"o��A�f�h�Ehd����`xM$�8+����B�A�E�'~�̚�1�^���B�e�����%���ݜ�ŷz����Li���7S:or�Z�BUo�y�[�^q��!L٠�c!uÎڛ��~����ě�M��i�  k�:�#�*h��?����&PT7m���Mހ�}ܡQ����1�'�� �~���oc��z��7g:3�K�tqGTn<�����E?��ü^�3o���f�v8?�?�Fkc"o�f{���-E��%^'sQ�8��c��G��"Ϭ���)��`ɳ�U�w�!�ZQ�D�A�I��(+J/a|\�;�>x��c!Rp~����Dc4W796t<\�"8�]����z��4��\As� .6��\��%�A>�Qx�o񜖍#Ӯ���?8Ǒ��H� E�9�<9Z��b�Ւ�o� �� 8uчU?�zk##���V7�<����Զ)� t1�U��c[Zd,�=d���GNG�����Pw05���#h��`�E�7"�H��72u�up�_�3��m��S�# �FEl�bs�s�4��%��ot�+8"��r��Fpg�ГG�%�Y�m����906`{ܖ���g�Ob�H��D���r���k��Ϲ,����cи �{��(G�J���+q���6G��j��\���:vc��D����]fl<b�7�]���54�S8V֓P=s���Q�Ɖ܊4/��9�K�dg�%�0Z�DL�q����f��ź�k2jd�E�G�+������z�3"}�G�X��S>��j��XNOm��J��xRP�e���a�6Q�� Fz\��w5V�ց��,y~�4�]4�$����x_2�te��pұ��2>ӽvъ���Y/#0ߓ��<1�fى. N����
ߍj�&����Bg���u<�$�X}!�6ku=e(벍�74f�M�y�N�����<3[ғY_�4�~�n��A���+C	(�²A��x��(�� �_Ҹ��,������z�=>գI����Bg�S���Xۋ�K){� �I���s$�/�g���u���u�KQ�,}�M*۶P:�=�����[���>��W6d�F��:��4�[��@�������3�9A::�v��m���s,�0%^��$�N<��2"�վ�}��_��(D77<��Ҽ�����t92e����yȺ��3��V��x�M-����p�����/�xe���Se��?���9��?T���8�u�t%`�f��x���^�<7Ĩ7�/N��y��z����E�m3�!c5f��́F�Qғ50螢�����C5bпr]��+F�3��<y�5��0�����됨QA�l1TC��e-�u彎�x?�sFrQ�V�>�С����85F1��Gu�NM�#b�}8�İ��)�Q[.��{	.�z9���5���-|��O������%�+�N�N ����v��y���j�Lbu�e>q�}�!���b�!|O���=Z�����ף^(TZ�Sf�e��J��kJ$��ht���
�5Ⰱ��(�?��y���-���~A"%"�93�-�[������������>ݗϞ=� ���T�R�:�@��b��l����������׾�_}���iX�Є�(\��
�j�B�pz�����.�SFe�fZ��}N��xV����(^"���`���``���P�%�,�R��!H�Bu�����nqݬ�W>�>#m�ͤ� Y!⦳i�g�5�(����|9)m�=Zv�5v�-0_�xWo9x�6�;��`��Ș{ �ha�����Q�x#K�M���ۖ\ �S�W�7�lX����O덖ƺQ�@7����ݰe��Y��1b7�!o�$`P���/ru�>Rۦt�^��Ji9,?Z��LJ���Z���*T��j��F�n�������Y�f��
�|��.Oc���9�0��X<~�!/n� C2��g"Ђ�#)��Q	`��	/V�Z�s\
�-�639̴.,��r�s�� $����rE�^)k����9n��ι@m��&$%��3���-�;G���Ĝ�*�@[���t��^��G,����i���&]:���7+"��iP�=��א%9�eKy;הs�7m���ow42����_c��?/*9=��Y�FQ<V\
q�`E�0�c9�M>�}��ʋF�M6�JQ�LA~:cq��㎫l\�X�̋l�>.��N�6vȀJc���q2�Mu1EFn2�冥:���s��#�p1����o.o���G���x�F�/�A�(��{HX�F��Ţ?��4��rLH~7�$��3�(�|9l��q�mS�n���k�*�� N�J��9�=�6��}o!�'	z]P(��I�{�A L�X���;NB�.�d#,�,�e�WzO1���;�%4\�q�t����\A̋�����I��%�aB}1Á夜���f3��ʿ ��'�'��xfK�}S<�� �Oi�O1�r� 8��R�s��o���T�6a� �U�!8��?�w�����Pc!�u�<�ō�俀@`�=Ƃ�D����y�1>T���K�"�����䶢���l#�	���"+P��9?��� P��p̲ x�S4���|�j,�e!�Ε<���zRs�ܗ9��6R_=�:Z1�f�54�:��2g|!���9�[ͩ�T}̩�d&M^W�~�s(˧Tv��l�b��t�����"��X�'P��N�xlq��rIy��Gd'|(� ۙ7����'5rM�={�i/�2�y>��$k*݀���m�F*E���S��Sf��φ��<C9��<6;^�0_H�H�0���鬏8��BT���
�Mn�˖(u��2��j��.D�Rӑ7xz��&o�glC<!��.�2\0$���Z�P�Șu2����k�e��X���/IX{֕DhD�Q��E�������R;6�3SS�-�t�Zy�2��H��S�;H�E!D�&f��xPgٽ��(}���}�p^��PĨh�7�>̗2%��;���t\_C����B�A�s��	6�hd-K2��'���e�F@��6�uu��%S�-�]4>�6��:�H����cH��k�v�����S���B�����ֈ^�U.:�����������p$,'�J��C�I�ul4�'y}XY�fT�\��=q�@�cž�����G�b�nX��Tz�ǂ�B���\�u_�'�a�@XF5��Qb��h@���e�<�kb��jD����h,�=���)�}�� �f�a�T�rn����90�#��&Ov��*wIy���_�� �>w�;(❐u?m �A�y�]G�ͬҰ��{8X�Vv��������9S�F��eF96\1��%#�P<��>x͕[�{���Z���]���s���1{��8zAs�˩c+�Vp�����AK�Q�DrNpy�$���-(�W���+EZ�z�ʹ~f�^c�p�6q��y����R����2�}�n��t/�����p�:�7�;�~<����)�7g|tcQ��{t��I0UYl���]�{ێ�u��Q������ɾc���2?�hB�������L�h气�V��\������5���Q�Sڑ�s��6Q#Q�ԑI��ZW'��Cݓ�FG���%��(�߽z��������|�Q�����AV�T�����^�&i�ڻ�˛on/��㫘0��(u��JL4L��|J6���&��BY%s�*	}d��-��F#�t#0/ꌗ��8�ěBXGT6�B�����rB�� �*�����:��΋ �f���;f�@�_*q�8F���K�ev����g�Zy�g�6aT���o�����M�)���T�&[�g�߈��@�&���޼����z	o�}��.����b��I��x7G%�73p�m<�q�bŦ��CcEE{\�j<r�S�Hx�>��sGB�I8IZ�D2F�͆4�j^�fkiG�Hy'%�,W�q2^�z��b�I���ǳ������Bz
���mԻQ�|�oq�iS�s�@�h���Q2	0�g�ݎ���(���jS�`����pͣ�D�4�yT�N�UC�!.Ӣ|�VI�S�^�(�� Z ��t�D�n�7��2�ً�x�i�D��� 7z��׃;A���C��E�	��ޣ�0/u l��,���F~F���
>h��0�ܧf�E�V=�	�q:>�=���8����<�-��O6���ܳ���<�n��e�ח�pl�_:_y���|֦z*S�e�ј�["�#����b=@��\Tm�6Ƣ7�F<�^�z��m�8�ӱ�!/m��B͜O�9t!o�	x�;d��P��y�/.o,�r<v�o����z��d��E� �r��fkx� ��r\�.5b>Fc�Z�[ ��`��%��=,^ ̅�BX7�����<�%ҌS@݂B�Q�4�ې{(��h��,T`�P���<�*/�,|��5��SO3�(p�DX1J�lp �� n��ác�a�fS��nPu	$w�dnJj8\ԧ�R})�]��K�< ��̍�$b����A����[�Oe����<^EF8/x��ж�H�ATDN����#c��K���pN����z�ҡ�m��fET�3�g��� �A7{D ��2�Bg��\�Z$Zð\ֱ`+Άo�n�1���a~d�|�S.�׾���D{�/�4V�P�|��3z_6:xF��5F5<[xM�"o�:�HZF���z�1��<���*3Y��<>T�u�xf/ ��YiC�+_��\u������1GRY}<�k@�*�>��9!ۧ �ս���7���O�V�b����_���y�kS�fw�MCj�;���̑���f?���k������%�H��Z��L�{��"Eq��_��àzp��h��|���x���E�M�1���2p����k�	��h���)�����3��w� 5}�d���}S��Ag3F������1:S��F�SDǻ���Ǳ!����Ǔ�S�Rړ�(��(2W���rP����ԩq�3lD�G\p8��ά���vب Dҝ��b����5ς&ض�z�hȏ���'�^��ϙ��x4c��]��ٱ��1���,��ĵ�u��]��O9��#�� ��otO-�xo�	0�Ķ�t8�Ug�я����H�Q0���T9�e�qNPx����Y��yH�ae/�ݸ?X�0�@�A~_�gS�5է��/Y��}��������Dur}HG�+^�Y�b���v��Y�6e22��#���y��<L�"��	��yE�����W��?T����CX�d_�dQ��4�g���A�XW��Ƣ���~��e�5����O������(*��6���5��Ȏw֝�"��Ƽ�"�ʹ�<9��:L�m��k�92kj��,I�]Ku��Ca���Όړ����Τ(Od^���EX oJ�]�''��W�����D�~���i�{M����H��/��g�r{)�oybٽ�/�>1Ry,L��Y�##`ym"?rͦe�E
V�}[/kH����դ,��b6�r�?g#r
��c����j�k����I�cK��y�2����"��C�I��h�,�W���$\_�H��[�D��"z7���zĬ���뫛��ޗ>i��0���R�J�� I��K�������{ow�O 3:�����'e�48P!�1��n4 ��FJ6-\p��,�p^T���7�P6��:VIr�Ez����sy#��0��+�C��w[a�.T|�Q��@b(x�͋��{�B�ې�4K?(H\��*�s�L�TPx!��m��H��k�9������ yC2=�+x�E�}�H��,)�	&�����bu����A�!� 袋�'gXS8a�`�u~^�ifڗ�+���l���Zt9x��or����+q�I���LW���R��A�.�#��}�}�~'E�|�H�F�VC�K�����Z�v\s��!˱xV�� 6��x�B�o�'��ta`Ɯo��'�>��T� �+f���`_{]E�B7Ǳ�go��AB�;Z(�1|Vӷy4����M�B�,����.*ƞeo���۴'��ʸqjٿQ�g�8�OK<vX�D|o�/!�L=�y��7i$4en#��O� @�z�0VHa;����v�h ����Gn���&��vi���N%>g����=��`ٻ���eC7d��g��B���+[���������vI����=g���1���8(�"Y|E	�rAr�@�����@��!��A\ Ad�ĒŇ-ǖ{�3��9��^O����U������;x���9�^�Y�tWWW�WWW��iMp���y����X��i�d�8yu	'���2���}���+�𤑒��is�ϏD5��,v}a���5��;Én0h8$T�l-dI���E�]"m;�̧T�l�OAw_7�3 4'��S�O��0�fx��iq����x ��W�<>*�W��9��)P��6,Q�MD&v*��y�|��\M�R���m�����L��g8�7k@H�z �t!�B�˼y�ҸZ���ϴI>����)A�^�~t�:!}�������5��9��Ԩp����8H�t]��;�y�kEƺ���f��	��E�gW�/6`9��A����)�+Ng|�y}�����/H�T�w[�ʷ��"�o8�@����h����x���R�M�����nT"�ek�+��ST;/�\�iw���,�=��t������ym���䁴���ىІ9�˳����,ø^��Z�����g`���Yې��������_��m�	g�
�SF ���`�e�����r(���W���[���K�fq�;6�/�A�`��s \o�-(l��܎8l
�i��+��'w�2m��!׮��R:h�'�ߠ��$� �q
�m�6;t�K�d��Q���B��٠�BlTq�c���� 8�ģ���#�'��-�gW�|%:S��<z�Ñ6�u���2!@��^ֶF)�Ր�nܡ{���>�߷.Cv��9U�F���^�ӕ~|�)��d~ٲm�6�����ݑ��t�i����N3;ސ]��#��N[�um���m�u������Y�L�K�x��1׻��R؋+�d}��6ի�lT^�}躬R�x�8��T��zO���뿙�1���f�'�}�`�u��j��V�W{?a���N�#�����\/�l}3�
�n�)�����c�,s||e��%8��IV�<a��}����v�y_�xN���eb����fy����|�{�����J�]�V�%d`Օ=?�V�����A�67������h��{��D��x�_���?���&�1�G�G�����A?׬��:<�oFֱ��cS��M�K���C>���/4�<�16��Ӛ�uq'���liw�1<�m����B��5U��UBߦ��#�sK(����������q@(�����X��b/IL/!���h�ÐݶoA�ްawSp>��?��}��v�����\��3�ꥼ���Rn�/" ��z���_���w��K_�n��K�n�lc�c��=�7*W?N_D4����V����GG� �Fvto��gD������4t
����v���u0P��0j�C�������
9-PTŅaM�����B4���w(c��
�D��b�)`E��=�F�@�ޭ�_˥=�'���}���_��ܱqV��wjo>��0���I��Pr=�� � b�l�B��v�h
��{l>����Pz����+JI����ɀqD��F�E�v<N�W>�lp�1��d��
�J�R����k=�ǋ���i��ԍ1���i��ĖW�� ����a���4������4�d�8T��(GF����ݝ#�yAt@��js\��ޕ�8�F�7 ���������f�X#���k��D�8n6o�л�m6&e��w����l�RBі0����wl��9 �8DJ�6�	7�H��i��s����i,')�:'�j�f'sŲiĽ���2�.�û�&g�j@��D�����=�ER�@6��9�׮��x�4q��8�l�c<`y=�^�C�aM�#�7k�I���Y��e�K�st���u^�©�N~Ž�X���c�fx�+���\<(.����ǋ�E��洏��0,E�/�]�p#�6�!�'� CH�������]�lc���	�wQ[`��,��Y�H�����[�Ǧ���D���p�Rȓ͍_3淬����z���l������{�e4�����22���[���!?�D'�����uH��6:ݦ��4�͑൱��pa'�U��v'N5�Z\d���dGj����{�m�Y���ψ954�@�G�9��1fǯo(l��L�0e�z}p3xܵ�Y/L�p�؃���{Ж$|E�c�OA �]���W"cсØc=��l���UB��n!s��
��(����A��+z�����cۜ��M�e�7�RM\0��)�!�`�w�#ܻt��F�@��t���0�t��k�(��WЦ���#�U�\y�aЕf��FM��&�B�lsG���|�{ӵ�nqj� 4��m���ϡ�bM�����٢څ�QG��6���.잮V|��s�-W�X&N��S<3��)��/�2�u���	�ӺѶd
�ŏ�Gv��z�K��F-2ǐ=tߢ]Z��q��N���]�A�n6o�]�����t�M1�A�g���e���y�_�'���t��P{l�\h���Q��!o4]>x������Ax۽S��Q�sώ�.���+�:d��y�����m?�<�u�t!?���:�y��=�����Ʌ��N�7��?6lb��ql��i���u�W��}�\bE/�K#��h��]?�\�@��43B�f��C���.�����ʥ=�~�#��|�I��\v_��7ׇ�ˀ�o�%��1f<��@����u�X7 �ܿ��A�Mx��y���8�-A/Tz�#�����])������K�w#3dy�Y�|KϸkTς\8+�[���l��!�k�htZx�D@��A�t�$�~��0�&��B.f>�A���l�<ٻ���1#0���oC�C��
fP���.j#u�{m,�a35��&UO���Kw?����A�%�KЮ�όd9O�_��{(;M�o*�)|p��BN�ؐ���7�G��ǂ�,h�D�C��F��^F��i�N^o�Q���Mk��y^�2Mp �<YT�����v>��R�z���w��~!3�׉� O��Co����6�Gt�;��x��v�1`�M���d0�����3�]���@�[
�I���U���ś�j  ��IDAT�t��{i��l��)���������_��������/|�Ko/�?��!������R~��4 �[έ?z������[��o~��?�G��zyb�##���a0�K��}(x,3�R�g� �(��)�0~X��3�؃�F�E��*w%{��w�%4`q��SRL��ņ/e�8ּ���?���Ve ~47����M�n���q��a����+p�``%)���0V4�]}�����u��ƥ��t1{�?�Cody�m<���~��vg��	���5>vR<�Έq�Tr��p\k{B�/��֐+�ǝT�qvld�1�3��w*Н�c���L�`A`8���5�6��H�~%���<F��~�GS>С<[�Nt�ckv� <lt�%j8*D8b6R�Aє�n�:�cm���k��ʑӆ%�����ؑ�L���#֌�~����c�u�l@v��q|��׫��F���;xG�/R��u��y����Y�	���h.I�Yr�;�px�.�����b;��Tl����p�$#)�����ˠWK�-�*8�N�Xk���/��ԻE���o&a�/�6l;�xo�E�d���߻�~m�FN&��l+�b�i�l�#�BS-����؍����}�NN�I(�(��~кq/����(1��Z;��1߻7��N������bwt���p.(����H׺] ,���S��г���ns1hNFs� HЌ=�C�O��Ƹ��^��2ߖ�Ӵ��ͮU��mffw�w�����"yl>I
Z��0ir{�I��f��Q��a(����߀�����!��t�)�#��<'��;�1�����9Z��,X��Y2lL�#���9o�� uhG����BD����F6����;��,-Wj
��e��M�����q6o� 5����J��b���\�\\��.���Bi{̗ӧ�-
�Ӵ-�x�?��5͛��#���P����׊S��i3�w�^3=����T��#=�9�(��g�sK���d�fGbv>';��N7����K�"���i�I�����g_�}|#^tR .T�P�sY�������\6�$�ӽ}���3u12\g����l�{1�jB渢؉7�(�G<YQk� �>���@�^������<�Ty��lp��T�F��}��b�]��#m0m��r"��[8Z�
���S����.�v���+��KM�]�u��gۄ��z��2�q7����n&��nɶ9����u�kc��c3�gQ[��ta��ƻ�t�1�h������i=>������@c��v�;�7y������s�.���>���2t�������pu	~ >+]� pl����7�ۺ���D_v��Q�n4a�9Hǀ��]'u��bW%`~�@�sF�!E�1�Qi�Z���x�+S?Ƒ������W��alt �5M���ۻl� N�,�u�����ưxSL��i� T�>ǜ��������md�K%�R��6����H��r�@�4�;H7l���=�z��C;o�P0p���O�lXz+��@0w��۫��Ơ�=t%�)f�:v����n�Bo�.�r.�8�D�X�G�2:���l�Hǚn4!��<�N�y�+v_C�Q��5�#���-�h�&:���?n�T��5�ҹzO��1G�B_˚��`2U�N1�F���_=���OcY�\��o�<hk&�$�L�{s~�،Ϧ�z1/Ot_!x�����Lه�M�n����`199�^��XQW�� ����A?�����W�+H-KCd3�\ڜ�2�� ��c�s,�%o�s����gg��_�p��L��c�s�cDl�k��sI�	���ld4�^�E}��ۄ��Z#�f=P cu.#�5�u7�G����ɸ�s~9�lsC��E���T�V�`�˓,��|����������������|��q�ģ�H���R^�K��Ed �~�~�����𣟾��c�_�Mx�we'���v��K1�ٔ ܍b<U�LCX2��N��i��t�6�8� nbj���	�,X��
�:䦐b�C��:)�͕� ���p�!Ջ��s$�,�Q����х>���m�~���'`�!�����Կ85�e��Q�::��a@o~?-������wS(�ݭ�!�;�5=�M�.�lĆw���g�h���xd���C3,!3o�)��C$�c��p���6N?���|���I�0�^�[�i���S�ݰ�&F�j�'�)�ad�dDW�]�F������a%mSe}�\(m��Q��H�)��������2
G�����n��-��~��� H�W��)v
�A���y��B����-D�8�ʋ8M�Y���A6�c�l8%~'T�w�,��e���n;6�Z��k�y���<*��a3['���/�b8�׺+�����<����p�����6�b�ļ:e��jw�n���48�C�u�G�� �Q�{L����x�@ftl�c�(�x�5hf�H��v���8�Dsj������V��w��.a}N�B4�Z��$9fw�3����bG���|�|ΝѨ[��A�d�i�~@/N���z<�g�Hq/��!Q�����ej����l [J��m"��&�U`��E"���5�*�#JO�B��u��Jˬ�S�Me��@�V�LS��ѥ���m�.@R�c����<ؤ�	m��Ϗ��2��G��c���TܱY4�$�u�A|>��������թ�:���H�u�����kv�A��d������:u�������XW�:�:�,8GXF��{��2���kCl�!�X�O܏��3��6��T�f�wIXb�i�Vk}[��?"	oNW���M�]�t\:6�!���~��$�=*=�k���Lc�+?�OB/���si�?<uvO���� �0�2�̂^� �j����պ��Ѧ+<��V�x�����SP�G�
S���v���-t�w��Eа
�'�t�_�ís�f������H�e����k3N�D3.�l���ּ]�cu��T™��F� �%NeR ��<l\�ߢ��?�`-�S��9J�?6pQO��k����0��|N��Q�Y���]7�U}��F�u7�鉇�lh]$�?�}��8�f���p�\-��CL]�	J#���tI�%tX����ç�4ڬ�>A�'㗱v��c���ϒ�X^�\֫
��%O7(sْ�����%�K��O�D����l��t�xLi��:�kd	�NToi�+t	jsG'Z_+<�����H�=ڠ�!q]���z�		�F��7����!�c�K.�v�/bt/���D�`���H&]��8
���5?|��R
�C�+u��6R�v��P8j�,1�*���O��{!����a�!�ഉ�\=,��w���CQ9
_g�4(;��� �D�6�����T��PxDeF-�C��G3� .O�l��@�5Ք��֙2<�N���QD+B=��O�޳��mPa����u�[�I�c��M������z�],�֐��l3ca��Ma�&q��]�uM�@W06���80���vZ_']q�#L6w.���~�%s���,���ܔf��l�y5_/��{�籮|L��NA�̟�������NO�/!�����{�������ڇfAg�ڻX@
���ߦ��<�����_�}�G��?�w~�����׾�����|p�o�g�^�Ky)/%�t ����������|�>�굽}}���^�����H&��`x|B<��`,� P�aL�q��B�R7f%R�y�Omc�"��p{���$'Ct@	+w�Q��=�Z��|U��6��p�s(�Y���{���N�	�?���"�?��z�^9�����uz?�:a�~�{�Ӥ;N�0 ��~�Th���Q����g��͢�A(�oG*�fA���`Ш��?BRV�;a�/�#��/��m���� {l�݋�(\�����pb����)׈|�~�95%0��q->0�x�R��4������aw������PV����u
���6��t���%7�L��{�_n[76Z|���k+ki8��T��?��밎06�ĕg�	���W��b�j��8��sO�AϙKs<��;�b:i�c�K������Θ=U#[ h���)��cȋS�⎬����z<�Qޒs����o�4�M$|��U�Xj`̙�莧���D;y�bmPz�eDN��Cm L�!o��P]�;�v0?�Y�؃�a/��Z��;2UF��8m)�|�f+6ʝ��,<,�7�������-�#U$�!�<`�&�hM�6�ؐ�'�w_�pVZp+�O_��k�a��!��"���'��'xl4f*|ET�d���c��U���X`�?�D���o�lԂ��c��ՈVƘw"˖���E�=g4�28-Z��W<��XCs��i�?o��������;�JdK���).�/���e@�n輆OB���ǆ�ea���5������I˧ݎ�FO��x��0ɟGCX�6~�VQ~�׉��:d_-G����Π(�Z!�6Ŀ�ݼ��e6�gN�d���i/ �΃��ue��v�y�$�/�1y����4�3ЮG'�!�?�=:��6��`��ʺO��h�����k)m���I��v��]�;��5�ՈN}Nl#XBK��:�l�6K��n܅�M�C�+�N*�tS `���<#�9�Û ���\u�L�ֆ�<���y�vti�;?�-��;/V��;6��OBz�������H�5�\�&�'ku�M�q-���St��E���^���L��4q��]�Gcqw.�E�R�pwYk�mY���=���	��g�~#8|�#q���a.��3�]4s6�����u�`�٠��s@��M���=~h��C�����[�1yVM�j�M��I�p~F�D�կ��o��&�n{��j6�Α�V��,HH]�D��iz�=.�����c�G�K�!/-?��w]=����*����Ѭ���dЈ!j����É��~�F�*bA��@/Uh���rf ��Xr�s¾�"����\3�>���nҼ~D�`���lR�C�"3���2����L�7�]���H� ��R���R�J�h�G��Z�\��i�5��a$t@��m�ѡ+E3q�����a^q�}���&>WAׄ��������$����D���}9��\��Ϻ?C@�[�a��o��3����e�/^�=������S�Ӹ�o����e�Q���)���u{�Jo�K:��hb���Ү�z�L.��<���r�����o�;}��ׇ뗟^������R^ʍ�Ed �?���/�~����m��N���#�.I�o�:��8w�#B�Ʀ��bl�#��0�,�P�#PL�l�T��M%����Gy�^�*�ǽrWUp��`�W(1�� �Z��{"�p�(�
{�%a�pYEZW��}���;��7���_+�9xAaki���S�ޏ;��ix����]��"�4}-ڹl0Z����}%{�E�c:csǝ��S��	�j@g<r�e��C�| ��'�M�Os�ϯ������L�	��^l�i�a�����5�k�t�"�U�ZԿD]5⛏ɟ�����������|�GM��&�m����ϕ�y3{���&#t����'~����v/���,G�O3^�4%���9��Z���"�c�"����L˵#��we�qtm���5�ݍ��Yߚ�o�u��h/����~��ˎT��I�<p|D�w�'�y>.6G0(+��h6�ؠ��b�y�W�6�׸�ڍw��i��O����v�W8�gР��7#�º�8m�$����m��U�t�ֽ�a/��v��0���6��`'��ܾ�]����]T7�4uZ�T\GPL����C�p�ߣ��M��a;��k��t��\V^�Q�Efog��'�7ޘ�>8��i���Ȓou���\2��0b��EZ����V�=6�.^���^�3;�Ӷ Ś@όw��Ra<��ڳW��3絴
��Z�ԗgLK����K�:?�آ����q���g��rs�+�+e�ta��Y��hJ�H䇒��Sp2���<�
��B:��2����ǘ���`���ī��g<���a;�sj�6��.�G���ɰ����l��a��ME�e�(�@Z�Ї�����m+�4?�.�[8���]�N�u��ܮۤ�I�*����J���|��n�t�E�v�u�~�r�c�v}���6��G�N$��Ͻ�]�2��������a����ӻ��'��!L#����?��oao-q0�r:�73�g�C�6�϶��������=��3���R��B����Bv��?y����.�?��H7-��%�b���>6�z�s�r��{��q=�ȼ��m��m��m��Ԥ�=�u�}�u%��i�>�̟�7?��P��^�-װ����ґ!m(�q���-|!L7<��]��URb��W+��uo�d��g��!p2�"z7�������u$��N��s{|�&㝪/��| �4��<�F:e�q��q�K�;�D�D�.Z�6P������V����'ҋ�}i'��u5�c�d˺<�tӡ�ZGup�ut󕴤��q�h8�`ؼ����ҍ���%�`��&�%�N��>4�,յ�}�1ۚ���ݰUb����ϣg�ߴ�4phx0���5��D�(��6���1o�o�'����C�V�W]��g���m�M��1״�z�ӭ	�_~/����3�a��O�5���G��Mr���y�{�a�@��W���{ֶ�>-	�]c����y&�����9ɽS�;f��^)l�� �Jo�����DP""\�I7�, �a��XƤn~a1<7�f���M���Y/X���E}����%��ha2��c�\����~ԫ��x�m������/���.o�"�B�Ky)/�x�A .�����O��?���>��gʮZ�{dM��B
u��?`���,����9K�P���VFkw�@�f%�G��Q��uKD�����¹�m�M:����m(�kޡ��.�7��Y�����o�k��~���<	d�2N�\�9΅�L��a �B�V�,�6�U��������CX��v(泩r��D���Y��؇���',:q��HǦ8����Jp�z<�n���N>�0�@5Ԏb�h�d;p�l�I���[��Yk^�2�(�M�Z<M_#E=M����E[��5�h*�m��B?���"pY�Mp[����DX
��(��ʖ�
��S308���Rw�2p�}Ŏ�K��F'>��8i���O�����0"���F��IK��
O��c������q#�0�|����ԷO�$��Gt�w���Cz>><7;��(hu�JvC8���i���ll`�t�r�lKqB�9�m���p��ԍ��/$'�!�&c9�W7p4��p����G�Բ1�^3�#����qg�F��g�s��ׄɘ�;AG�*��K�+�s���p2�B���-�Z'��{�@��X�w��F
�3�tӉ����ojk�a^�ָ�A�֢O�h�H�����9x�p�x��]��uE��Y�����������d�Im=�+	 �A�)�}!�Kr�F�nd�����4y��
J7ǀx��Xǜ��~Dp`!�1Ѧ�ؼ�^�J��Ӕ�%�E�,C� ���u`�H�%^r4&���m
���z�N��9�q����F��[�[z�`��;�h)�:`�+���AirY�r�eO�0n�4�`j�rY`�7���O�4I�\������uL�M�֡���&qr����Vh��;��Z����g�ji|�׀��xX\Xd~"[^?D�N����������ɛ�o�'׍!'�;�5�%oӘ"h��u$q��R��F˰ۆldm������/�-��j.�{�>Ւ�OA��LŘ�]<��ۆ���8�`�O�Q�*6��Ë�3\��tL���㷫��_�968d{��N߻����ny�w9{�ͧ"�fyt<yk�
~���o����it�Pt���W�τ�m�=�;L�3)�l�z��"믡��x��Pt9j�dXD{�jy�Ȯ5����Y��w\9f�8l���$������z�J@�r��xp�A��q`*��ʯ�d8� �CI޺\�,B=���<G>1�;�7~}g� `��{��X�q$��6fw�p��gЭ������o��z��P��d\�i�^��L�x^�	 ������p6y�xc��%���x��%�Q�2�m*�@�.
��~��t�L��!|~p�u��X�]������h~�k�F�
A(_-� ]�c�iK�i@xjг�N���_��&�?�O���������G����A2?����\�m׳�hn�Qa�C�Pq�lk+��5Fs�zG����6��Q���&8,w)�d$^נ'��qJ�3I��ve���u;M[EV-��qܖL{6ϼk>���~d�C��4�а*c��We��n��Խ��J΄���C!�I����+�ț�a���naf�ŕ#�g��hTck����I�D��>
m�z��b�ͯ�� �$�׸:���!����V��2��Oib���Ѕ������ӵ�?����?�����<~���|��z�\�FQ����R~���`sy�ɟ�3?��_��_�ƫ�ן�>�C1|28�	�6�ń5Rzf}-N7(9��͜p����i�'��&�ap@�4K]�[��ӅN1�b�h��O���D7�Ȱc=�!x�R
5�΅RD	�Uy#'3΢�^ܷ'T���L�
�N�� �
@0檡�#&i�t��g��g�yLdT��oS4>�5?��Hm~�wN�GuSF�����������
��S��,9�1��Ξp�B�5���VN<�(�$ڵ��>R�u��tx�Q��.�e�ת$�)|}��)E5�E�aӶ�Q�1N9bw�x|6�6�bc�[W��Q�=䵀w��WcT�Xuؒ9��0���"2��aА�0d�N0�홳��S�����𷁷R���f�#0O7���hk�	Jt#�?��2gP� /�~�\{S�C&1�������d� �Ṿ�����5E�e�!*x���atԫ`pw#іn�5����x/�8~*W�F�I0:��\�x�5��w�ۅ��x}��&l`1����]Y��gΨ���5��q���p�\��P��,�w�a�lm�4�֪|�ċ�����<C�ǭ��|<ͯ��bx��5rH�@J�1����L<�9=��%�똦|n1����<>?xʐ��p����H�
L�6���2�&�\̼ᱱ�z�o�ʉ�np-�	wV��9��EP��\� qEH8 D�z|���u�5���?��������d�g�mMR�������:�����;��~���ء_y��zʺb�x��p��s��CE�W�dX[�T��G_?a?t�+
Ɲ���-�	�"���i��:�&��A���H�7�	Me;��&lM�*�[�}J�_>eA����e?�<����/3j�s �Q3���p�bX�gC�"ÚO	������h[�)����<;�!+�r�9qO���0O�G�["��ִ)펳� ��z-Pك~h�6B|�R$ �t*i:y#��?�U�� �Xؗ�`�SF�xN0���?��F��Ԑ%�������x>f"���1.A)˚GǶD{.ޓNO�t��+=w��h�u�8`E\�Ap��颩}ߡ��m�<��wy
Ph�Y��ZKj�5��Qډ�_�}� ��w?����?���zI��5IϘo�]�ƣ��[I�4OU�kZģu��3��fx����T϶S�(�J�������It��LN�c��)�ؐ��9C'6�6d�@�v����`"A;�oM���<�0�q��
��|8��:��`��<�t��$^	��K�X2�]�؄l4�n ��������*���/iAl��E�����zu� ����X��E>'��S���FO�sx�5���'�bM�xm�ds_��cz�YΞ�ފ�.1���u|6���=+�z�M2�l��G\�� �� 8�K�0P��h�r|�I�:��l���������.�i��rezf�1hp��Eʜ��W���
�o�彛Ӑ�t���/��迃�(DĀyu:���eq�����ʿ:�;��� �[yV��Y�����p���*9+K���DW���x�ft4p��sW��?ٕN�?���w�^].#+^� ��v͸f�/h2L����;m�6�Ge�_�����B+^5�}�ݷy��W>�����w?������Uk?~��3y	 x)/��)?� �'F֏��?����7~��~�����/�A��I�?��΢QHj�n+�����lU��:R�[;a��!`�\IH4Up!��qFǥ�#���R�@��;�R(�-�d$�>Ŏ#(L�ptg��AQ&�w���nʯ6�^U:��P�v�<�q�c��#XH{0��I���M�Y#�MǤ��@��� R���\j�-���>`L�6	kYmD�Π�z���l��3}2��oM�� ]���B^A0L�!�!'���ͲPu�|n�hE��6��y�P��JK��� �̓�F2~g4X��(��nS5�_8O��f�3*�BC�:�yN��r�+��V~���c�5,�*$~��iZτA��)��#u�l�M��ZW4�[��l�G�^����B�7rV��s�Z���2Q�s>y���/rZ���z�������w��[�I�W�Vs>9�LW.oK�yS|��Up��-�f;ø�l����b��G�(��5�M���|�\�uфdZ����cq�#��S��ܿ/�:�m��%�N�d������o[�:n=�Kl�_l�=cD�k:�.<ߋ��U���%ρv��u|��1R@_��k�jc���/��-NlB������Ms��w
�h������J�p:;g�	]3��s��˵�AS�\���V�.̃�9o�eZ�+>��.��t�47F��eC�?���׼K~�a�9Y�+'m��g����n��}����B&1�ݹ'���&��>��!HA�U��z�o~�ٚ��Y���C�Ջ�\hc#���tʟ��FL��t�stb82�ݥ9�D�<6ݒfZ�u�,��bQ�R��a�d���=��7�ɿ%Y���廰����.���2��z�J�}3�l7dP������G�I>�mf�i0l���Ѿɀ�'4�6�R?ŎB{�i��ls��E4�1"�:��d�����w���t�6�w�~��3/��U�Rc���h.��o��ֳ<�z�����6�	-���,�}d.��}�_a>y���,i�6�߄67Y�d�<|^�.��)w�:[\w��?e�q��y��n薛�e��P�M��ϳ~�Wlf=F�lm�Vg;P�a�8��$���/�G���F>�#A{[Y;���8t�Ef���������:$�m�5�d̬����t�	T���N~�?d�s�gT�c�X�[�#�)��І���L�Y}��u�^ �Lr�y�)�Ο��)�ɍg���t��ϋ7Ӌ��3�t�{M��&��P}d�A`b�%��ལ`N�oϽ��1Ǹ:�w�g�F��dZ�%�E�D�l^^G��i}v�^����U>�������K�؏|��__.�{_>�T^ ^�Ky)w����}���M�|���7��7~�����>����qTk�7�] �;f"�O��߶��Q�� �W"����}����8]�;<���ڠ��܄`E����?W7H<�I!��4&�)�[Y(D.�υ7D�K[���Z�.��ςo"�A�ݞ6����:. �ǻf| ŏ�P����gŶ*��]7!�}"�!��3#J�YQ�ަ�Oo��1��5<�9?;
6Yn���vf�q�w��F*]�1�>�j�Q6���W7�b������1�m(�Qw#�Y������d<�>��7�A��$��.����BsD����̋�a��3�^7��,O��̳yT�?N�6�<��%�Zᾮ��Xc\���rK��6>�<�+��V-���N������s�țl�7��Z~B�-�Mn��[��N�\�?�a}w�lFT�/\/�����Yn8l�W�@���4��U��S!ѯ�˶=��ݙ����|��˟:�o�|<�x�	�qp�Y�ר�b��c͕�Hgx[��i�7� �b���ݳ��"<�<%���f��o�T�FW_�N��x/�S6��k������K=��G�_��D�46��>D�~�S��mZ�U~�XZK�"˸s~��-U�YŨ>�Y4���U� /����j|Ff:]=��rK�8{��o��Vh�`l�/�rx:��l��>�6�]���ٸWk=l�N��/���g%�7�,Sl���xb��3gs���X�ī��-��C�����'ŉ[�i��N�r~y���Sf���Ϻ ɤIw%�����H��S>���R�I�e��' m\���aۓ-�s;et��t����C��o�:X�?�����R��Ŝ��w����N� �.���X� UW�����U{��t^��}�|��{�|O��U�+]��fD�GY���'E���jÞ��%�\�O�׵-�>��]<�^}p���P��y<���z79�(,lS�����z>ٌ�a��_ސ�q��W�4󐳹�������#�k<��,2��9�w��0Tt��վG��������mlk;��Y�W���w��Ozr���O��ߙ�^�犏V��0���+~�e��r��*7���k[���\m�3[��_a�l�A(�c'g�x�W4�~=��Yv�:�0ޤ�2�x��)��ԾW}`��V���q˺� 㚎�U�����v�k7��+9�BeШC~�Y(Dh��σ9��3�b�?��ǲPw���#v}H�S�!ߙ.��@�7�^Tx�g+=Ƽ�E�k?�S�����W����_.�Od�Y%�'�_�Ky)?,� �O����_���������o?z����G��9�pG�,`  �P��{�ٻ9[�\�Y� m�s7u���G�����;�?�FT�U�ROe�fW!a��T>��I(>^�T��F�.,��
���I X�x���̿ղr���չuY�s:g�<��l���\0���@w]�~w8�p��Q8p\6bV�f��T1)�
�w�i�:��;��!E�.v$����4�ڃB\��N���`S<ƪS��	�������[:[�.�.�R��h����l��F��9��b�*<|�������huRL���n1��NO8�;���'���ֶԾ��G/}>�a+�j�㷭M'MVm,�-�QE��(��e)8O���U�pn�2�n9��Q��#�<���ζ&�v���8�V�W��~�w��[����Q�X�_3$���v㳐�-��D��|�����m��{��`�̯���*M�fy����|���V� gz�8s<��o7�>�؉Dd��࠱��Wm*���0�,厜i�n{ʸs����&�g���<r���N���������eiQz\�Ȭ}�x���W�6�"�-6*�^��u�m'�ig4V�g�f}���7�Ӛ��u����M}��;64��W|��,���y�[�+�Ot,|�|�v���F�7�u��ں��:�i+Z*cw�k�N߉�H����U4��^�]�!�<��-D��!��_�k��\���#�Ct�H���X�����[����:~vf��&شt���������gM�[���y���c��0x�Fk/㩎��e<�>V|����y����g&�sV��Ao�YЗg;m5���s{�5����-��6C�1�YGZ��⁬����5.t>�Am�,�� �"y^W��
�3\��c���K��^�x����eNk.�y���ǟ'�Y��p�/�U�6qxX�Ve��Y�{0�þ�j����Gة�ԠA���i}���~iy�wCw�����ףW�����Jcx��o�'$+Z^[��В��M��W�:�����Y
MA�D?UGZ�����l-�+j��,�;��<<���I��Y�z;�}T�,�g�n�~�/�]To�uC?S\�'me���%_�苿���[>���nݶ�gs�����O墸�y�cv����4>c�N2��L{Uy������=Ca���e��ٍi��?Z��#���q�C�����vy}y��g��ׯ~���7���X^ ^�Ky)�(_H ��|k{{����w�������ۏ��2�+����l�b�̹эA���|8���	o����G$)2�`sw�%���é.e�Wm�S=�p��`�]`H��h�"�����u��C��\�[�@�B��M��ۧg�>6��$����D9���m�Z�n�cV�o)�����3��۷���á$��z#�3���oP�*|��?�Ml�>;��Cٍ���,�׹C4`�O}]1���b�
�&ܸRIJz6 �%��8�y�g�J��ʹ�s"���q[�ٳ�͛�<�l=1`���iи�=1^�c����x^_J�����x�v?�;kkeگ���6��U�<�ոW0lE��Y�r���o�NgՑ����[�hn�l���;Ñ�V��NI0?��,�/�o��lݬ���t�Y��f�p�Z�g�N�留[���.#���Aǰ�x˭�k���3Y��g���`�C���sX�7r�K������U�����Yr���[ރ��<Wcd.u��T���������]�[���)�x����������������^=�zj����j����o�!z�����[��aHk�~������z<����m�
������l��tF�Y���j-Lo�v�� w��[z�-Y|�ׯ�6�t�)�I*�F�W=���~����Z�W���=ؼs�Jm�L.ݚC�Y_^6��^ɺ{mq�3�ݳ��~\b-��u��Y��l#n�d���{kj��u���ܑ��ʟ���a�z<�u{ug�ƣ��Q��v��JW�*4��J��}�ܝa���=���r�5�3c��s��U���>{�9��ۼ�9���Z_=���ݫϼ�u�ÇG��ټq����{���l5w�~�c�\����ѻڮ�����$��t8~�-����y��O�:��pW�X��s�_ү|�2�&�� ��Uѿڥ�PN7f|�����ѝ�?��L�	���4����C��0֍�IWm�����W��G��v�ҵ�/���=��^�Ky)?��	 ����>����_����}�����ֶ�p����7Ӝ!DTo�y=_���8.���e�֣�C.m&,.msap�v���1E��U���]�Er�qc<N��`�#������¯�>���!�E���V>����˳���G
��8�<�ɟ��l̺���	�-��?ڽm������!�W�B����C1ņw�-@�1vkg�J<���}V����C���! �Uaк��\m?�/�Yi9�u�H�w�ݚ��l\<��u�i���v&�3"�����:��ߙM�I�{��Lg3b� 6�Ufz����>��}��Y{���ˍ�[k5����F���j�����]�3.b�b>���t���QV�銿[�▱��_�����8kC�G?�����L[�D�:<s`��H?��{5k-g�������������5@�a~�'���g���6*��qt��KW\7EV}ŜUz�x�9v.YO�c�O37�p�1�X����w�~3<�h��m���OV��uM�{,��39�h�׹�x4����zFsg�|V�\qvV�,�~��)<�VY�[���:�ϴY�vǊ��U��|�|�ӪϹoȞ�Yέ���������3��+�������~�ܛ�3Z����7�QO���e+�F����i5�����8 �����Z��ڽE�˭��x��J.�1�w�t�{��=ߣ�[�8���u�[��g�3~VA+g��Ҫ�Ug:%~_eŹGG��z��,#�����&Zm�o9�e����uم�V��L���W��<�'��离ԌQ���D�_��t_�v&o�.��k?�st�aA����?�4�w?s�j����M�����uV�1/�-��ۿ�;���w�Ř���C����@�3��Xo���Z�G���a��?�a�#�d�|n槬�r�g���2����(R[�z�U��mG��/}�y�Z'�{�_���W�y���d/6�C�������e�oۆ�[�ͺ�z�0��~`��o^W�a�o/0����:d��s�Y�;�,o�M.�*���������~�?����|����߼y��-�a /奼��� �2w�^�����՟�_�����^}��~�/��ޮzB[Oϛ�	�xiUسQ�)nTD4c�W{g��B@9�>��؄��nً�#�%�^��h�	��{��i��m�ER�Z ��q����!8����=N,��Fᠢ��3'�w[����*ah�b2+�wS\'��8K�c��q���3�$���鳸� � �ĉ�[
iUv��"	�+%���1m���؟�`_;�&<[��;���Z%z��8�`n�ܪ���W0δ0��m��=s֭�������f���\�l�p_�?o���m܃�������r��0���m�<��{���>^���-��J#����s��>j�w1���N:����
�g���2��N��9p��\a9�"�j�V=�>{����܇�o5�}?Ǚ��o��i/p���L��@�2���1�T�����G9s�Xk���ֻk�x|��C�Z����y�h������\u����%����u�V��������
���ݺFg��,z7xPn��e	}?��8�o���ſų3��]��sq��;s~ރ#?o�?��}-[3��RY�G���v�|�����1<�f+�p�>WN�z~vu�-�f'�����]�o˽�s�C�F]ˇ���Wv�λȃ3��g�˝��-}���8ϞW�^�uߙ6K?������~=����<��s8�˔:���*�!��V`���X�_����?�h&��"c`�a5��x�9�^�9��Z��y��74����W�C���OK���u�~�M�e��l��<w~�V4��̋�~ n���k�~��n���ߵ�Xo�MR��	+��˲`�kk�۳w���Z���������J�}�_ۄ�s��N�o���#o�� ˇ�a��?m����V�?������0�\�|�~_*-��h��q2�=4���;1�/���wۭ�,�^V��f�6��u���f�f �g�i}Πa�h��MMs�����\Oo����o�������/�����Ƈ�ȗ����ї�R^�K�/&�����������������������}��[kΐ���zu	g݉�ő��d����M΁��E����Dj&��8o���`_�����Ƽ*&̶^�N����DlA0ȉ�Zp~ ��3��i�x~^��ZYkE�	0��Q5��V���9Dz(����:��3�[�>c�([)RZ��D���u�z�4������m߸/VdQ�`����Y)r���)�R�W��:+���2�O~O�A��e�;г��4w�$�^�+P	�����^��?7�g'I���E}�~o�_�{f�<��z������y�eĠ��qY�:�V̧V���1���J�̓���sd�;.H�X G�Al��w��[���3���8g�����B{g�E�BK���Xk��d����Cn�ָ��X�ql��u�����/�Yz�ؗi,�Y'����F5��݁����h���3��>���������V�(�ŷo��n����=�o��3yso�m%���U�WW ���~a`�����yݜ����㻾ǎ,������ܣ������*�3�ø|��+[@��e�{s������v�j�h���.�����v����+�N:�e���/g���6���c��m����nw~��8ʽ���>�'�kg6�-<�γz�]uO�߲k+�Vu������~{�V��>o��}>g��������������I�w�Q�M����=��%2vi���ӕ���� ��m��g6�A*��3�8�ت�{��>���sF��s�z��s�������j����:1��;%˨��n��Y?����9[_g����]�M�9�8��z=�m��{�/��>W����u7�Y�t[�ܚ���_�d;p�i�cަ����-~�p<O��U���Y=�ww��>���T�Y�/�e#��8�Sۡw�6�>�#��Oq�<�n{3����D�ƽQ��ʷ���pEo\��Q@��o����md3�>a>���/ �R�i��{���͌èG��E�ǧ����}�(��'o>���د�Ư�����_�����|��g�R^�Ky)7�: `H����o<<\�����KW�><�]>�<�+�C~0֦��mۋ��l��=�v0vV�:ؼ�����7����F�q;�f 1F4%�6���\�%���Dc�QBJ����y���Ӿl���T�b��������(+#3��ylz%OVV*,9
����]�m���<����T����X!!��ʑQ��#�Y52��9I��2��M�v��jc�X�/�x��T���h���wvΝ���a��n�;%�&��q�P];��zʊ.+�3�Y�d�oYr pJ�]���Sa�]�����c�o��l�O��}�4>3,ό��ɷ7�(�G���}�	v:�}e���Y?�u�p{�a{N�穹�d-yc�e����S`嬩p�a��<�x��q���mY��Jo<�Sa[��L���]6#��q\���������8���|"������ܣ�:��`۞��̺OE�J	>�Ά�N��K����}�x��_�t����|���AZv��;�p�m�9~�&н��x�"	�!���Bwr��C;t���4
M�8>k��d݇��<�O�d����,��Wu��l��Q��x�\f�����|}�&���������k�V��f�o+>����t+X�,�v�:�{�SV�����z
��[8a8x�a�-\��W�'�n���0?�<��s�!�W��֊��=ث,+���t�ѳW�h�\�\�4q�.Z;[��ʳ����������q�XS����A\or�2󳐁1��߅���V�}�,\�`�Y��:e�}��g�2}�k��O达6W����vz��U߿�ԫ6��{w�Sϴfƿ�YΐZ��[��Zf[m��ʌոw��xܷ`�k]��|i�=x>������D�qou3~��9��3���k(�S�!��f�2m��WK0�z��{�Z�5`�s�ϑ]!��ch͕�bw���%�_(om39l{.�v���� �a-v�_���פ�M����q����o��9�ցk���boa���~}+o�7r��n��G����{}��\.�W�.��/奼���Ed �����������p�پ?I���M�DOmS����:�a#}|(��[�g�N�7�h?������v��dX讻��CY'�F����6����<�����|B��ƴ�3s	X����\��-K����f5p��ZghUp����f�4ҡ�ˤ�=މva�n��4�.��ڌo�}��Ws�[�)(ϡ�����Y��2�Π�Ju�Ǎv��b���`�j��+;A�G�Uz�)������=<=i2���}�h?��?e�1mO�5R �lȚ�HRd$��>����i��iU�;�X�=�FPu��zh
@��&D�M�-�N�P9��rPh\W�<��{��t4+~o�4q�J~|�݀f�N�������fW��;�����=��F?�]��)�j���l�����'���xX�5s8�zv���*�b��}�N<�yS����9ӊ��������q����4��������:Q����=�c��h<�dD��sY�������z�vRmZ{O��d���spU��k8�'D���"ո�H���<�5��N3���pr���|^]�bl��7�� ��CdP�V��a�)����L��;��\��+9^VtPǺ҉��fX+�з�/q�x^�L����s����:tbQ}5�c� 8�.O�]M�4�v��c~N�[K�[���x��ruo�9�N��D ����Zw��*�i|��� t�0��~5��b�~�����v�`����:'�5��O��7�_-t�����2ڠw6)��zi�Z�k:�sgM���<g|��yVq>˜���o�,N�.��ع{������y����b�V��l�zX�IN-��|��TCOB!C��gқ������������-��\Z���-�w�ϛ
�o�<H�nc
��ҿ��a��v��Q�׫g��z����z�����E��=�¦ȶ�\����{|*v[0ۊ�b-��e�+��Mڍ�`��{��|mK�'Wp�����][�r�O���|��LS5��ۛ�U}Xe(xbZ���l3ܚ+�7�5�0�Ưվ�v�:gĊ��8�6�~�<ƃ�%�l���?Ö����Wz�һG�@�ۧz�����c�1�খY�e�	~7��op����s���E�ɕ�r�����]:�M���s?g�ۄ}�Y�? a�Q*ߛq��+_�B�#�q�a��,�'�C:%|\��D�a�Պ���S�!�i���op�n��O���*���8���7Ým�L���~f���W_3��u��W��&���Bmf����ǋ�"�9���L�1��b���k����S��ܚW�Sg�-?�0h�D&;�������'��><-�c�b�|=V[�T�=F�:�����m�gv��sL�Q�:2I?����=���h��x�g	�-���u��!=B�V(��ް��Wl��E����<|�ћW?�3?�����})/奼�Q~� C������g��������o}�����G�>������2���]6�dk�D�v>��fʎ:A��Ŕڽ�;~Bc�)����,.Dv.�ŉ^ipTc�/���;MVJ����.!�'�hU{2�W�XU��ۄ��R�̛:�'��|��^1�V��:�=��S����c͉���N�j��3e�m���c��״�� �A�wz�������8q�=l�TDwh�{�,�}�&YL�C��UijS���>�πW\9�46�ɓ�*-�%�k���Of���^��q�Z���7����Y�am��uV��s�o�	�r��
n�������㷼9;��!L����Fqϋ7zϨ��k?h�:wWg��f�� ��lW�q}J��}-�m���u��I�)jc�Z��}~/6����[��x��r
m6o#��3Z����ͼ2;�B�Á��c���f�����m�N'x���66f�\��'cp�� �d��v���u!��8^�s�߱�� ��=��JO�Z��1��\�����[kdu�u����С�j*8Y^!"��G�]���S:L���pV���C7�r���,v2>���`�IWd�m�o]����I��gz�/.�����is��x�N%�&��fy=�\���k�۟*-e��{�x\�8t��z7`��ݯ�ܲ�ϻ����m�A��x�.k�-x7��}ks:
�h��*H�f^�fCR7����#��y^�Y�oӳ�Ol���9��<f�������̷�G�}�r�W%���o�sԱ��d�U�~^�͵��j�:=�u�-}����:I�)��~bEOUsq�}��p{yv��jS����2�y���0�
&��g]B�Ԭ���	d�M��ήPKߦ�׶g�[����Ѿ����y���a�~�J<�'�x>����O�����y�D�>ā2��s�4���U �S�{���Y�U8Ļ�s��u�z�~��-��j7��6�{�^ϴ1��2��b]�9k�������5�N��Y�O���.�u�>d6��պ���Z�E_��m��ln�u�0�d�$_�3�ٖe�F�7�+|վ���7Ϯ<&��>	�d]�c��d�D[�Ee���s�͑ѹ���KG?&H��Mh�uqX����3�>���,/�wA�qm�as\�L��d������?�����_��K?����;�^�Ky)?��� p��O}���/��~�~����ӏ>�����z<�	�GA:̕Rq������
����胀k��S��P����;�݋�����_TL���k�H�sk¶֤��H��M� To�˅�n}��n���B����U��>p��a�c՟:
�颡��X9��aj4��ڠ9Sn��`<��I)`�OvT�|��3c8�:6�߈���C�7����Y���;�ռ6��N����bLʼ�����)�/95�!���#D�Fք�}��2�hoӾ�6�P�̉�4��Z���ÁS�SNA��3L+|q]���E��	d}��ǉ�Չ�Xx�����\X�ʸ�;���5OE�/�'�o��1"�9pj�u86�� ��W�B�4��y]3��11������+}a]�����&��s/�����	������G�Y�Nԙ��o�5�cW�ǈ���d����ų|�e�����������w+�X]u�����N��s�����J���-o��.�ٲ>Ex_��uk
�7xQ�EM+o��D���}�3������JVl��rn+����q���z	��9@<��])�g}l���|)�܁Wa�O���m��\���C{l0��{"��u��,dlī�O֍PI��Y�rd��\�4�:��v˭2;�k�kz9iM���:�k�s�a���UC�D=V�ʑ��W��|���@`�O��' � ���&x/���,�s&�<�*+����8r d#����ϘC��g�^�5c4쥣DF�o��^��6�Vzm��1�W���s��o��HO���f�����KE2�������oa�X�
s;�;�?�u���~����ҖϠK�-��u�����^�@����Bֱ��*(��i�B��3�W���_�y<7�r�|E�+��y֜U^�����/�����u��Xn�_�c���*gmܗ���d��h���V�)�a���q慑-�����'��+�m��*]�{d��r�y����R�PǡyV.��5󉙶r�2g{Z@<=�eI�gz��W���'4p�+�\�^�Z���6;�]��!�A�|5���S�I�E+�m'�@��ON�]����o�}�<��*�v҅�G�#�~�׻�%�Ed�DPz(0��zc���:��I릫�$U��w7 ^o� �~�85�o7�J�!n]��|�B�wu�Cgx�u5�^C�_�뇫���<��W~�?���z�}���}���7/奼���,?� �'f��/{{��ꓟ�g���7�������o�g����~�����d2(Y��ӓg�Jg\�O낙eSg��?�����'�������o�`|t�@V�7�����9g����J�J��B����p������ـl�������~�k72�ǝdd���l�UyY����Jh�}E���!c��2h7����p�Q�P�7�i�q���jD��F������7cfeP7.�:���1�h<��1� G��lD1=�
�tx���4�/�������O𷳥|n0���ևcݜ�T�Ż���9�>ϸ`���sn^�s�_#�Ρ��Ȑ&8g�����(Z
;=y�W�Wl�V�i�|�5N#��vpZ/�2�^�g�d����1�7�kv��6��3y���pP�D�-�׭8��)���ʡ��3��Y���M<.�S�Ӽ�ΏXc��6nɟ��k���-9�e��q�e������������xpu��6c�3�a�����S�4�M��`�iW��q�S�XU?�s��!�*�f�d��n4dI��9���2Md��%6(Hϧ�SWB�xOc����_O�yly͟������T�8�;�|<�u,A+�3oc����������N�����2���:�ϰf'��Q�⢮~���Ѐo��V�|߰y��B�=�a9�p������dNJ�eg~1����32�f%Ɵq��6셣>�.�\6��ֲ����}/�+��:U��%�W��w�g~c׍�h�� ����W]��KWA���c��@}�d)����P�xb��*�KV�,���Ri�+=�8Yu�xJ�d^��/�N^�k�꒡���&��̺5��Ȍ��fzūH[�AՃ������Q��s�CR�W�[�n��}�BW�T�s�d�b��ʤ/g]��:��e8�u����2���ê7�����_ˎit�ϲ.=�2�S�������^���V'�Y�IZ�����pgY��k����u�'>�p}������O�gY���+�<2��V��!8{�������	]-�_o���]�T��5��w�V��� n��|Y��l ��"[R�éM�%C�Xb��g��4�5��[�N�|�y�����j��	�x�;M4�/�_�s��>d9�릿��n�4��s9��^D�����ӿ���o}����o����*o�X{)/奼�(_D�������?�s����?����w��w~��U��j�Av�A8�izo�uDH�b{���1f����d[�^8�;�/��:���j5IgB_8O��NR� L2�ҧ[:<+l ̂�ʁ�\`!�J.�Ԫ������f9}��_)������!B�A�@���3��4
	E�5h���:�կ�v ���{��~����y쳃f�-�׉�3tdc�3��;{U��"����G/�/�x��۲kn+d�5����X̋^���9 Y�<7T�i��a�T���~yC)����o�N�w͊xw�*�l�W��'�C�\?�.u�g8��h9c�}1�y�u=�umrF!sE�!�����bLy�i��wI�}&j��i�3�-n�ef�r��X>�1�7��tc1nvϸ2���78�s��J�ggN����_�#Ay�>I�x:s��ZI!8�,�ΝLq�%�-�d��J{�����؃���|�e���%h1�'-X��䱜�����pK'���ɑihuZ�i3�`b^�-�틬y|\Yx�=��qYq�b�yWd˼4��AḮ:E�_�p��j[��`�}Q�vT=4���[�^�P�*�~u���F����	^
>�m��t�G�(`닾��Pu,N�}f:\9��ɘ��LNc�F&T1?�LS��u��[�>�F������<��ۯ�Ldge%��Ι^s��x~w%C3/9�h<��'�W] �����P�y �,<�������Ŗ�a:g>Tq���3}$tۜ�-�*_m�������k>�Ͽqf��ӌ�����;m�g�μ���~�<v�mk|�qN�W��o���*+��§��s!y��I���t�l�q3n2�3mr[u����Y���s�!_C����������<߱��ڙ�U_֏bm���س�\�y�7��gV
��x8l8�;�M�?�pe�^�?�3�P��ם�R�x���{�+z�	������T�X�K|9��EN�e�00�3�g�w8̺pm�=��YG��3�۩~;�w�}3�u���2��j��EQ�ʼ��b��Ə\�����������������5g+���g_�	��@N�!Z
���m꛳Y��(���ix�+�ӺA�3��4���a�Yw��d�#xm1�tk�K��+��F�m��N7A��pm�����p?�e���>L��뫮��6��eu��s���k�o����c��\�� ���{��m��1�� b7Z�:i@�y���^����O��|�O]|�r�|$ �r�Ky)/�f�" �kO���������'���]����8���ul��8��{l�W-�,wR�#J~-P� <�PE,�Z(Ӄ}7�ו�آ?"�48�2:덍'u�oJ��w�hj���,U���E:�J"x�$��qv��Sa��Ɍ�x?@+c��(ClP��^������ 6x��P��Ϭ�g�I�ڕ��j�rɑ�l���M��Ӿhi��
+4���������9�8]�ꐍB6&�5;���i��w�T��B�w����3��#}RT��"B�)l�����]����(��ֹ�Fbm1]e��v�0Txnx~�(�J��O�H�wbs1�'Ƶ��P��e��3�1�d���F��B� �u��D���x���a;���6ف~�c��#m�4�	Wnt���S��yso}Bm��o�{5��جm��_���v�2����!���c,3~�g�n�?���w�ϲ����5a#0oRV�u%o1&vrU��OHgG0�uv�g�0����7��沞�^�:�[���yP�wu~]W���Y�?vL`�1����2�|���=�ͼ�ev�d���;�M��g�R?F̫���40Z�Lu��>�K8�V�UʳXK��|e�-Y��G�C�Rb������g1�w��+�羹�g/�~o!�ݡ�-ôZ��+�w�O�}ή���$�ȭ�ܖh�^��[��[�n#����{�aj=+�E��[ev�p%�6ќ�%�I��v�Ɨy<�˺��ϛ�a��zg���(��yh/�1�[��f�I2)�S�����L�t��?��7�y��n�e}c����gqƿ7UV3_c�:�	��m^�+��P�ǰ�5��24��ڜ�1���	9��zݬ�D ���S�\��3�	��>�Ù����R�!�>�MBOY�d��-�df����,d/�@�)~�qf>�u��M�^�|��W�fm��l(��������ǖ�Ě'd�3�}��x�~+��:[�D\��:���9|�kƳ�|M�b�G�����k��rm���'z��e1�r�7�Y�3��~W���h�����l�g3y�y�<���F?�.���.��d��0��q2̲#˖�f����,�g>wo��|U����8�}��}��1������B����#�.� ���0��P�W�Y�f^�|}���Zgnw�C7"�U�h:��ZK_��
�[�!y����#������Gϓ5_�=����	dS�f��Uo���	��u��U�������L%t|V;��q�\��������?y������������ |�[�j�뫿�w��W����>�l�^���e���9ӻ7��Z䡀�D�l�A���q���LLqݠI7"`�`ٽ_�g�I8�l�K\=����.��5�yP�~���w��l�@n�Q ���P�I"R��Af�2BL"1C(��H�EB ��  �l�8��ྸ��w�]����z�g������	������w�U�V���U7u4�tD:p�˹J��!^�idtHGۗ�+й�Ɯ\��D�}N�U�.�qG��u���oW\L7)�X~�
У#��N�ʎt��y�Ⱥ�K�#��(��r�Qa�|���|X�6^-�X� y��c�w��;d��	i�r�e|��s�H6�h��bj���6���m*�������𢑦XG,��ש�Kxx4�����eMa|��c��h�w�P���1;& ��Տ��A>�w��mk޸�����޿sǞ�~�d��V�eAm�Jv�ʻr��������m.A*�u��O/�	P�Vǜҩ��UW���0ҩ4�'֝~�����^�6��k�u��������!Z"��)��q�U�G�ƶDY��Q����w��J���`���E�_�Y�=�;�WGN�~�|��|�鷫1�r5��H5`m��5.�X�]T�������2�!�0ᾴK>���<I�߯'��q�w:Wg8)�~��#/�&����{�u��՘Ļ(�Fi���=ǥO8�LŖA�W2p=֮Rƥ�8��������
K��k��1s����������|E��l߬����^���J�d?T����o��`5�Z�>��v9�9���B�8i��Ĳ��&Z��/Y�����Y���Os�D�:�Ν���*�ʈW�%���7����m�-1q"r��>'?|Qol�*�p���8��Ό���k��2��2��6�4�?�Z�q�^�O���/�
��ݨ��=J�n�yP��[�9N+q���uq<d��D_�b�Oz�{����ʲ/�]�9`,�!�����s����5NͲ�N�׶����[�:�Mr�X!/p�4�~J����0�ᏺߨ;��������ǻ��YN)&�����ٴH��w���U�'�ʪO#-X$s��hU�r5�T�u}��m�Z��&yC>Җs�-��/�~r�&x�..Ӝ�G9" }�Ӹ�r,����J�����sP�Yb�'?��^�*w���$8�����!����>�$�ϓ�΍)�}�~�~���g�/>��_v�������:} ����_�����/����>�[nZ�Cq�n7;�ԃBx֍�^t��MP�
�ݶ	f&A�td�vq�W��'�U�y<ґn�WGǷ�>���#!��kj�j��s�red�N:+k�����5��g��,�a[�nr'O��A��Sͼ*��g0�e��>���ʈ���G��\��A�����Y��?
 Yv�@�o����N�(��w
t�nM�9�Šʵ<�*�%��9�9_�i֤6:y3�I���^��uQ�U��u�6x99�.�x;���e�5>�k�ן�V.~zԮ�q�@�;�|��w>^t\�#ў�;���%�������B�h�z�������s~��w)�k��o!���Z�+�4��l�7����7�a�G}�⋠��<��q�ej=LE�<}e�^���X����6����	�F|S���6N9y%�u���W$ŝy�k�|��F\����OE�I�c�:����X�N&j��c����p��~Vܑ��6��ne�]W��E���y(_X�����;��zqʿ
>G�ĸ�u!E�*��+;�y�N�+�3=`�OTt^��ox�iW�F|����>��:��7��a>ե�M�]O��v�<���&�p5���>���U*��z�m������:�j�E��S���Vޭ0ț�#ݷN��/�_�>k����?U���*ϣ�]���q��s��=	��_�<��9v6��n����&��܊+`[��Q?p,�3�F����jOS��δl�qD����=C�C�l��q�ܗ�+�9y�76�f�w�o�!��/�߭#d/c 4�W�1D����u۵�{�AtAqԻ���}�8�y�q�J��{~ih�	z��u���Gc ���-��c|�+?�*/�扈�k̃������[ұ:�GS]8����ٕNu�1��r�#�r��*�mL��f��r�!nG��/���Y������-���%ʋ�)C�z�k�U�_Oq�5�ԍ���7㨬);�Րo_�B�>��1�z,�*��;<Sڻm����B����r5���E���ي���H��?Ky;��yz|����g8Ffl�����iٖ�b{_`���;^����������v�G�ZA��rw�;�m����UX��8޷�ê�+��ا�S]xmS����xeD7��xЌ:j
��@J85�T��Sf_`3��d�)�s����g���g�ڑb�:������E���v��N����,��j�������o}�������/������ʻ����{�z9�%���t�~� Z���w��>���˿���>��l��j�W_�w���e�a�� �O�c�1��K���\����A�����:�]�� �ȏ���C�J� ���+�[�� ;���"�?�����,	ME`s�&��k����Y�&ߔR�ƛ 96�?��V�?�9��2;��}����0
o[�r�U�?�y���xT`�w):A�e����q�F@J�O g?�uB���vEIm����'L@����-�.�.�Hy4��|c^� � t�LǫB��ځ9>�KiJx��w�'��T6�r��e�\;�N�O�ǣW���)m�w�%�����7��Q7E9[��C�ΏR��w�L�-�W:�Ǉj[�Q����
uI7�v��ϣ~�����wZSg�6��ڨ���7��Z�-L��Q������ǹf>��e�[u���Zg�	�4���O�Չ�(Cl'',@X�9���o4_�i���>B�՝v<1�2p*|?�^M�Ŀ�oŇ��뻁�����4:���v���v2.ɶX��8�Gۆ1�d�~�#�[_s�;���=/T�
�>�1|wE�ixс�h��\a�8��-�B;�z��m��V�-�]�3�tڇJ1����X.逜)��J02v��!��&o�M���<r����R���o���vx���Պ�u�xy��0������m����w"�7Q_�ޱN�@��s����x;�;����%|�\�]m}�8�o��ٖ�ީ]�}�m��}�]�z���hT&ANׁ��XF�7Y�nH{��֫yцb|��p��s精��i������|�Gkqu�:�4ѷ��^�|�V�g��A�����8�1�WW��W�9�s}�r��3���t�i/�dߨ}S�_OC Jjߊ>��ەm��8+�X��5�Z�<�`iK w�]('���WRɕX��M݃��S(�Go�@�V������	?�ي/�wƷ����n;d���vd�)�9/��!�G�S��G���_���)�h�Hk��)n�G�kceOc���z��`��&ˉcp~�����q�B��}���+m2c~�4�\
u�2�7�5%�7t3�m6���r!���br��e��k�=�7�uuƩ�A:�T7�����g��1�l�q��	���p.�s�Ц�2�Q�S�l�wmo��n�����3|ö��M�@��3�T#�%���<)�u�ߕ��Qm�.ؙ�T|J�؁����ͤ�ҥK<�G���a;yhҵ�{L�Y]tye��s4����V_}��G?|����w�¿��?����_�������x*/�%���� }' l�}������w��T?��g��~�����q�_�7�	�K�`bߟ�AݱV��'ƇSQ�=}P�ƥ+e���_c��M�V�J�i� \�6���8� �nU�z�ㄇ��e����}��So\�j`���A P_A���'�t$�y#:t��nw�ܱ�N*���E��9�11��>�չž�v�}���8�� ǟ}�-�>J����i���ߏ	��NK,��C�8��ODw�i��qIK�!�5�qW%�xM�AǤew㵃o�D�
�O��m�i!���<6�JMt����n�Vo})�8
>ϟs,��oR�I ��bb�A"��c��.�E��8Q�c8�bD�v�z�}��w$��p��_�X:�e��Y�Y̶�֜
�#��m��^k�_l�+��G�2`I�0�Q��`r)ܥN}��x^&x��z��m�����S�it�W���5�!�6��N])m�q�@�1[}�w���!�C��ݜ�(9��~��܃���cgA/���-�9֩<����䡖���� =�����*��8�.�G�_�x`�Λ���1x�ļ�'��a�[��d��>NI"&)�mw���<�?'�t|Qx�Ġnԁq���g/�@�/��$�1����|�&m<m��6�'?����ߤ��s���u�!��l��-��x&�!'����'um�֎���q'y��1Ж���0*!�hƾC�r��sQO��ﱝ��!,��q�bog�"��r��
d�N�����;O<7�P�"I�Ӣ_R���JG�}G�i�-�9��^$�+���$=��g����~�׹m�0�x�6�c�[�۫���ex�`��_ŞA�$��h�;�KI`��:Ku��lo�������xЧ���{F;A��mǬ�D/�=���Nl��WѾ���Ue�Uk;�gS>�~�؎z��B��(�c{��x��Mv��ev�D�Uy��pt���|��������X��'s:\M>w̓'�Z���"��&dA����U��� =�����J���B�
��ӆ�hs�l��M�H}d�qE��X<�E��z~�u�g�s#>����?���D��)ڄ�:PZFI��Y�ǌ1��B�'/���0�d/�i��o�f�u{�Ͳ��d�������S�T'w��#�-N��C{�ٮ7�崅�{�L���h7�X���9H+<)�ty�<���x<R����yL��?e���[Y~���}�v\������M��>�@\er1>OAC{��
Wĕ�(����&�AN��>[\��'}�����k��(�0����S5��lg��DC�����7�?�01��J����:�nr"Gğ�_�����o�����"���ie+�+�8X�O���!=������o�C�݌��}\(G��q�S;"����D����]�n=�����1u��|�~����@7��q�R=v<����A�Wb�m>�5bf�X���3*Sc���w7,ؼ�(��������9��5�Kc��s9��p���ž������~��_�������G?�'���?*����/� ^�KzI��'� �Po���;�>}�����S�������n�z0 F�t,E^	�TA�fu����h�|:@������|q Hu� ����i8W�o�w��^ x�<!E5h!$G؝�U��*�3r��:������àΣ;p+0�Zާ��dn���`~��n�8� `i�D�dH_���@��S=��p. �4�Ϻՙ��hG��IG�"���r�Dqj�;W�M��)��
d��)�qi��^�HPD���wfk�|��i�G�CVK��4u�<�P��ͲC�
��ȋ/�wx�7:�O�du�x.GZ��;��Ϸ��YZ ����yg^Й�r���V ��'Y�bv<�c���U��rTE6\O�� c�{�A��V2�+�Q���c]��zl��������\�Ohju+��<>���{ߗ�ӑ�������8�;y��������w�Mڇ������1�]S�du��ۉ�z������q<�s�p�7�0�t�;���1�>qw_����u�ab�z]e��Xa���(Ѿ7���M��� T�GH�:�z.����3�֤�ſm���.�=�Pq��G0p>g��Ɇ�1L;WK�U~8Q�>�I�Y��l�ر��}�u0^_4�r���k���:=W���sơg9Ң*�(b�U�J/t�j!xXG���x���� �b/��L�T'ޕ}�)���=a���>�{��-N�g�﬍iݏ�1��ש
�l��"��8=�:������������ק��t��/�k���N3d)u���3Jif�yT�jA'����g����VƱ�M�C1�~E��ʦ�YO<��[��o��ޢ��+r��Q履ĝ�xݤ^�ܪs���z��^�#�Qn��o��>Q��@�ǿ�~{ǭ�� �?�=�x*&�;X�1��%֑߷m�8y+t��o��\��H�y��GyF?�6}K�f�:/�m��@�E~����\�Y�4eެdO����V��*���cQˊ���S��V�v��D��v�i�;��c�r۫?s;�;����x����m�~E�8�V�+��ek����o-vx5���2��>�v8M�3���l���S����y�}ڹ���Z�^_�������I#C'�,hi�(X�ֱiT|�o���>�����?[�(���գ�;�������:|$辽ms�U��� �.ɂѻ��z��w�����dvo�����c��Iuu�gM��<}�t�EV�wRB8]�z\��:]�^aؕ�k{].U�Fۑ���<F�����i�Ol���b��av���[��scQM����v�W;�#�d������q�	E��}�?o|C�0����en�|�������W���7�===}��w�KzI/�%=H_�	 �������7^���?~���S����C�����#�#KwL�N��*_w{������(�ۖ��tCq�D�b���~�=�U ��}�U��+VQ示�h/�X͑��a/�������������O��ȸr2܉���?��"{A����l��:cÀN���R���\*%p���7��c��s"���M�\%-˃�d{wJ�N_��e��*��G���N|���Ǿλ
���H�F ;d��ɪ�x����x�l�8>X�@�c#I�d��"��zч�F_	NR~�W)02M(�4�3u��@����'#�u���D��7k��c>,:X�6M}1x�`�D�����Qh�5��M�Y��k�,���,߱S[�P9� ���q�2�x)�tWʴG�@�>Q�u�璃\�A>TDP�.�U�g7in���ي�+�QG���X'kxU�Nt�^�НL{Q�jj]�]���7L"�"�>9����b�,�<�	g�Q�y�V�������v��U��?Q���Cv��1� �u��(��1(�}K�z<���i��/{��q�GL���z�2�������N��X��V{���y�m�|B �.�Q��W����vP�0�%-D7q��j<�1��@>���֒���� �q��C���r�ߴ2'�J�*���q���.���Fƶ�~��?Jט
��I�9�������~@�ؚuG��Sϣ����"�<����C�WwE�D�#������ʦ��f��7��I!�F�)-^օ��uG���Q�'��Lo?�E�+L�2¼�
Y&��*vt����z|�߽O�?1Eڴ���iN<����FJ\�C�Q�?T��3���@���?Ng$��%Ѷ�e2���)u
l�bXs	�M�\S�k�p��S}H�m�xe�}�<��>H�|հS��C�'��{�$6C_�/�7���h������X�X%.�s,��	|��
W��R�kF]�XD��
��s{J�L��,d}����v=����Dq�%�fǧ�9�,��o�à}%˷�;�}���y�;'��Nm���Z&���}�~���{��N��`��^1�6�o8϶�]����}�ۑ�dYǬ�_mu�ٗ��w~��]�fԃ=�IO��$�x�B����g�N�1�����~���h���g���1�'.���1��/�oJ+�e������{�/�U/���Țn�C�����\���_�/����uQ�X��˺�����ccr���͘e������}���t��S&�`2��Gx��/���~�}b�Qk��&2��:t�랧��o����#�/��?���{�aP�����^�e�I/ 8���#�p�G��'>��_��?���O��z��_��~�&g r7v��m �cW����N��lظ�X"
`�Ƴ �f�tC�ߢ(�&�p�eS�>�ne��l��
�����6�rz�{�қ�mu��NUM�sz苠�H�^�$x[.۬�4�;O
8��4����F8�8z7��`_������,J����m�uB� 拎�;oG�Qɨ;�ai�>� E��!�:�BJ4 Fh�%�C� �@�}q�GPu?�z�m�Xw,��׾�����]R?P"2G�c����Hw/��繾z)�'5|�A�\�m�O 8ƴ?W��+|G��۲N�I�Np�V�%�����g��d�=�K߅��z!k���{���/M��;��cY}	��.�#{}"F����π�_Fy7��o�xns��˛t2h"�G2����/��;v2]>����J�OeB���F����<))� ���+=��	#y���Z���	m_�z�j�����e�I�~�2�\�_��B݅�����#��m�z��u<p��p�@*ۜu`OX���VcuX�G6��^QY�Sw2V��p-�,~�ߙw��Q��`�E��z��G�����UvjB&؆5߮�������ꯌ.cIIƑ#.
%�*��.�0��|=���DF���6paQ�}�粵nuĉ���aд�;��a�1�V��&��+��@o�r)��)�P:Vr}�ɑ�/}r���`9����x��[s�o@��*��s�F�E?�|�	Q��q鋐���c�u�y[��w��vLn���qz�]���q���q���)�+�<�k寨?�E[���>qj=�e��y���{��ٯ�3ƣ���O��=N�Q�K�4zdj���+⿵>�	�l��W��D�O��I�)�R_�o�	-f��N��Z>u&�����ĺ&M�~���׵/�?��N���#k��ƕ�`=����A��{ρS	��Ai��{�`eC�h;�6��������e��CK>j���.�,���i/�>f�bE�>�TSBO���8�ar/���꘷�v�h��f��9߃�7�z>�1F���П�C�~;=������Pݹ�O�g�;ۀ�����D���(n�i���\̟{X�٘}�O��c�<��'�o�pmZ��O�v�AZ��(�vY����n۹�4�H�K?�<9�xV*?��W��������z�Z��~��d�KzI/�%I�2N �?x�O��/�ÿ�_��/�滿���������^���S���7��籷�e�#��\刾��Ծ2 �,���1]e~1�:=WXU��x<|A�:h($��9����� ��h1i�^��r��zS
Z >���t�%�.����@�~�FN�6����4u���o����I�d��X�݁�O�2���L�ޏk��#�i���,��ҩ%����e*N���]�y�w9���Q���l���2^9�+'���	dV�D�XN��/Ϡ��6�i2FY=W][����6�Ϻ���Ϋ _����Q�}<��x�|*�L��t,���v���XvG �(�I���[�D������X۸
)�ۊ�~_�D{P���rW��ez<N��T.wc:��Ni��t�g��M1x��5��έ�T�3�/,��z|\�b��o�o�7w��9ǽ:�s�Eٞ|�<�zb����x`�[�B�-~�˩)/��<��hK�q�	�pG���W�̾wYYMFv��Q�9���_���������Qe/���� �`�u�M�����
Ay�����K�xEu��rf}�z�cX�Ư�`PҏJmF�~eUu|�1�g=ү�����u�N
ŅE78�����"f�Os!^)3�b�
6��|n�(&X���`ڛ�<��Q�4��.�}�qv�[��H�ƻ6v\M_J񜖕��
��`��bC�&ϗy��S�J��د�˯=�;�Ap�Ͷ�2�ա�\��`n��ծ{��L���3�U�<n���G�>;�5�Y+E�M���/����]�R�c���d*��}��UY�j�5��x����->�yƅ��N��>�I�DN^ȵ��o�.���t��K0�^"�Զ���-_MF@�F9���c8�z'�@��Y~<!'b!�M����GrL���_n��ԝl�`�Z��e`,ʾ�v�z
�۵J˕�ۯ�����[.��zUq"�s��~ˋ�p�:m����"��"Ɵ%��gW��%����N���*^ը}J�m셾��rT޵n��I�:H��A���ޏ>fЖȿ��cR��Y�õ���.j�ָa�ZʗuM���(\a��<B��js�,����_��Ug_�$����(�5�D�M]��m�;��Zx�T���l�:��$�;��.�f�xjG�o��RB�����T<8��XD�z�}u�@�J��2�=�3^��>
W�t#�ӻ��G��;}dYq=겱��^���M-�����Z��|/��2�#�D�~��h�e��,G���]ʕL���k�@��бj����k�'���-�x3�k��lR�n�!/_}6��Ν�c��� ;�^�b��O�>�7�̿�ɱʰ�-������gO����V����釟��������|��;�|��GO����%�����,�D <+�v�W�_}��������?���������/������S�s��j�'#-
Рw���� i �`lt*�!��#T�nΫ�A:���y7���� ��م2�]$�Ǥ�m6���/mA�:g�%0�dLʭ��?z��
x���'0� @^� P�\הu �����C�'�� ��N�h��u\�̣�Q �}��K��� ]�rpR����6k���m������y��*К�4	�Z{�,�����Yc���	���K�5��"�Yo� ^�=�v]�������%�2Y��Gg��ȴ����	������[���t6���ߨ/�'�pt'Pt	���}m'd���
(#��5>���Q��A�<0����۫g��Ƙb`�������D9�D�ö#0��-}��:NJI2����^_c�fs�T���?��3ml���Μ�u���k�g�n(]S�=z̓�%�y�����q�CY�s"(=|~��$��3���3����ٙE���~�c��A�&�|��J�k�m�����i5�Vz��6��dC�KW�Qy��7�����֭��	2�~��e�����O���&��U��
:�~U�87��N�͜웻�FA6|��й7k��؎�@��dN��f�m��(32!?�]��׍�۪J�Q�������j1d��H��r>P���M�~p����H�)'IoJ�\�鬵f��xb�Ҵ|��cAD&��ݸք|���2z�tcwс���=M��)_J�� �l�?w ����q?�A���y��x�f�qa��hV>��-�[-}�~�~X�E����<�K�6�%���|��^R�e^RW������~��5�S��o��Z���QWE;��L\Hq��o`	L4��WL��U=�Xs��O݄�v��j7���m m���t�!��-�o8�&uR�bO�#�>������&�u�mS�"vU��=SL�+�;/V%OV�8�I���@|��1x�I�Y��1ʧ>Z�(�z���1�8¿^���Y��:�>����\\������z�j�畏�2��G�ig�l� }�s�ZA�W�m��vYiv_}"策�}(�����XQ�n��Q;���5c�h�V�O���S�4	+s�i��P��A�H����F��k��ﬞF��W+4�x�/�м�;�/9�W��]�Q��byXG�\F�K�o�/.x0��`~xh���cέ�����Q��o�C&��s^/b��s��O=4hi��j�9莲�����]�>R�&�s�c�么�8����������>~ƕ���������^�ӗq@{zN���s?��������G_����^�V<Rq���Mt���
T:}�lC�f�?�;=/Q��{�ȶ鬌��&���U�u��~� ��@�5悉�w	<+�۫�f+m���G�*�玐�3�o��\O����N1����XW,S4 �]^odWN�'Lt���Aг^��΍�+�$��O���N�+�h������໵C���e`͟��AM㸌�	:ώ����m��dj]�DPcW�f�|� �z|���	�4 �v�V��1���&�NArT);�s@��:F�_1e�Z�b��J�~up�v�Ye�r����ܲ�9��r�A�=�Ġ�W����8�nkE���k|ä�棼����0}����(�s7�u�r�U�o����ܞ�&���!� դG�g�;ϰ��x���R�u���pX7��V��h�6�B򠄎m��J���}�Nl,^��vo't��(3��z\>�l+�Gp9�
LW���`�T�I	*�����.@�G���B��_Y��q_�^yۚ_��}��� H�wĻ��ԋ�3��v<��\���*#��|ᐗ�*x��k���;��wʠ��ű��b�;ַ�/��`�[���vh_��X
1\5��8�8�8�����:��g��Y^=L���ʏ�E�U��*�J3۶��^���|�)_�[S�d?��~F�1�b��zJ�Y�3ړ����G�Wˏ�� G�E��-��T�t4������/�+�_G��>�D�*ˍW��>�7��aS�O1(��z�����+����>P��}V̢�3ND;��r��V8�J,p$�j֡폘z�o������4��RyUL@�_R����,c 镰��p�ǀ�U�/T��'LFmW/�H����I�u���_��ԿS]ʶ+���x�dV�e�i�'��,�ً|��'�em ��E*]cʨ�U�'y���]<�Z��&�Q��[�=����'.3_�r��K�W�a�I��Gˣ=�~�.����ن�q�i����~��>0|�����sk�z����>�����J-���R��ǛF�L�Ȳ�Y�j<�s���I�G�'L�z�m��^���:���:��ڿ?�(�hSG+��ҞV�7��G�},��m���ےq�]���Zȧ��alEYfY���$.rn�㲼1�n�cOq��h�<r�W,OL��ZV�G�߭7KY�w���60g�IZsvN!(&����2��<7{�wX,�r�m,��W���A
�)�
�����뎝��i���'f�P�qz�Q�W�������������j�ޫ}����{)ˡ��^�KzI3} ���ӽ>�O����O���|���7��T*�>�ަb����(��@�8����&�;'��V���Ciw�{�;����>��ԍè���y~�W��:����6�v$��r`��tr0�����8�+ �)��7��F��V�9�h8Ͼ\ֹv ��<��x�z1��!�%��)u��vжY{4��7Ѳ:�>	��[w��d�d���'6򖁇�W�C�� �W|�d�:)t�����c�x�����r���-\=�Н��NN�:Ϥ���<�vt�߮��`��:���N��U�De��5�1̿�L��(��>���F=2�eӁs��߻>�s�q���U�3�
����4�m�ímt0�U�*��z�6�W�4�sM{AP����A�c<K�<n�A���wt�ٷ�#8���U�u|��b��Y�\�R�4h�A��q�]�>�Pv���cu�������� p�|��r4�o)�W}ر�b�>&��3-[u\�'�c{t��wG;�&���1E��$��GZ��n�+[���B�V"Km��X�28�[�c��T]����}�|@8_o�ߐ��N�2ֶ�x��c�w�+���=�'����񤓘|g$�8�2�Sۧ8d��ľ��o� ��yYO��_��q�8J�l��2rԏ�X-'/��,s�uL��:9q�۵->Y���4�]�]���g��6�w�	�j���r�x�czE��k�ȳe�����b;R�u���fu�@-�G�ùώ;�]O�6��}}�3�O�S���G_T�,��2�[��qI�'���3fns��o��.���<ۥZ���=�1����v�Ǿ�cJOr�߱����e������<�����؍�V�r5���ՉZy\ѯ�������ϠW�srm�;�跫�uگxI߯�,�j|AF��]w�'�:F�����&u��	�_��g�N���F
�>2����
����)���2F���﷓a��j\78>���u;t\�������F퟈��;���f��_fn�g)䫎��'��'����qv,a�38��X���Ŵ=��joV�('���&�MhG�?P�Ȧ����온{U\O�q���O��{�1�����h"[�Z/�l�j�5�W#.�c0��ЩC�����\��m�yr�q�>�k�z;|�[���c���g��ȣ����L�����x�a�w#�y�OЍ~=A5~��ª-�G��Z/�1b�.��X�QV2�b'F��5�(�v�<��Q&�ķ��@d�5�����z`<��U�^Ƹ� 8du]���ˉl��E��e���?����W��gй��?��_��;{�����է�O0])��^�K:ӗ� ����������g�/���k~�������;�tL�ygN����W� ��Q�+
&a�Z�c
7�vԡt���q��=c7Ew�oϺ�v�Џ��F�W�N�:�N����t��Ѭ�:<���hA����G��N`��(e�^�����Px�oU�M�w-�����*H��D�ol�]n����:�� �ک��3�q��i�OgW�ͨu�����{������ּ���㳤�|�;N�zP�L^*�La�<җ+l=?'�u<���̏cM'Y �ԙ�Y��bm�@̊��1p5.���x�N��Z���'�V�g�`^���=~�{g�L��r��䨔R��^�����9 ����i����ܚ�X;�W��͜����{|��w��> -�n���3��o֥+�ݦGg��c�g�Xh�T5 ��@���]�e���P��ߩ�a҅0�uz=��zspa�S�a�w��0�_MB^u�z�͊��O]�#�e��q�n��w�ރ��,X�T���h�J;i;�;��N��:9�������2&cv��Ol�:��T�1�����ǃb����zo��r��h����Щ�ٮt��;��_jվ�z��v����O�+�K�B[Uɗ.Syb�|��#ZW�Y[�s��F6X���q�;\�~R�«��2��v3�JGa�������9�N2}�������U�=~3�>3c9-���IH1Գ˩5�GY��jx=Ay�CeyX�a�}1�-�u\��zꖚ����ߊ;;^������qe|�Skb���D�vx��hP>�)S�7LQϯdAi��_���HmO�}�У>�^��=�7'�	�O��L��=����{����׮ �r�qyr���I���+�<ZN��7�'.4}S�B�!�E}J(�_�S<��y	�}�%��<fb+[Ǜ�ux�]}�X���e֚�z�?�x�]���i+�&������㟎�k����SB��n�y:lö-mO�e]ƛl02�c�BV�^�{aW����4ᓸ�C��U��16��V�8VO��:���������cpj���m1�.��o۞�u���f�y�>�u罔�m�'�ǿ{�i�u,���}Ҫ�꫽ŕ
W��0����(��@Y��2�=�Gۡ}���[�B���ղ\��ܣ�g�g�&s�sDk����*�.�]��%���C�_��:�ƚA�!�8_�� `�c^�lo^�4�ć�ف�q��Ū����y0|������/>zz�����w�{�=�dxk���^�K��_��. hcF��������_�����o�����G�������م����0��W]��q����.�|�T�g%�0d��߇򝠸̟�<���w�yo简�|�1�쎏���N:GЦ�,����0G1����ʾ�mk�_�qjG��FIxjΠ;~� ��ש��H�^���I�?�V�������0��,3��r����uy�3�)��獻ߋ������U�g}(���ht�K�U���.}��=~C����z���h����������wї��2i:�����H�O���
'�V���_^������
��D9h��4|o���=� ��Uu��q��\����e��s��|?��'eo�u|�L���,�g�(�~M,�3��Gˢ��/��2�ul����e� 촬��6�2V�
�o�~v=Ǿ�����sP4�������D=�2z~}��:���#�9�Q��w�T�n�����O��vu��S�7�A�Nz��A׭ǻ'��t��� my��=ߊ.L��tL�<]w�f���A�x������7�B~)�`�)6#��_1@�`L4o%M޶2�X�z�|v�wLn���;)f�e���O�nc�CnX���3[�W�f]�ȟ�v��|��t�%^)��2dp���M�Pf�w�s���e������r�����пc����E�|�q���W��=S9��lE��H�Q��=� �^9�~s:��ˤ�A'<�ǀ�-�*��+��
�+�����9&i���V��*��;1���$�?���#\��l#�x�J���ڳ�'=O\V&�q�*|��z�S����Y��F�w��ɑi���`.����L��8��n#����jG����Kb���3��<� ��=�娲_ç� e��v�F,±W&��4)�wG�����ݠ�׷��~7,�6��ۥN�ђ�+�$�4��3�߉%;v��-^^�	9V�8�_�Ŵ�'sy�N�5t�.|:䷟�x~_�xf���hb+*�FO�T-qږۑ'�K��`�x�6f��z��?�9v#���CT)�yA}�q�V&u~�}�n�eT��gn_��ӱy+�(��m�E��6����@���v��|~�c>����c�r���8Q��i��z�����_�h;�Ԫo�>*^IX1��z�_�������V�6f��v��x҈�]�b����s�s|�d��������Mq��m��9ݖꂠ2y���Q��v���K���cq��	�����8o�X��ϝc�T��o!�gIu��z�v���ޡ�����O�})�c?Җss�c�-UfYn�f@�G�cϫ�G���6�q��7�~#^�����Xh��:b^O�2϶:/ж!OJ��V�w�/�9ar�س�QGCa�t6�À#Շj=Xwj����\+sc,����+RL�2��}.�]��#���X�9�4�o��g�vn{;���ò�?+?��}�_�7��o��?�/��?�G���̇q|*/�%���� }' l�����o���O�g�����g�T�9vK��9�?O H��P��k��ʻ���7%K���*�����ø$�q`J��ɑ�V�W�=�i@��<}��VL����z�A.�M� 8�^9�We+x�ߤ� |,d�I�W��y�����Tj{�=��m��{��P*:KΣh׺	� �V�V��8v�zۼ��pd�
t����� /�XW�G�;˔$5�؃�g9Ƞu�r�=��ȵ����6=cA�uJo�C�jX]i��ߚ��N�&�TrZc��u�BhQ�r%���Y�H��<�4��Qn.�t�0(a���S�U_�V�D/���W��z�{�૬�b�<i�G������U0��~�J�:<j��L'NɃ2�3_8�t#eou�jP&tb�m]�({qG֛���g�F���,F���D,���� mt���Ȟtw<��q��_���VV�����?�� ���Z0�؞��ao�g�|��S��A�e���o�?�v�Wla_�Fl�c����.��3���|���65�J!ϑ����a�Բ�!��O����(����\����z?��&�p����|���6(Έ8��͚�O��R���%�>�����ے.����k��|@ݴ3]����w
GۥX"7��]�C�d��u�s#F��σ�!2
�T>2-Q��h>�}�y�mlˬ'�����A;V�2��h�TX�d!��zݥd?:�m�:'Kq���'��g���Az1-����tx��1��@�?�l+�Gt�D�"�_��=��='�F�ǿ�m@�em�Y�bI�S�4�,�W�!�i_�A��±�n�KΛ��u�(�*=hG^4�o9>P�
E�����ӥ̾UZ�c���Fe9�Ǭ�?�	}�����5�E�'1��o��� ����i�O{���mr���<�����$��v�uxB��^|Z�E�xE��j�|�`Ҕ��x�o��N}�X����^�zv�\��9�K]�26�i��[����B,���]gy��X�_D�V�m����V�W�^�%�W��y��E�c8��7��^�2NY�y��Y�M/���_����X�S�#ՏrʘW:��F��s@É��/6a��V(Wg�nK�#�v����n'k�t�Ť�3�}S����babX�U�{|�㶾�Y���ʻ?��{?��������>��?������կ �1/�%���4�Oz�������~x��7������?xz�T�Wu+p�pW���]�� ��aܰR�J+اIS�t�:v��}��GA�O �lh7 S������+z<ۗ%�� L���񉎪�7�e}e��m�#G�'��� �F��t��t^�o�W�h]1h^�u
R��Sy��ӓ��:,9��2�������y���]<�:&��u�'נ�y�o���;�����t�K���1�����M�����AA�{���8�; ;�:vY�M�~:#1t,�1^�u�ſ�Hƶ�9���\.ۑ���W�`��z�C���?8=��	u�������~K�t�g��@�o���A
��ߵE�
�y :�i���s��O �v.;��Ffy�6�5?ڒ߯��||��:P�����A9����Nk���1���:v�S�Z�b7��~_�z�}W�蓧[����<���Oi/c_+)��Qzl�����P���pt��h+�^�t��N#8y���]��:���f0�������a�y�0���<)�vIyN}LYq���`+>Ԑ�u\֟I���d>)'����������+�O}R�@�ʥ����e��^o�u�Qj~#y�X���w�TVz�y�����k�~���Nc�����]����zb�u��ԾDL���S�Tvu����q��λ�#�-��'t!Ȑ���y��f�V�X�ˀM\����|��R�G�V��IiK��n��[�Z}�1��#s�=���`��eG<�R��w�N�8������>�wц�����O �����sխ��b٨���}i_Vz$�Ĥ;���޾�}O}�4y��7ڿ�A�.~���_��clx�88ӗ'XW�����og#{Y�wWvX�~eK��^.������h�r�Z���vf����tx/�vi�>�����y3��*To�r�Omk�q�G��I�"/ww����gԭ[��<����Ņ�B���y�������nֱ.��W�M�L:}!"�d|�j�hV{�z�xul^(�X6T�4ncf�w5��.�yHԑ�<��n#"������c1�h������z�����q<۴�\�Uu2n���_��������<�Q�Pg9����T�626k������'����m�~s|o��Y��ݧ�?����|������~���W�_\^�KzI/�A�2N (����m�o[m���^���~��P��8H��J���F��~�OP��� rU&N�O p��S�3�9������s���2,187:�mLl�`�t��e(��$�2��aM�j����V*EÝG��:�����ݨ�Ј�A�����0�r�Wx;�{t��hkoiE �l��y��*��Ǳ9�VR��k��⭗��RKr�e�����c2G�9�l�ۢ�jQp�t���W�P��S�M���H׺:O踐�1w$L@f���G���lz���ȣAռ��ͼ��G�B�$��+�ѦǎUv̑Gi��#�)��[(���@`�g��b�u�|2>�V��\ȭOR_��Z��EtUF�?Ƞ/P�!��8)���(7�dȝ�ǋ���YԷ�����W���p�ҏk]�j�c�˸J�M>��Z�3�!?��*�&ۿ�Iߌ�(w��AM5�/����xl�5�<zyIc#�ı����X�_��g�pqa��e����Mk;� �5���]�*!���<�8�㏧�d��J2��%/�Hd��.^�����yr G[��I�OW|��@l?��vKu��	��XLʼ�ʔ+��u4ej��y��j��y���?���3������̴�pT�'��r�e>���rJ�h��>x��3}������k�6���n���v>`�Q������>��:����y�,ߏH�I�(W��&��ҫ�j�^��`��9��	ms�Q��1��7�y�����t��[jϺ�"��1�^�Řc<�s�k=�t���?���2�?E�yc���i��y�8��7eM���� ��J�U_�{�{5ycl���.�_��؞�s�/&�OD`9��PO	m^�[a׳�(K�U�M�h����{��o�cL#��mT����R�3�'V��m�]���K������ţ���mc��m��ݖ�t~xf��3��W���e�ک�t#�����*��p�{P:qm��ם����~����^��[�4���c���\��5�x�u�3�R���D�xX�D� ���Ѭۣ�vFD^�r��xmԉYg:��<���,��%�[�܎��Sϰ`�6$c���u���>Vn�wl�܋�m�L�9�]�7�`��x���a���� |y�}�7��^o^��uF?NOE����gf��T�[۾�?�*�������m����������^�KzI�KZ �Ώ�(�|�k��}�|z{��u/ۡ��"��8�����y.���� �H
z��qm���e��t��\xP��?{������Fp(���Y�D?^ݏ9�w�)��yRQC�6���Ғ	���]�VI'��	4�.�� Y TW;5�����N�;��I�(_����I�����Ռ+�)0�����wq��M����3��^H|s��.up28��7P{��ȓN�;���p8�~ud�+ʇ~��zp�V��{�{��̿v&�����&�4gǕ�����&�$ok,/�͑�8Y��&�pǞ:#�w.�Z�}�v:��XNn��X>��4)���sy��9�����|wZ#�h�(��C�Ɖ�O��_�����;Խ�؁N�𝷽��7Չ�'��^�x �MPJZ���1�����w�g��-@�	=P���O늋�b�k ]��oV=�&`��i�s-;�3{��0�����>�r�&[���Q�r�����u��'�u�:ޑ�+=��3Nj�:�7zG.l�J��~�nV�Eo��J�GS�:Y���Mmǖ��~.��QN��_�OS�O>b"��
���:}���ի2���%�c��=Q�F���^ۉ��?��<��y�[�W��өP��� �5?���<]}��B�ߌ;���p��NQ�I��_������+�eyllU���=o�����6yV�}�=��A7\%�7�7-�����gl�v�����P;��+<�ex�bG�O�r9Z�	�.���I@�����#���!����u�$����f<����/�F?9��O��#,�qw�S.�΋6�7�{w<����S�:�<2����l5�~�g�O�u����q��GRS��c,�x�?�^�j�=ַ=��6�OAO�}��c��}��͌��8c�&⅕��.�p�4ΐ�c���������H�<�Wmk^1��D_�o죌U(^/ڶZp���4`"�2G���y���:)�W`�d���;��l��I_�����kĔQ��P�{��9fma�g>1?w7��p�����{�9v�ߪ�\/p��6��*�����>��P^�#��&2y��3���}��"�f�M�$&��y�K�.o*��}�;1Vq��5��?�ڳ�/����o`�Q�y��1�O�e���=m�q"��3~+=�~��s����~ċz��X�l0ĸ�8Ť�N��e�k�Z��ƣ$NP��1����6NT܏�=c�z������w�������K����?��/�Š�KzI/�%���^ p��_�C��ٟ���������o|��w~��������\�.�p�p?ۑj �T�g�{��fp5��/�9;ui������Ƒ�p:C`gX�����h���	�p���}N�p�7����luw3��7�V�jv#�s]��{�� /:=,���Fm�:��C^�0���Nw���2d�,���@9 �A����"f��@!{m � M�Gy]��`�M��rD�,�^��-��䍰�Ip%Y�+箞��8�#��o��w}��� ?;���v 4��|�8��������\�Xg%8Zj� �5a!���1���4�v�V��v]5�'`]�ƠB=I�F-�O��̎�����<�OyW�����E O�o<]aR�N��W��ѧ�i�Gwf.Y�,�fMu$S܁��2�r�r��:�YN,+�9�LN3���T���u��k��޾j��������bԤ�����I��AMǷ���w��C���]G�t�,�[��l�,r;�m<��òc�]�x���G���=}�0���q=T������c �Iޡ���G����p�5��ϣ ��N��E�D�A��)�m�e\Ʉ���8V�@��zi��Yd}��='�˱S�T�SZ�~z�|�W:�Iu9�u�T^�ȇ�[y�o���~�68����KĒ�c���m[��yP��zɿ�UJ�a��������Ɂy�}E�ZUl�$�U�a��
���E���ئ�۪)/jM�1�D}���+{�ȅ��ϫ�o���I ��������m&�k�P�7#N�SP:�~���Mz��y<�x��=bub�G�&,u���,�FgM���=��e��+X���t�PF�$��N��c���k�~�O�鐍*��>�cr���U
&�շ�q�^�^K5�_b�G��u�������)�G�!�n��u��"��/��!g��-�P�^�a�'y�i��d�F̣�\i�������*�ǛxLUTh�
����?296�oϧ:�ݘ��T/��?��\\�qS �hGF�E��j�a��kL��m[˭L\�NcR���=l~m�%�[��������'��U�+�'ʱ�[��Z�',/ڀ=�g��m,��~������7��7`��<�������m�ݎ�����QO|*�;��:�D8���,��zIp��\�:�s�*U�]�jc·j���u3AԑX��m��I�\B�A�����dZ�-ᑌC��.%W�Z�1%���xֿ�v��x~w�x���mkEd�� b�A�gMg?�#��4e�����϶�Ue4u���. Ҟy�3����ig���n�ꫴ��q�v,Z8�~n�7����?�w~������r?~zz��������^�K��e� p�_��'�����+��~�;��_�����9����v�@''��1ЙW~�o:$>��^�zV�O�8"�R��AH�b/�n�� ��T��}s��/��(\vӏ�d��Pֆ�ȳ+��x����DZ�t���n�s0�NJ �ҟ1��{���&��#T��(�[˙]
��.klj4��+�=(V&m3�h�zK��W$�b�
ǵH�d�&�;=��IǊ�>�� ���X 	ΈR7�� �; �[u�,Q��|��6ױ������R�B�9A�f�`�������}W� �ֿ��Mtu�N� ���~����}��>�&�ˌ�jוЏl���6|�䲵�ȥ�6)��K�?K@ۂ�>
t�3��:�����퐏6m��K��*��١^a����R�u����i��;����T	����*n�:���j��A�I���!Ӆ�l֝j�4�j��6!@\��NC�n��4�A�\�'���}�U݃&7�1�.啮�>�	w��2K�v>�'�l��ٓ��w= ���*�E^��.7�9>&�ݑ�21�ŗ��X������Yn)�~_@00S��"���vS��)L�A}2c������H�J��aLi�ҡ"�h�6���U�Y_��]�E���N2u���5�~"��`(��m�!۽�hó|�>Uk��2�U��2�(�_{���3�7��7����/J�1�L�q*��H2���hi��L���	`�%1kY{�����!j�FV:���O-���	RB�#jU��lp(��TuG���_�"ʤ���������]�1Ug�j�G�]�(��%��zy��	u�q�NU;�5�2"�����89��U�4�e�W�VQ�ƿs���8c:ړ�Z� ���Rnh��M�9��Φ5�7�A�{:��;��gq��|M-ȋ�4�6�ǳ�I�����'=���A�����7@[]=p�h���tMZ��.CCȂ���U�ȷ�S���شkD�al�-ǩ��c7�-ت)o�#�4�lb6�:��.X�4Ї�qA �1��;��:%�۫go�����11��w�aQ��i=š���L�"��xUx:����cx���s�9�5�R���u8t"�S�g{ʺh�d\ZҒʄ��k�+\۷�W�'ײ�I���Ք���`��>
c��=Q��W91��y������S�G��b�IS]��¾�_CyP����.��M�`�m<q���v�r���:�/�'��F�?���0δg�Xl'�m5��r�f8�Ίf�k���N���ͽ)�9��݇>�������~C���K=vt��g�b��.3C����N�R���bd��9�Bl��/5��c��yc�n�雜0	-O���sM�����_�_�Ձ��\�O���}㯴b���.r;6��r���;��	?�a��~�@>Xz�>6��1�%��1C��s1������r{����|�۟���'�����'［����?���v�����^҃�] 𬸞uY��>=}���W����̟��_������|��������c��O�;XWCໜ��x�������D$�VO����� k� �2��U�e:jNk�N����6�9V���ͦt ��D)����~���qp��E�4%��Wܩ�u�����V�	�twߊ�0�?����}+��r�W|j��SG���� ��H�����D �K��# H~%�dMt�6�G��T�cР0h0����v���N�X��Х�Kg/�8Q4�J�KM��o��Z˲-p0���T���k}�d�M�wh
Sv�x�'*\8諡�@G�X �'��ߕg�HOX~_%tW-�N]��+��<P��X�ˡ��710*�'�?�����=�F�H��n��6��fPf��A?�ѓ:����r�M���Z�n�-ǝ�륪;3�P�w �m�#��O*h����n���e�>���3�:�s��B*�R+^#�o}�z\}Y��c�]��@Gi��L��Q���̆���`���ǉ<�q��&cd���H��&���)�9m�,�y���#��T/����MO�A?��Q.PW�j��W�w��I��;�_�0���5ܑ?�١��jюJ�5�@�ƣ�K�� |�6\t��3Y7�Z_M{��g�U�r�Kc��\N��|�=$gCK��ٖ�,%{X�� ȹ�4Em�Μf���}�Aqt�H�6��3��Y��:���/�Y�o�����.����`|*u����ۍ���8��9>!o���4�@+���"������"�N8�jS�8���m��
a�ob���#\9����\4���˦=!.$ox8Y��.��Ru�&�Y�fo>����,�S�پΡ}>3��]\(X����k@Dj�)��!�xo~���mB���)_+�f�f��J�&�"r�J8��>��fuG�Fqsc�S�ַ2�{9�p�Y�MC?�<�}���ee7������;��<mt�tH/m2�Zy^�d�+��&���*ɣ��S(K�'�<bq�ʹ�41o�'󢅿���H��[���n�[+�������׫�Z��WX���hh�ڬSg &zZ��,m�4��)}�s�+<�>m�Oˌ��6A�^���X��lL��;f	��7S�߅�"1*�e����������|J9��]���dc�[����;����& ����Ŀ�`(���FF���^N�s�J]A�Bf������礮�9�Z��ط�����W��x�D�0�rN�ˢ�P����5��-]�G�G[㱷:��펈��h��TP���d<���h.(ڢ������wO�&
f����=�eU������U\幑! Ի|7�z�=�kQ?�Y~H��5e�3��1���m`�z{��i+�>x������?��Ƿv�����k��^�KzI��9�}���}v��'���?�͟�����}��������N��cp�a�k7�
p���ܟ�d?���?�������K�=�d���y�#�4$�F�Uv�Q����4ܝ���e�#���ĵ	�:�f6�FMWjq�'��|����)�<���; rڬ�3�M� ��G�����s�(K���c\�p5� 9:[4���X�{, �kq�����^xJ>�J+��zq�8���:�
���e�3�<t痎#�M��؄��Ǿ���Q�7���z��{���U���7�t��]������[����c��lC����N�fG^��^4�k���E�(Ԝt۫e�1�� "רW��>tyqDG��,����(����h��-��':
���ע��������~��S�_�3�,�L���c��Nڥ��gԵu�)�
��|?n�z:��w�k 6��.���Z��]O�7�&_ub���>ɇ����� b�M]�R�m�8i������Zq�u2�l���~��ȇ<��Y��5t�z�4�C���*��)w�9�k�Su&߂��`��'%�w�Ӂg�V�Eh�7u�޲Y�b��v�8���G��־J:c^T|G��"��q�oA�W��sr��n�3�(c�m���m4p�;mZ݆�N�����8��3���s]>�9�'+�M!o�
���y=[Hk�%(;̳
Q%��>�C���0��9v�f=��e��ڔi�]_��I�@U��'�Oa�+��0�R["����DKi���C�W�Ǵ�y�!�r�5i��2�k�� i�:��O�q��>s��a��&�Si�sr��A�hkS�Ao3^�-Њ������Rt�֒���l�lv|�BJ�Zu�Q�r���񁽯��2Q�#&	�}�]2T���l�����&���"V72(�U�ʏ����!��1��&˸�:pj.˗&I���n�D_9]�WS>�����%3����ۗ���ap��|�W�E��֯�q_Mub�zj��߰��]�8&1�nԷ�.b��E-6^�w�O����ӌԟ����/�����2yd�2��t
��P���w<'�Pۙ�3)��W�ɓ�v˸J~g�j�E�]�z呦1'�ּ��4yo�O��4�3�k:VD� /퓰��(��'?,?c4�۴?�Ge��2<�n��J^ہo+]���m�=2^�1���#
��?�h��w�|R�_��N�B���|p�\,ﴥ��c��)]M�[Ș�>u<��~�PtR=���l�.}ٟ��#���)8k�k�^��'���>� �8�]�B,��Ѳ��y���il�X��H#I�y���l\���CU�餤��|��6��E��:79<�܄��y�ƻ�<4�l_!���&߶0O�4Z���@��F�����S���8���Z#L,4��N�0xv���׿��׿����le���/������^�[�/c@y���m�ߞ������w������u�q"¬�m�~W��'�E<���~?x9��9�{*ڝ
��3�� /�*����pb�'���H����0���XT�p=@9o��&t��0Ntb�99A���;�i^L^��h0�� ��x!1hP��U�ufG�$���D�SjЦ�^��7�Op��~e��:�V�]�a-�t
Ž�� �\ʀ�zp�=�!_�::��w2�J��]G���K0A��Vg���>�8���RJ�(��]����Ӏg��7G^��ᨒ/l�ҀwL*W�GwH㺂^��e�n�g�F�����O'䎤�pP��b ��Eʔ�"�{���o�GkǼ��
�;�y�;ʟ��^L��]�p�|T��_�!^��c�u��J�@��z��KYu��˸���X��b����KЦy��ʬC�!g�p��Mh_�s.�S�T����f���d�J�P>'�خ/����ڞ6����6f���G�u���J�6F]D�Zq}��S�zU��Z�����z~ߥ�cp,�v��Fο6��ἧ��Č�<.�+��<Q&�	}�$.��/tb\�v�4�j��p����Y�Ss��ߠ�TGy=�NO)��Qw�o�%*�N/��b_п�oK�!��2�����1��3b���j�c�Q�6�m~�������w-^Q�$�h�].V*�5B.�_�?[��u^�]�C��>)�~�	��l��a>T&˰U��?.J[�/�(jeb��/�k�k�K�+M�O���x �*�H�qB^F�dXqioS�<j_�W��w6�6��j�L߼*~������Z�N\�V�����`?���u/�c��'*�K��~���\,]��a���T�!��}!A�3OL���3�&m3멳���?��8�j��h���s��
�r��xKy�ر��	ʏ�y��q��{�a�/���$5a|D�v��J��"�~���y�}!��cB(�v�"2�)q�� ��^�.eG>�J�E|*ϼ-�;yI��|�?��	u�
�h����З(��}Z�4\�Iz��M̨e��Evmr\�6����m��+������G���@� ���
�����p��h�<Ae�������Fu�����Q�me!o�~���z3�R�J�⺎��)k��d�Mq���Q�����4��*N���:��SҢz��9�l��(I#aC�٢Ť~LQG�_���2�G}?�O�5ʪ���-u�*��\N�.[�6���oe�l�a�X>In���ҏƅ4U'N��#'�`��ҟO�k����+�e��3ލ��!~��c�2���ZN�:�жS����^=�ۧ�޾���z~���Y�����^�KZ�/e��S�������?��>z�^y�����T��Q�	��j��N��S#�2/y$�0�U�mDdF�XE�(����}����|2�0��}�=D�@���X�
�&�hy��K�QC��ҪN�K�9~�=6��^9.e~�4�R`���K� op~�|�\�ɶ�;Ez��ϵQMi�ů1��
gd��}��f޷x�ֽ����L�:y-�R ���(��ɖ*�`�Z-8��ʻ�z�)9�Ǆ�e��ՃX�S����� 9�o����?'������H��C~��Kݥj�	ŉ=�u���"�����ء�O��2� w��	 X��Uޫ��;1F���Nx<;��U�:o�)d�=��i}g��d�V0A�����8��|� K�:�2�H۝���ӑ�*��G�k�&�E��)�����0/���>��[�����e�Գ҇M�*]f��0Xg�ڧ�g��=i������f]X�����R���&<ՆAvR r�7��*��Z�B}�F8ָ{y�|��O��JVuT�sm�������q�����V�)���WEW�X�va���x<��}���ƙ�6:`�T�RL�u̟�u`���:&��3�0w+ı.����0����YsB����u:��;GޛL�d�v���e��+��_�.�n~��B�X�x�Y^���F������A��J��G� 2�N�����dZ�z|�,�h�4��zR�ǺM�������Ra�k�3�PR[LAk���*�S0�E����&(+b*����$Ե�7�gu�h~P}��:;s�����Կ�GJH��إ4��Vbb�<�_��á�&;e�s�����8���m�
�c��Gǰ�(�o��Uo'��r��'Zǻ:�����V�=p��3��F��}\�4ii녂�i��'�sq�&��ٽ��;��������c~�u��/7bw`�t��7��lc�oCv8A�:�?R�U���؆R?L\4gm�0`�6��.#�E��z���KJ���ܪ|L����X���p\ej�̴~�!/�.!��������ޔzG�Mhp������*�k�����y�R.|��^E&�-�&��E8��S��J�f+��O�Ъ���o�_�M��b��%��|j�l`�xᶱ�N��8�����?����9�l�<9Fg�܇6Ɇq)¿��y�ִ+m6�ؿM�i��_�_5�_�]�������J���ܸ�|+ڟ(K�jx?����rd��I����60f"���i������ԡ�Q/2�l��c�0��Aܔw�������'i?��z<Ǘ4>Ы���+>�X��w���RZ�0�6�w:����r����6,��9��u���XeS00@}�p�b�S@vݟ��7� ��b�>vq� �>N�-��^����o{9����쌗��^�K��e, �O�=}���������[�ϻ����~���ի3x��Yy�G�1#A�
��U�j�t��% �ap`d��{�^ݖ$=(r��܏�����]6m����d,f�̐�!�� �����%� �B�d�$�� ,fH Fj����mWw�ǩ{��+�����D��oy�;a��g��V���Ȉ'>2�e��º�t��o�]�x�/!Ͻ|�L
葭�����e��n	�nTJ�MW��5.�
I���E�T�����Y�c{V��p����d#�b�7@Nw��|7��R����2~ ��s{���ԝ���,��v'�--q��YgI��Ǽ
"ȧ��F��fP�=B3<�x(�����90��	�#��r���c��gw^��UzXm����V�wd�j���%^�5Z��-� ~Z�;�;�W���j�9O$/i2B�A����kGvE�ًw7?��|�ٱz���VGQ����kWu�RY�nq�[�5��}g���9M's>�T-�6�6m�ڶK��:�D�♵�!�9�s����/�^Ot�䎏��y&?��=��zo���6���A"ck"3���h�A4���'u������]�0nZ)ׯ��S�8T�`F``ɀ(�8�s�gL[[Is���c69��ҷr�2Ǹg�������C��r�y�8:��$K��֚�jC����5^qN�#}��*S��z�"�[I��\�:��s}w�ǰ�����~��}l1�}����c��{�I�'�<[�ifK6�XENt��|����|b���L��+�P���s���5U��vY�m��"��ː�(Q�@�H�8�B�!��	'��coC�#��=��ܦ��8�9
N�{X�����6�Դ��-iv�H�l�Pݎ9�c���5��A1߼����ou�N��C�@o�~mA~�\��k���&|<.�pL��r���wg�㘑}�n0���.��Xދ��hb�{pvZ�C¸�{=o:��ܺ��]}��T��A�5 ط�醋�7IQq���@���Є^��q���V����kt�����i� z$�'>
��<�$c I��@�,u�;�<�y/:�p�/qF&�U@'=���H5-'�������:V���{}\�n��>��4���.�%�k��9��s�'��3���L��9�7v�A�R���32kV�
ٮGA��u���-G�Ř.;�OVi�1el��ߛ�M�`'�ʈ�')���s=i�X�-�
҇�����_I&���u�8�Xe�}9/I	^��P��8H�B��`��|;X��`�<���<�,�ZZ7�+�1�`ہN��팴#�;��uwqO�@�YTl�d����Ȇ�6K�c �.���>/�N�3�r�m�OVp��#��Z�Ů9��63�����W��0І�[1�C]g�{�FЧ���[�\�`� ��d���I�mlO�؊��"v�|���hp��﬉���qm����~�\?�'bW躭���@Σ�-}[��Gk�;��}��������ӏ�#�i�;�fJ=Zr��F�ۂ��ϻl��uo����y�O��FL�8�(<�S�Zy��-���T�h��>�qr�:���ɗY��׵ ��__e��e����7���'/�~׶ju�v{���;��������M�K���V|D5��k<�gr$�`�~�g��C>t�����cQZ��Z�L�<�4�z	�},L�E���yA8��/>�k��_������o�+�_��>������K	�]o������j��z��y|��_��?���_�s�����}j��#�[��y����m�uw��_:�T���l��#= 4��� �#�-�Moe�}�S����8��|}��Y��g��h��y��Ʒ��{��F�KP��d�߻L51(����(i��<�X�w�$��3����? ���l��aFY�g�qd����zFK�����2�u�hx\A���(i�G�����èwf;�?&< ��e�0���m����x���rr4�p^t�w)���ҹ�������:��O��J��x�>����V���`��d��WA侖��UV^�����[��=;�|^�c[��/Ըk�"��G������6�&؍�ܽ��m-׏w�]�
������V�ڔϿ��R�����.gk�X���2�������z�x3�vZbx_'��>f�{�Xְ�A�Юm�8_�>�;��<0�V�Xcuۃ�c�!���ꋝ�@�����f�Kud�Gҏ�"�m�����){ϳ�#��~x|�;>���K�Rv*�������]�ǫ߬X��:�q��e/;��5�-�p|T��Y��(VQ9���P;ϲ�T=��Ꞗ���s�����`mk�Ϥϼ��:�t�6��ʻh��`�W��	���>h�˳9�\�W�s/DM��H�A���C%�߲��̍@wʩ^������:��ݣ^縔����gv����Y��+�|H '�VU���TV�z���-Ŏm��nv/�]���^߯s�{�'� ��T��r�&�Q����7t8�����v���D���|C�Tv�	�H�<�U�t��$f�|�ݶ��|�Q�c���wm�/��)�E�65�o�i�Xu�����;�m���#[꽊5���o?c����qP7V���V��{�s]*rm���ك�M�P�\u+���T�8~��Ԫ�F`��X���e��n;?��2�W]������?u.�X؉�<^������e�m��q�.�w$���y���\����[Ƌ{������>�Qu�^u��^�J�!�|�B7���U琯�u��۩WtmLy�G`(�7Iaw���7=�9�������$�G����i�R��q}x?�c�wG_e�=�c���ƆK��eT��<�]ڱ,|+5�î�Ue�>G������cDm���\8[{�+u�]0@���W�0�>��nWlT}a�n�O��4pLL�����j��v�!tB���5��Ե�s�I�G��!+�X����+�ǹU}϶tm�s��4 ��]}׵C]�>��j����~�I"��Q�FU��}͜;(��Z�۴��뚫�R�����;?�ɣ��h��ϻ���cG؊ăwb-�$��Bu��&U@�ņ�m�	���+�;��bʋ���\����j�-�hP@�t��+�4~�0�k]�;,��/s���X2/���������[����џ�#���?v|�}���]o���v}���T ���OO���W/������>M��h��b����IwS1w�F1!��HƦ�`���t����!�� �h��@S@��w�W♖=4.J�.C3ϩ܈Ӛ�#2נ���0�s�H��r�c�^ϖ�zWgB���Th4�Ԩ�9�8+��(����i���
���B�Uc��u�σ(��ⱪ`׳1�Y���D�[��f�_��O���;f�4�(�J���N�����+��PZ�l]��w�>�w9�5� �K�<����x{����9�]�/���FW�Og���%�w>q��&W�Z���X�Ȃ�|��tg���.�"�*�4㜈���|�����*ƺN�@����X�3��B8gtm���X��#Z\
�����r^��; /�e}-g��w4�ϝ��7��\?�,��v-9sූU,pЏL��e�Ȯ��>��J�i��wP=�ot����r���t��<�[���cY�����:Ncn���o����V��6
勉7w�ǜ%}$��1϶���o���{���eI|�M��<׽��YY�{�4�?���=e�4�(Y�I����%�2�m�b8%�pt�����b�8��u��V.��e�U�j�t�������Y�U�YǶ�&�CǓ'��|_�XH�9��d��㠞�������>5��5��ΐ���6����k+5z����
��O���h:�=�a�痱���Vq�,粥\F��{1���M�~B-G�ܚ���K�X��O���{��Pe�.�^1/c����?���?��DyGȭN����/Or���G������)�^����[����pܓh�6cnz�7y_t�,���|?�\yw��� ��{���5&8c�>xĹiG�\�[���,�+���!�{�ܣ�,���H!q��.F�g������|.��aEϯ��wgb�.m��X�gqx�,+�����.b->����W3� 0�$trb�B��8
���#�d���fG�%�@ŷ�+Ig��2> O>da�S�?S��ĥG���e�Ux�n�P�e.m������-��!a}�:�F�T�KO]c�m�����>�t��p^�:�*v{�D���8i��M��#�E�B\sщ�9�N]�.��ݑ;�G��	G�2�c�-�Ce��.�M0�ߍ�-�sOO�M���F\�!���e|�>04|Γ���N��:����uor,����K�z�oX8�y |~L�|>��g^���}�t�N(�o���vzzz�$���>=��y��]�@p~�{K\^����
�x�/����w��I�V���g����ʃ�a��ௐ�H������w��?D�O�DL��_d�n�.���4��x��&O?���-ʜ���o&1�N�5�*Jô�k3��_��7����k�v�l�>�2z�y7y�G%��w@�vp�>A��;�=�-K��aD�D��g� |�Y�-�*¾F�j������m*��ڪ݇������{����;�W�u�'	���L�}��3�&zv�u�<�*��I�u �1!N���C�qF�=��}.Iמs��ۚlu�O[��^R6h��՗�C�8D.�~z/,m�? %�]�Z��n"`n���'F�1�}�)��F΁��ߥ�mFȐ����"�I�#�x�˄��ب��}&>�r���fiK�6���X�C!I t�F��"��p_�L��m����dw{����o��:��wϼ���˵�������3r�Α6P��#f�}���n0����U/B��6-�am�.6��N���c��椁ǆT�H���n/�9=���>����?~�w�����o��oM�p�Q�v�]o���w� �����O�_��ڗ>�iD��
=����@�;-�S0�P8ȖC
B�����P��KZZ���;��dB��,�M�ʙr��D���a�V�D;���]��⪣�P�vb���ʊ�
lnM�\-�c;}kϕZG��ܸ�����ߗ_~n?��oz�M�I�[f(�Q�z��s�4Ҁhun��β���@����̘]� #wQM)����i�4qH���s���K����Jg����k�G�[w����[;�.ʃ�� v�Pi��6ywp�5k�s�2�VxC���ϑe�hTp�b���.sm(-���#��;��]y��>��E�T�����Fw;���^k��k�n��8��T'ٸ���e�}�X�x��v�+4���=ud�����~g�qy�n������J/\_�/J��Nw8_��
5�Π�U����y��C����,ec�l0���y:$w��>q�S������1k��� ������z���c���8��ּ\�k��v!�{���:R׫���>{5��d�k�އ�y:KO-'hn��Fڌ���	��̏ʁ;}�*>u��]w�ꮀy��`_�w����mj�{����w������:T���{I �ߩ�km���s�#�v�#����w�nM�����Y�!���Ft�}�����m󎉨���?��Z�A�($��{t��`l��񰜯]G�������NA#h�Z���9-Ǥ��ʣZ%������.7Mڹ�jOI��7c����Xq��Ͷ>�&������^bO<�2#���g�߭C}����{��9�1��1�7<�r��h.��*K~յ�����F�^�y!S,d���{�?�J���)���kblw2~�WۻkW�箷�����86�w/w��,��=��}B�J"�E����e��:}�C�]U�39����Vۺ�J���z�x�.w������rG���_߆v,q�/���>�v\���v�l�6z$����.���e��"d��x�p�m��|G���"溗��|'���;��1�>�;�|m��隨<�|��@��ެ;��%|7/����޹�㾶z��\��ɻ�:�Wy�}S�]���׏�EZ��}y�>Jǽ��_u��t&����!���?�V�>�33������v+��q�As��sluZ_}�ιҲ�M�A�x�c�3��.�����i���ß��=??��ϟ�Y�0��]C�n�r����ח�����N4k���q��8�Eð_��//��-�Y�(�I 1�٧.I^�2��s4T"˷1q�㖍��~I*�,:�gP��;�q���,�\���q��3��J�[O���}������ӻOϟ>�x�܍����z�ޮ��. ��?x��?������7/��Qnw9s�3�!`[*�Չ��� e��\ҐAnC�� ��ٓ@`fe�]�p�;��c��m����T�sL^����o�hL�*����/���
�]����*�!�+�9�P5H�8_��A�O��_���>��������gޢ��	ͫ��=�	�sT� �Ap����Mu�ذ�ǥ��RG���^�{�����ߑN����(k	� p�w� w��~����Md��B2�a����	�XK�6�a �Σ8/�P:����"F  ��IDAT9jɺ~��e6~5޵s��䓙�n��}F��P�<���yz<px�ش�lu��Ұ�jdg���$�������G��o M���F���aY��3�u�sGY������bp���H�а��v�,~[;�<�<����Ĺ�H�̃��eb�U�;�u�@?��L}>6�x�8P�p���<��4�i����3?��<����v�s����vp'��������ߝ%KQMa���a9�9����C"���m�;��a�Ya���'ls��;$u�;�9N��а���c�{�6��q\xW���~���X���0lF�Qu����W`p�������r�4T�sV:�6�5�E���.�̤G�6v+��^IcصϾ�cH���e����gw����>��<c�ɔ�~����D�]��Q]��]�M�=�݅Nۿ�dښ�7��@�J���Iy�"��s�4�,:��a'f�uRp@���;�L��Dd�Ơ�r�a��__�9��wZ����;�����:�oF��ǖ��f��2o"����8w ��\�+�dD�w�d0�4�D\�N���y�I$;}�{t*^�_��B�[���v�5j��~?�[w:�rOu8/�ݧc��S}π(��Q1,ڷ35q���2����؎�vsu��:�3���>bȯ9��𙾽�4�i}hB�޻s2`%��Y�(
�+]�)��
.å�P�Ee���$�h�{<y��y�"�.G��;�d��U�D�|��d@f�q�l�L("�����YV��r|ּ��,v�y��#�1���臉�
�a���n�<N'd%0�0Z̍�S�>�l�P�i�-}<�xD�Į��q.C�T������P�E��N�#����oP�ʞ�=���/��jR�Λza���oM���D�Y��]���$^��Ă2��:G�3QM�.��������~�&��wıs�
��֤̻Ě]�_���c���2��W�m��J`6�t����8��}��ދq�s�~$�sK�%��+�H���Y��Ef����<"�,�2�[4���}�S�]��'�
���Y��: �	�.�I��3�d���p�9+]|��ɴ��4��ݦ��M�ǟŻ9ms�ך�#���j3���Vת9=��5�n��q1�#mB�tV�{�>���k�+^��t���e=�qX{���{�#�p��I��(��ae��	<���ԑ��n?~�h?�����l?~�/>�|��g$��K����q��}��=9��ҟ��l��,��~��ׄ��"��۷��G_���u�]�{��-e3t,l�O�q4��t���6��L֮4-|a8����.���n���������g�蛏����o>���ٍ�|�ޮ����;I ����~�w��������/~盟>�����gQ#�v�JC43뭂M�T4�c'��c�J"��T:-��y�8R�J&���@��ÍVn�Fw�N@4�Yr,�h�AK�)��r�Vo���*�C�a�w��B���{�'�g
�n��������_.0��bt��G?�/��"��Zf�~u�x	�:����T�UG�ʐ%�;8t7���w�Ή����-�`��9����@�9ޛ����h$D�+�{�h�S�bp�]b�'�e�tE��V��nd@>Ey8N�#w^�]�d@џ���p:} �_3���#���<����<�=-�Q�h�Kw�R�g��z��2����~��@y����W�(�Lͼ�_�]�#dh�� �]�p�6io��c�u%�n�CC�>iy쇌Wqn纆���P��%-	�A�aU>�#'�|gkHF�pnE�̩���ɔ!��zp�kچǹ�cźA���p��N$��8`P`�����y�� X��p�Ji�vW���gn�;�g"��Ek��B�}9E�{�_>����x���-e�	����4x����P32��^�|���n@��6�Y1�5���r�>K���禮j��<{έw�yr���w�#Kv�F��oZn�Le#Q��P�>���>W����{��z� �`w��b�Q.4��^.����s� KB��_ë5I��H��Z�1���#�)�v�𵵖�I�¿#q@vEx���oQ�9���)ϵ�¢^�\�����!		�/�Z�CG�#:Z�a&����)�A犉��8�=Q�~����
����k��5i1u���#�}� 8�O9�ę��=(�2����G���%�@�%OqtR����s֚B��$6� LA�e?"1���a��1q�A������G�r݈~7lR�e�N�&���<X}U� 7�����&��xl����dBI0	�%�7X[,�˅�J���,O�)Y�jې��LZ��O$��*1�YZ��y����i� �od�ȿ�^��Y��T�k��X���r-/a��-#n��������.��+�C��js�%K��
��=�'9�(���2o.�6��0Ǳ
�X����c�b2��Hԧ�qyO[h��C��m��Ч��\z_ʾ�m[k֒׬6hQN����,c-���A��|�_4�k�ӹ�zD�q�(
,�r%�qb��|��bc��p@�s��#��09,�-�]��{�q%�9���=O�C7�_��2i#h�2�+q7��{,�2�J���_םQ��$���ï���Ď�9���ȃA��'��+�ϣ���x�f��Ҟ��Hr,��jW6�c��C'��4�����9���\��,x���Go��x��<R+�7��c����C�'߭����D�N��g���a��Z�� 軋�'�ȄEuMp�.1�u��ذ$��j������2a����	)pW�jky>v�!�ŤI�ti�ACv*Έw�)�΢�uD�����<_Cpl}f�GE�s���2S����1����Fx��䃞�l}�P�����;Kљ\�s�����3P9I�
|���k�?�/B�4�ݯ;�T�D�u#��b�|JŚfC��	���`�c-|3��U-Fe��P��r[�w�t�?a�rr��=�Q#g&Gßr@w�n�=�K.�~b�����(����b]�Zm�Ħ������,����~n>|\�x�x>���/��g��[�$Y��U���SE��M�� �`��I �])�I��B�ho��F��xE���KFM̄����hi/-,��8,�ƛ<��{m�ݸ||_{�������z���g����������o|������冭D���v�]oW������׿�W�ܿ����������{��_��x����E���=���bt'���m&���#�X�s�%�NYܗJFUӌa8���
M��G	���M�v���;ˢ��f.���q����A1,b�s�j��X��,4*1  "�%@�z�N�Ucw�������̈��7����z���K����~���4�1)9T���r�fM�����P�,�F��IK���)��XI�J�1�|�6�}��F��&�#i��`|�#A�8�,�6�%����|oʗ������l�;O7�9��T�`�8}����)Y/�Lh�VO�A�.��t���#�%�V��SPwՋF�j�E�6vu�j�;J��we��'�V�p�AQ$����+��x����t���17~2�~`>t5(�G:�Z�B��G�c���>d���Z����KF���ѝZ�&e}G�c��D:�.kǢl\�Q�w6�.^_W8�X˘�xndذz_�3�裖����Y7�{a���f0�� [�uXh�h� _�&�=�.�|��]�-�s���2g�d>�"i�������	�Qٶ���>G�n�cF�3�$��p���ז�Ny��3����&N���1��H���#��
"�d\_�c	��#Ý��}��
���˛)B����;�=A�12Y���;֢'2@U�i�z���1gw��81�q�&�'�i�bwE$�X��G��L��^�8��Q���[Ɯy����+?w�`dY=\x0Q+)p.7����8;6�6�rbbP�*�Ô���SVS�*q��V��L�a<#s���@_Crt��_P�T���r�G��I?Li.J2)l�'+h���9��&u���у((����|&�NE0�{��0kk�,�ov�8.��x?�L�/�\�h�3̿噡��a<��@�$4&?r=b��3��o!�b�8. ����$�β���}b��U��w2@BH�$�SR��V�������/գ��3�Z���G�&�m�̄�F" ���&1�~�h2�:�)O��[Y�������A�fĴ�	R�l7�y�|�?�쮌��dW�p=��2ulI���F���j���v�%2�F��o��9P��ɐT��G�&<ɕ8�34�_{� ����q<���b6ᑞ�se��ѧ�u܂��`���#I3nzf1�L����r:����
g+�VtD&F�ZV���v6�I�a�߱������B+o?~?<!+�o�Rp;!�B�t�u�D���%�Bގ�Zʖ�T�w�r��c���r<Z+}>=�4 .2��I/ϳ�A�Ɍ�w����P�w���5�M�˴�F�"uY�38����N[#��:Y�/+���(g��7��;����*����ەe�{��d-e�
"�������w� HK�\��T_1T3ce����@�:f�+؞"����#�� /a�PVU_�Y��RF��nٖ�q�߃]-y4���Q}�ہa���j�7И�ދU�*�LXյ�"��0�z>]��>)�GE�s��)nc"�(����v�3�Đsm��<T0m�7R��F�>���+�h��M�	V�m�,*$*���E�ɼx{嘃��^2C%.�C��#䟅6� HN��0�
p8�7�9�$:<�F����Ae�f+�+�߭vTG�~v[&��\qs��X1���������2���m�8IU|��.&oD��+�����E��$�_��_���c��Ǐ��_ӧQ1*ޯ:T2��b�^ܯ��R��3�*��y��	�c�>��V�6�'�;9^�� lj4�u B�y�Z���ܟzd���!����܁6�h\]�Jf�T�/B�ׯ�q�W�g��g��?������{�����o����׿���޵�}���� o���v�]��?���9��z���?>�~�����;��������O�8,���:����_��f�[�5Wv�
 "�}!}0WZFT_�l�/�/���3W�O��z
vy����� �S�]��4 h8����+����P�F �lι���ӧҿ��)�q�4ъ!+�3���}^5��{�_ԸֶX�YKmi�^/8@ @u7r�[x��R�j���X�Gj�l�8����'h*v=�rйg��p��1�����d}�~	����:gM�l"|�,K�?;��Oٮ�R�M>Gy :i�9���<�* �1,���G���[����ۄF�����&^pL�_ܵ����@�`�w�2���q��K#׹?? ̅��1����i�Ξs�췥���\��L����������O�s��K��ҍ�{^��I��Ms��/�����g݉!s�Ъ(�<�{��Т�lx��n��ב�`�
Y�o���??Wy�ױ
��n�9��G��~Į'M~��B~��r�q�~T=`������;����<�0�:����3��Ht����7&1`>ד��O�c�5�D��0\EN�>1>.��T\}ʒ��c����l���90��'3��X�F�p�Ȧ~ȮK��2g,���;ܧ�Ÿ#Zw	t������<�2���c;l�DC���9V�	~7I<2�F���������}u����N��ӽ��4��\F��DEh���0��0�)�|�t�'����p���j�*�J����q�Xk"�(0�E����b �u<��-bn��8܁�	�7#�}>��\V<��@7r5���ւ�z�Q;v��F�V���5���6���T����D�1�oo�v��w��bC>��*�\���6�=��}v�Ԝ-/0(oYsգʉ��6������̺Li1O�cF,p��ϝ�,]��O!��w[�j!����H��w�M2s~暨2VB�ƈ� �x�$)	�R̒�y=$���wSc��%ݍ���-_��j�y 	:� H���@讬7���&�[y���b]�ر���:�� h%�����p�� ��A_�}�қ��"2��A�o�G�E������r��zWjX�ėg�Zj��h�An�dW��C�R�Yw4ch��#0&:��5�����7�g�'������f*��ÑX5�M�#a-��|��c0o����`�7v����'�i�������{Le����{x���פ�D�)�[��Z�1�����wk��LD�?͈=�������G(��-fLXԤm~��4��+�l҆c�s�[�.v}ח��^�o�s�S(��R�+0����bR�$�x�H��8O�Q�����*�Je/��	6�y�j��H�_��)��*:ֲʀ�(|0푺	��f�̧���y�pr��Xt|l:�zr�8[��&kK������8�Ѧ`7�4RǙ$��/��d^��y�(8,��i�gŘ�׵��3߈N�],`������ޜ���Z�l��T�����`U}noC��7������ໂ��t�eh_~����0+"�g�ӏ�Q=R���}���>�j�}�����8
��ϐ��k�[qj��N���������>��HyA�������p��Ug�~�*���f�uf��;:A��
nX���if��t��iV ��n�7�͏~�����x�������7�� �v�]oׯ���
 �̣�=�_~������?=����<>�kq@B����-�!T�-����4 �j��vC��J':�K��i�i(�#��'�e��Q��]�������ޯ�Q�qF�T$Hm:~�Ѯ��w�]��
���s�>|�F�m��lKv'H�_�Z��o��n�d�@�<����5�iW�ʹk�7�_�9���P��b9��a��^����
�Y�
�`$�D���}c��Ύ5,�a��P�<e5���|�-!y��Pf��4^�X�](ٛ��ȈV�T+���i�T����w��aɃ��v5&��\��&wϵ6!�ŧ��9 �k���>z�Y1��C���W�k[����j(�̒�f�=<��B�b�9 ���XQ&�Q��vcx>�F>B��0(�����.����s��*�zcip��:��(G�7�#X�5�`c����9��N���!0���H2�0P
?� �l�~&�`א�5EZ�o�7���?±c0����4�v���m�������$�]G��?��y�<ޮ�Ya��BW��_&QV��]�N��y Wנw
�Ƞ~�Y:������A�o���?�KI��������}����a�.��ڊ�a�[��6���o�����M�2`�>s�6��a�4D�����h/�b��<��G��f��9���3w1���<�M��U3���Ǝ%�7���N_���+�}w=����W� ��?G�B΍�$�,{b��3]E����-�(c?_��F����ܽi�^w�J�
��긜�&A+�ΐ�w��Y�,pg����w����X+�nu�]�w�����9m����QH�_	-v`���9G���V$@��Wzb�`�]� ��I?mH����-�&��A,;m��FP(�Ȫ ��x�RR�F�*�SY
^����[���u��G���A��S)X[�58��gౠ��績e�罞�(�6��X�O�.Fs!t�|�;e�ψR�{�P�KtO�0s>�����G�TP}���͈�*8�A^E����[�myՙY(���]�=�ELc�[��a4!m�0[�đ�=~ �,�;$�]�Ki-򛁡8b����{�Db�5~�����ulr�{������Sp&+/Ļ��yk9��!4�׆Ud�O���3�EK �$f��_���X1 �	%�U|��EW�%n�Q����V�Ҿ��.lA��I�Wi�~@�п0m�=�՚�5,qx��mB��@���!��խ-o1���V���N���7U��,ӊ4�ϴ#�A�&ϋ�r���9$����P�}�����Ft��m��?�Cƿt���@re1�Cd���G�U��r4ڷ��I�эl)/�\S�c�k�rSA���e�7�L�lr_��X��3oߥa�]-�����;�T��6}γ���}�{�d�^<����6��s�
:��#W��� �6��g?��O
m��}�/︴��β�%�[pY�x4�8u��.��]�\��Ah�ݤ�Ί�f��}��m��ֲ̀BNH^�$c���a_���>��/�߿�>�Al@��z�ޮ��z}'	 �9��?|��;�w>����~���؞Ǿ[׽�
K�i@͌�@��.��dfK$��� ��$�@��,7�N�����{�l[���� !�(F��v����h�c�����6A�v�~��o�O:|���	TA)�w�;��!@�����A#~]?�Aܫ�����;6����q8UoA�?ү���Sx�z��0y
�	�d��$I7�� �p.���%��0����Ɲ��~t~�8K�UX6
��u4�A���'�hC��_8ۜv�1���:g*�h���"��4���(�ZC�� ��hD�F�����#vt���eQ�$X�Mci?���BPj��y�{)w��h�3�4�B��B��^==�D�<����� Cx֊����V%ݱ�?dv��A��_��)��Q�]��b��2�b�00W�2�F]�Ξ{����6H�aYv�Zhz�`=k,x�Þ
�t|��C�P�)~/J�g��m�wM94\�G��4����e�>��#J�J)I�� ����p�#�<ks������O���A��n�����p=�(����8�������)��1�����冣�Zȋ��'��G�NF��\Uk_���g ��p�ή#ג	0rL�#�b9��b���x ��W�4�1��Xb�!�N=�3�̊;��tF�הo1_�IW���)3_�i8.8��,�J�>�z����`�O� ��!D�	u^���� |b����& ^�����ؐutR<O��<�z�4`����Uu������j!X5�se�t�G*�]�M�_�
����r޹N���{���I�2��I�L;OO~�Ơ�%�Pth8sL�|��tR�)u$�4ݲ�M�Q�$��&C�F����񆁯��B���g�?�~��j�v�T��w���Qw�TL�c�Vx/Yl\�W�!��;���	t��v�n��{�m���_��2�\H����@`�k+�"_�!t�{~�FR�8=�:��˦���d��	o�6�1�D#I Y��3P�����v�Ǹv
	�:��-���v�i>s�囑H��/�#�F$�����Jh*����9{<U���L�d9��g�$���(�9�p�:�y��^Lܮ�@źX[Un�t�}c�y�ݐ�z�)*��S�A7B'N�1b6���H]�8x*��fɓ9�a5�M�Q'Tp�"��7���\Xo��J�f�?�i��}�Ob%�dI}���ȫa")W��؉�8m-VP�s>b��q�le��%��2Nv��$h�Y���F�لNz�&�%��8H	�J�0�1};�A_y&}Y�l�v_��K���A�ʠF�ׄo�.x&qA����_�̢��
j��A���oج�ׄ�2������C�� {����E� 6K]��I��G�=�4@G�-�e�������#��Q��[7�\�)wLy'��p$�D�5L3J�cR^�q�Xb�k���N˦�i�Y��9P16m�=p��DG+O��8�d�^��ږMs�_"h�v��okdR5g��0.�m�ۤ �`��Q�:x얶?�!Y$�t K���P�yT��7���!���k«�O�П+�n�O�@tM��������ɰ-��1TN�
2v}n�޿���r��g\�S_��	�M¾QN�}�Dc$�O��Ĉ9K��G�G�SV4U������G�c;��o�D���}C����3��n�HzHL*ޭ���N�g���(m���C}x�t~��/��K3㮔���z�ޮo����/�������c�������_���p��恆M�3_��U���.T�@�� �3hi 	:7A��X��㖊��u�(e�\ O���%��Y8�a��<5��az���Ѱ�w
V�YǤc[��.��UA�Ne���� �AW���|v�#4�	3ܴ�x�a�$�r��1&�3s���w�#wr(���?s�u9��`�`i��u�~`�������& �4ϳ����1���� �G[�n�� lȶ��]��6c�g�����㌶[�V��Ęhr����^Q�h��ޔ>+F��.J�{`2�c��V��9:�z�Yy����Ėk��ڔ�
{+_�$|3�٘�j K�{� |D	2�w9C!�Ŏ+m���1��<���۳��<A���Ĺ�u���{���7��h|4F38R�x�`�A���C��弄�Jox�#�lg�r�_3G�D�b��p�k��o��I	z~{��8�:٣�����CX��w�5ji�Y��0�%����O�(;�� �ͶPΖ}���C��n�=���~��5=Y"����\e����m���X��3<��v�W���̓��;��[�\��;G��k([���f4�g�!yL�����6�@��!�[�_�������l:=�����H�I�#�7xv~�s�#����.�;&�',�S|х�q���N��1<\��c=�M9���Ñ��ι�`��a����Mur;պ��f���ђ#�IO�Ksq��K�-͝S�[J�*&�z�PO89u�
���� !�0����K7���orO�8�]q�R�K�>�hG<ȪIX�mU,hѷ!�t��-�����)$4m�.}��ܿ����Br���{.I}|�������l��yc������W,s�ץ�x'ާ�;�)hp����Ne��zߨ���xv�����K[k�Yׂ��uI�B��Vv\ך��������8B&���V5Кs]�k-��X�ޢ��F,���e:�[�e[��i��:EM��Hb���E7����dx`5�_��j#d�0�����E7?�_�u?~d޷�<�w���LZ����<�.?�2�
��F�xYkY&�e������$��`����_�#7�	��F��
�c��ne�3Ĩ��a��$!�3n�?�_��`�r�dNϵЬ���ّ\�* ���+��x5ȕ{� ��\`$Ȕ��쑌�Q��y�����#gTwkC��C���9<� sa�?Z���9��ɫLޝk��!��})-��lpM�����+AF����c�R�+�P�	�܄l:-"�]ez��&D���}(S�h���M��h�8u�̙�E$	��3�A����c�AA���4���i�I��.��;��.ky�g �b���^;y0�A��H�֭���R�y��լ�=�+���p��+>���u��������U��)���c$a;a�!G���볕���3���0���)e�e��1b�%.cO���H�
!K`�c���GK�t�g^͎O��tP0�+M*&�!'.z����9�D���k�i��+=68����~��=8��M�»{_�ǐ��f�?���#񚎆�"�4/��*���8��V��e��9�n"����li�۞����'��G<Sv(��S���|�i���~���7�������W�}��?�|��ު �]o�����?����Y�O?�������w���O��}���TzjO�~A��omܴ�G�L%J�h ��)N� � �n�P�ÈN�/iՀ�Rn���,=
��x��F�����}�-������[�)�e�����	\��S=��ʳ�w���%Ss^���޾��i�$��>� j��&+��z�����y�#��H ����U�܂�:�� ��#F�e��#�+A޶K|���^���x�W�a0���^fY;w� F����Ϋ=�u`=��%�A#��Y�f R2.�l�f��Y��Xr@k�����5���a4���B�#ۼ��|o҆3�N�|���v���:4Y;/�I
��!��%�ޝs}/�&մz��|��f�)�O�X�:v�����at���%����/8	�@ؖ$H��9]��aτ�q༙��!�޼��y���9�&]�c������8y^��Ŏ���Lϻ��u9�4�|��ޙ�`wa�9vȺ�5G��9�x�qj���,vR#��e��XV��I
ɏ.1�V��&�R�;�R�e4�ָ�(���]S�˿[Tux�����宣_k|G��j�K����>7����wY5��G���G:Y�j�sl�EH �����k�1�/�D����Y#+��(���l~n,t�eP%VKT��|d��R�3 �|.�y�z"�%d�`�bK���5i����|hV|K��I5F'�q��fm����9Wq�vqX8�������:�T����e%p�t�i!�z�6G��@�a����鍬h2�CuʑXPCb�F҉�KY�����L��N
�f��Cr��ш:�nȃq���m��3�4�����f��!;V1���I����26eU���ߘ����f�p�J�wop]��ss��v����H�ߵ��0B��s�b� ��� �5�C��d�n�;V6$P��g��f�je	j�/q��L�:�1��۽�)>H�$0���pD��師���$,�=j��߱=��BT(	]� 2���&!972�h�U�B/8��܂�G�j&��9��mB��/��8�M��g��̵]�����d!����Վ����?  .7[$?z�S����A�C~�y�)?:j�&��9}z�~�'O�9����4�zO�U_	��T�F�5��\�V���/f�>@�I�J���>/��Ʋ��8�.�XwO.�1�f`��H9�ep�B�yŧ�����5�Y�9��k2�u��C�����%���9I��8�f�.��	=�qǏy`�&��������pFҐf��rR�'��#�$��쪞�:�ف��I�g�=x�U1ސe��ر�m< #:����UB`��q^�_Ș��Z%B0���H��߶��MY�)<����R�F3�g8�,�s�㰁�L� 9�K�,���.�%�+[�g5�-kr�$�NW��<t���C�Z'&U<Z2q��扤�|M]ʣMoGU˭�G� �i���VU)�;�M�Y?��1'��J�j�{Α�=�˹$#�>��ir��I����2n��A��aMalX[��i�J���������1x>�j�In't�<4�F͇~6$��2���T��[-� �*z�.�	�ƕ*�7��c�ZtY��G57�ě� ?�?~��l~�~���1wҚ23�'~�ߧ��L{�����[
��3S*me׿�
�b�"��{��G��E�r��&05�vkSAM�)pZ�*:��C�g��.�ϴ�G 6����=��>�����������o~�[������ꫯ�A�����v�]o���]T h��'��������������О�8��1��g�c���P@�{�4���ST�鮀�[��	NR�!;��t���4jp�#9��t�Ip-Am��%Eh9:�C�SޘP���)��] 8�c��
�)�&{y�>a�	4��K���U�	H�ƨ����Ǐ��g��YG���fk�/����n	��je42��~iD1+~K �x=בـ�<9��$/�^�f�pc��50(�~kb�%)`�	O6�Y�2#��z��*/A[ǆ<�ѝ>xe�sHI^�q�wz���kN�ԓn����!��p4�O��ݹf�wT���^@ϴ���t!+���,Ku&��B�T� ��LJHN�܉d�d�{ḅQ�3��!��r���wNgL8f@����AW���EI\�+�%e
�N����M��85��06����%3�e�5���	�����{�yޏ$�'DG��p\1��f��9�͍l��L�N���b��򓉱pP����7�F��������?8�/'y��4�у���9X.ηt����2�(Iނ�g���F����(Z�u~���*>��0�N�#��G��n�]�R�b�?d��Ǔ'E�r��ϩ���m���xlvՃ�Q�8�D�������[�p�㡥��-v5��8j _V{��#d�N-����->�� =�ï\�L�s`��M����ӝ1j�z=��eM`/ٯ;.C1a)�X��KT`t&/�`�N$u�s�uc�k�0w���ğJ}`��<㹡�����T�M���Awa�;�tpi��Ay��;���\����I��Z�~݋]g�A�ٔ\}˞P7�4J�^���S$���X�9�9Oz��SBSgrV������#�3���ּ)ִl_���,tiN*�{����[��=�/�8R�#�su�՚�{���g:a�ZH@[mu�V��&ɹ�7'!e�f�Z�%/M.ȑ�&���%���~iߠ嗛JTN��mb�K��L,�ʫ��|��M~Ȝ���n���U'��	�,S'R��F+�J�0$.��Tl��1�Yv+FE�y7ys0,m8GvL�v����1���l�+�D�Q&#v}�˟Ag�70��gf�R(}�5j9��1�:]֋�,1������L����ZCx
,gEw���|�6��������k"�ZƂ�T�������J_w���q�����ة�PO,��0�hwPvh2�ӛ6[��l|?��K~�Q�f]CC�<����?*/�;�|2q����;��� O@���
����):]����^p�����0�"u��B��jA[T�Z]F�䜞H�k�F�cF|N�Ό;�E��|�RV@�ǩ��/Z�� #��&���:@Y�wzڙ�HލU)�ǒ���K��΃/)�xS��: 	�g����E��S9Ǡk/&6�W�Y.c�zp\Vc�g�����{V�KY�4 ��#xX�`��P��0���P��"���;{�I�Fz7�>�=��l����'��RT����A�,�w[��1�G�_oHB�t�=���R�^a�H��悯�A���!'¦�������� ��c➮|��	��dFM��4鴵WkZ)�K���*�`{x2"b?�60��k	v������_lچ��pɢ�4�B��3_U ���V����J��]������h<�ſ�����ܿ��C9b����z�}��-E�G���7�T���7ďTH~z袎Dnc� ׇ���e�߁FS7�8<�{��b���/�������������������/�������{�ޮ������;I ���>{���G{�#/��p�+f:�A����e�����@C��W�CT5�����C	g�%���y��w�1hcܨ9{,=� pP+%TM��$�サ�^緛�:�^��	�淶������Q�:��o��ƾ���e&�峆e%a`]z�A�Q�y�t�gUk�W�t�ȈD[���AC*���bp���!�x���0�����[�/vB$�G��U��Z;H��ع��>�wx&P
-Ki8Y���0$� E��٩f��/��WjgiP�t�|7���nt���v�yw[��FF�����ݭ,�Qv�ѐcD� ;��N@	*�9c9�Xˠ��։v
�M���RI$Vx9x���s<!� o����.|��o7�Zd�x��{�k����t�
����y�ri��b�u��:r e?�0�k9\�缻<Y�w kY� �n�s�����<�gJwa�N)��&���R��0�0��G���3`k��#J	x;���:�9h�x%��8o0��c���~������Zo=�x>�I�k�w�xU�s���u��|��H�*���r$@w�9�>�H%��q����|���#J�8�bR ;P%`��9M�^޳�J��m�)�V��؅����;8,`�w k�h��5��`���ȹj����ހ��'ۦGP���E���X�'=�L��hЃ��	cA���Cp�Z���_xH;��yrg͑kwt���l�Sc`g�F���H����YE!�f�Ɲ�Gv� y"���n����{�DvqF2��I�6<� ����r��9�nHl`E��8ֳt ��o<�+��a���W��S�D@���C���*b�Ջi�6�C�c�9��~��c�<��g��ξ!0�8�@<�C�[�%H��K3��B^���]���	����S����½N8��`:qә�ʕĒ�,��t:��ϳơ��d�=���/;�������г�4�Cl�|W�H��/���6���1(��5 B����<�~��5��1`"����>����g���}f���`̪f�����Cz�:�ҝ��I��$)��P��l҆$Zs	x)��.���F�:W�o��Z;�s3����yq�g�w��y�ȇ�;�n C"�<�_�]������$���޵��F0	�OV�!��`�Z�GMb1��!;�8��.�����c$=ב+aہ�\�-Pxz��g��zm=�4rEb�H���3����o�/D�$.�q$�������� /b~Bv"������6����Ǔ��k�9&��'l�0ϣ[F��ӱ� ЇeR)�W����J��L�kHJ|�"��#u�"́�L�G�ƅ>�h�(k��>���:8�
���G�3!+-��^�MlN�yRf��хo�sVQ�)gC����fVe���;�;g�=�E��8�G�<��?�ލ��2��<� u�u�C9⨒���?%�9���\'��q�VB3��9+�'6;ţ�{y=j-�-�$�r��c8�2��F���["�i&,�֚'	^�J�V��]◃�<�g)8h_Ki��^���,y�cG�6�+�4���	Ƶ�?�!�g��`/yw��4�v�C�.l.r���Z��h�L�?m�\���&?�ȼ�����r��}z'�9b�c>��U �G����GT?��?���5��$jEf ×�0�x�DP_�N���2<�����|c����>$�,������*���Q�e Z*��x�Xȭ�����U��Aܴ��z}j7���"S.L�������?��].Ϻ~��Ĥ �&�]�`���������w.}P�k�� ����=�����L��R_���Ѫ}�7�|�9lD�e�����u���~%�~w��L<_��m{��"u8���/m?���������}�����g�ԟ���&y�ޮ�����]$ X����wO��w{�i����v�DP�@� �%�]�>,��V�=-�
"�5�@6�iW��w$dl-�����fyt�nK�.��#��BM��A��-��R���9�P��	,Jo�v����Q^�mmz��ñց�К��~����W_}e��{bI�4�`x�^��pF<�斷Ae� @���t*X�/��[7��{ @A�J��E�-��Ȣ�����|�.����m�����>7�{��2��Ԭ�u_����Z�3
Ah��@���ݐ��x�a|��z���'�`�(s-s`y�|���bzZ�2���3��#i���:��&x2x�r����eհ��;j@z��A�u����p�.E���+Ȕ/��p�4�w�g��|��bnD+8�}[�� ,�,�2�nO�������X��v+����ɧ�F��b�G�e�R���8����V��_A�I��A��J�VP2x��d)Q�9h,��U��g���G�h���s���R����oa��A%: w�g9����D�у�G�n�o�e��FQ?�x�^"�aw���ؐ�0�)���p
�8�!e<yg~�G�шH�6��uy�� ,|�s�� ��#;�W�v/������m�x�?~2�ٕO��4qf�w���n����qY�~ș���4˥䭳�y����Fi�
�uz�������%w�Ļ�G�"�G��#��-�K��LJ�����K|����>p�R�/��p�t:�CE�U�,�ę	g${X��	1&��u9'�9�ɛ�]N�mg��_��rc���О�������en�;�@��#��s/:xN�{!C�w��Ym#���� ��p2b�?0Y��v�$;RR��"X���٧Y�7^�:+���>�s��q�@u���N�1V0!�F�}�|k��U�#x� 0�w�P�9�����\�"�#mO��d�3�OKlG�k�m�UpT��D�1��ȷ��1���y�����,�>gb�NV��2gy�X#	���5'�(b�DI��O�k�?8���p��G�dD��]��L��Bl �{��U1��^�y�oZl������s��P�4J��q���xc3&�x{������@�D]7��|��Sb�K0��U�B��o�28:4�Y9��F�L|C����?b�ֽ�,���	�)�7f[Ϟ�e�͘Tۂ�.�8n�~�R�J]jb����y���;h(v�:� �L�$.�&��8��{��xUr$F֤�%ΊmL8��?���&բR�'��\G���kd �y?���:��N��K$Ԟ.�Sf�s�!�Z��%�c#�	Jœ��2&:ju�30RM�m+A eW�1��2����:�8*ǹп"G2AZ�u���Vc��y�z��e�s���ɣ���:�络;"���¶Xu-l�şk�EUMT'X��t��5=��nlA+���~H|N/zU��SC"��[_�0�B���WW�cK��:80��%����W4jwҸ�4�"�@#����n�`/�\;2�8�z�p���u�=�Ab��+���ܲ�i�K_2�g�;��38��	X�hc=������{��C|[�Gb���s�>bA�E:�'��L�oYEe�d�6V9����$2l�<m�_`�z��_t����l��J6Gʈ�p�Kr����mX/����k�ŹkX�}���c#xn�#�<y)4��Pl�_r=�y#�Ys��b�����B�/��9VbKܔ���Oc�MAH�ˣ�|б����N���<���+�g�՛�?��<�qHu�E�#�u�Z� X9���Ǘk�3G{2Z��Z��1���3��2�O�>��_���?��� ��&}���EpT�e��;ŚC��U�T��1�&�IO{_�w��O\k��n���=�����5ig��U����8��fk!�@����B��� �Ү%-2!}ә������������Ӈ2|��Y������/8ػ���z�ޮׯ�$�w?�?��o|�������'ہM�����48���Y��	P1��t}<�΂������Z�ڳ#���
ÝA �8�X������@۩B�Ӑf��{�l�q8x��\��J3#0ԁ:�2 ;�,���z@���4ϐ� P�W/1��m��P񫺷WxyS�>|�������_G��ǚo�Z�s���~�;�����%#;w:�����Ý�<��@�t�����<�ґt�`��`�?�~��8�d�wD�Ov�!��c
��(=���s��s�����go�`��-@X�x���]�˼aM���A�wI1�o���A��[��|q��"���VPw��!��)(�]��E�h�1��9u<�9�=Bs}�k9��S�=�i{��#�̣W��g�ҡRǁq��?�x�Y����o:�I��f�<{���o�޿@�J�畔����N����}���7K�F��
.��y��&ߪ�
���c�[C�ä���}mb��,�18���7����R�b�����8V���ppB��~��!�K�W^�}-߁��~���9Z&���|	�0�9��G��	]W�E�����O�w��Uy��B���r�&O�c��E����Ȅs^��t,��*�P��[;�Zˑ%�-�k늉N�k�N�^��H�5���d�Yɗ$&�*��|�!Q�0蓻e����T�q �>>���4��5~��Sc�/�o�p(�tT{h�C��i�sс=v�K�B�G�N��N���Q�Jg�E��7r�ř���z���S��>�LL���%�A��w�;۫��D�{�HT�S�Yuͼ�Y���Ƚ���?�_��!�K�D�W>�u#�U���i�ӄsńY&��8$��1{���޳��6��OǢ�y��)Z�޳�B�k��^Ǩk��a�mnsa�B?��F[Iu�l����ʿj����Z�馻�Z�΃�@�Փ5m�G�	���gd[��t�v�:��w���*6��0m�A�ԮX�����`G�Q`���0mE��;�S��V�Jh�%5���^Х⺤l����3�3x2"�r#�nlP[z�8i���%��2���R=&�λ>l٥�jw��@�4�mوN�*��M���ݶG��b�k����Ȁ�.FȄN�y_V��
	t��M����@i�7a�X�;ܖY���f3�Ӽ���Q״�%�q�U��v�Gi^��U�(^�=�o�/w~�;�::w��w*��?���;^���H��Ϲ�\Y���vm����DJ�]���us	��8�?�<�ͼԎ�ul����;�fws�r�"���T��>�~�M����9bҎ�s\�:r�G��χ#fY�k�O��8B7����і���r��>�������#lx�:�NO^�>(��#Ǿ���m[�/�V��r��5"aG�E��&��.m���[�!���Zn�6ᣘ��������c�	PQƕ�`���ع�T�5᭜����ݴ��>i�Dg�S۰�ye)�fj��^�Ǫ�U��}�:������/k�iV�|�^<�O�IT~���d0ǖ}�u�U�&�*q-��=����.w����.׮4&M)�0G[�*�B"&�����q��s~��_���g�����3�O�Q�����z�ޮ��H ����o���/�����������������"���ܱ4��P* ���%�N�
v	x�6F�bF[G���x��Px����ܩ3D) C�EҀ`��(���Ѹ{3��{��Y�el��ũ��7�~7H�ÿ�Ҿh��N�9���7V"����6�^y��f�2��]��� ��i�xԄ�:�M� L�cw�Ɖ�g�KW�ȀI΀�M���F���l��f�F�t��q���b�~�m3��Ns�� �gx��<��r�a�Z[������fh�9�	���U�8�G����ɼ�H#��8���؎"�&/Z�ؾYp�\о�m��k�8��F� ���N��~��U�������ſ����#�:R�h�&�I
Ggv�=߲����������/�O��0��dz�@O�!���Y�>���]I�A������#P��,�k��I�ZwK���ΐž������q�}h?�q9<���"dt-v�#[�Uc4,�V�ب�ʲ��ߕ?Q��}տ��A�#p΀>�Υ�Z3&�AG6���6i�����k3w�����v\N�X���?t�ӕ�q����S�X�tL�'�Lޓ��1��8��Py�:-�Pi�;���I`��*:�.|0.�ތm�}dBK�Y��3C�$Z�d!Uոli�������IE�qY�9�-�V3A�'�w���\��aY�6��AG��4�w�=�$��ۄ��\x�2�e�I���m!'b5A+ݖ�'�w���J�.���D����+c��c-�P-YqQ�1�;�!X}Y|�Ir���ًmn�<A��S{���0���>kU(M�{}�� �ё6V123Ib��d�^k�w��y!h��a�ー��~$)I�8A�a,-l��&�w�*�����s�i,��b���IP&yj�Zѡ��M
��~q>�Ws��ri�a�OXǻ]�+�>��Y��K퟽&�\{���ϋG��������~:�3i븾��mA�@�d%�=�	n������v`b�7�|�vU���f�K��Udd��`r]���C�r}`Q�1}nd���{ʴ�4�f�[@S̗����n�O��j 
�#����d_��?�8�_��󻶨�fJ{e�.r�X��l�� ՝��k����@q�m#���pW�;���H��t�E`cA韖���u=^zL���֯Wj�����<����-ɫ�X0~MJp;Q���*�)WG��J��_~G�v]�9+��Vt*����ؾ�{`�1��rI�ܱ�$������Kk�&ڪ(��3핪ӯ��	6Ab!d��u�g��W7<?�[���'߬�yɗi�:�-��A����t�r�Us���}�ƹL�&�S�Vx���Q���Ϩ7䥕B���뚕�,P����aFY��e��s��اɤm��m�(�0��JC�e��{��ے�E�o�s�}գ����V7.K�@�	B�G�XX������	&�yH0 0�-� 	1�	0�����v��2�]�]�y���J������"2׷o5ԝ��ꞽ�Z�2####~��Ndcq�/d4�m��
Oc��q�t�}`^ȼ����|6�m���{䇮�lx��ۛ�����g���������߯o��������^�2�T �u=���������_����_�������/.��w�[��Z�<0���e�Q� ��G�
�W���0�Y���m�4��ǄAc�AW�p�j~o�V�a5���ˀ?�o�O�úR6�<!E�o�]8t�g��S���43Rq6��ڋ2 �FӮ��`�����$���.h�`�P,-�*O�:g�GK����^8��މ�NWv
w\�ZI�J�=$�X�Uc%� �e�K��0����6�`]s��nP�1�� u���?w t��h������Toepp �S;����<qRf>N����C�:;�#_`����sҟUN�u���/N��܈�Q;x]�}��⎇����G&cs��%-�ߟ�{�o���͸#��}�;�+���<�1rD>T��������9m���U�KO�t��怃������Q���.��w���r`�k�%��3�cm�	��Xǧ��m��ףY�G��3u�*���e'kL$<�|�]T��e���H��U�$I�)%f*�'�1~�h�>�!�l��a�p
����҃��7;��c'�F�^���]N��e���cgi��� �Uk��<���m���W�! �o�,��<̂�=�Om��� `L�	(t}�������ס�P�=����%���.LR�]�~��sQ�O� �vAe�*Zو8VH�9ŭu�+���"VK]Ɏ�v. %��m셔����ulc��*?��$h�
 �"��k���R�D���zz�ҮD��~]&GG{�/O\��Y.��Wx����L�)?���I���S�u �	Bx0E�s�cE���,?%��v�,�`�$��*3n�
w�M�+6\�B�5��u�t�kZ����ŏ��ڿ^���>�h�t4-c*N�P'�~��0��>�d������u)Ǝ�U�(�ǘ*�϶�<��y�/|�.!]�*&��Bb_� ��Ed}r�z����MD)�S�z�TavU���np����v�/�s�w�~�q4|#�>�cmm�;9ݞ���^��y;�rM' �v���q�'��l��[`��O����e\c��������A��[�[�[M���� /G���N�����|����?�\��ǘs�Ͷ�
����]�&=-e��^f[��;�K�� �n+�߿�"*N�-T�u+�F܋­�������V�� �g�iaR����>�eR�������-aT����0��O�M�<�Z�%�>���r�U�!_�!��E��/	wT��֜��4��Lڊ���긬��&��S���հ�'��w��$�����m��L��y�C�k�G�	��*�!;��T��<8�1,1,����Z�q>K��`r��S�Ɍ�B�4��<A�OQ��L��~,8�	pnE����5]/7j�.5������Xn��ktY�?�q ��[\ԅ�V�3��2t��y��
����o6�7�]n���t��Ҥ"�{��3K���^?~`���w����'����W۫O����ց����^�K���� ��w_���O�c�w����������w۵P)�� aR\-�G��j���qҒ�\���U��c�ܡ�7w&{q��i��}8;��:�W�}U���`�[����ջ]���:��'�XL�̪�~g8i��������ӭ�ek�A�8n�T �ϰ^����}7�(&ȷ���`C<�]x>�5�>��ǛL1H��W�n�F��A�-��΋�l�A>�UO�оTG
m�B%YW�VN����v�^#ʆ�O�i���Ղ��ns��D����(��<��19��΀�}�գ���ǚO,�*X�j3O�8G�;'+��h�r>;z� ʺ⾵��ƚL�;7d�A�VY�<����2��T3tǯܕW��T_:��R׹s	��+�����B��u\�������C������8iǴ��6��<Y��u��o�d��A�ˆwm�C*�HgԇhK�u_Tŵ�;
'el_�S:�,v�Gu��M�,����`9��c
A��}Y�/ǜC�}�k�l`�m�B�Qv=#�o&�nL��!�Lj9��D�d�+d�Ns�XqzQ7h۶8F�A�*�[��`,�o�]Uy���y�#hl���	��V6��_5,�lﯸg=۟~�N0N�,�D��=���,�Os{�'���!�h����j��h��]MH�5Rs���z����}��N
:zM3��f����?��W��C��RS[dR95�40��}�g�����1^��Oh,mU�i��n?X�4F�H�<e���O�u�H����&���+�$�XYv.a�5��m���|R���/���3Ҹ�	�=�\p��B9Ԗ0\Me��A����.�����i�#i_�Iذ�y����ޢ�#ݲ�W��oɿт]x�.�f��W궒m�z��w�^�ﱍ�vu���r��Yz�{��%�d�/�0�ڔ��M�tB�k�H�ac��&W4�<�x�u��nY�!�����<�M�_����`��na��N+>9t�>��h�c��O[\�Qn���U�?�.(������Q�V��y�P,ϒ�[���o�u���2�l��T�~����q w!'=PJ��D~�P�x� Y�偧�A%���o091,���ܢ>�/]��֓Y�w�x-�g^�F�:V���߯g'�D�Bl�:;������_dH��M���Q����>�_0V��,��HO�u�n\��i��:�Q�����N��mХ]�7*�~�����[�g�{�ˬ�c���uĸ�����-��CO�)[�t�E�ǯ���5w��aO�Y�����8dg)N�J�o�l�ߺ��.'���$�E@X�n!f�Ӧ'���0��Xz<��]�L�M���}���EY��d_���O�֒Ǫ�ׁ��w�O����;�۰����Um� NS=��e�C~�k�
�ө�G�/Ƹ�#�7����5�o?A`�D������ꎛι�����~������_���|I/�%����u, ���3O���߿��G�_�|���z��~��ށ��Մ #AO����Z����B�Ԇ���v�b(һ��$��ʣ�a�Z���;x�jw э�0s�>&�{��D9�`�'֫�1� @��lЀG�����r�N㾚�����P�^���d�� �7��i�-s���>�yv�Es�վ�b�VZ� �t\{�uɓH��r�e������t�s��).Wd��o3M��'u <��V�]T���KG?l�z���"�V׿ؿy��h�m-���xf�0Cq:'7��&�r�D��>"�Y�A;�%ugSN�(��־Q���5O	�P^!��Y�e唠���3�F�Cc,�`�]�d@~���W�ds�s��g�O+>���:�<��x��7[�����W��.�D��Z���Lt�Y��O�M�6��r-��W{�x0��LW|�}��ӿ��~+�8�G��ۏr4p�|ߣ���)�;@��Eڅ{
����h#��Ƈ:�(�v-��L�d�?�N��z��m3oW�)�@)���Z����iZ����l|��}
Nl_(#=��+VQ۫�LW��>��@>��bz�i�]��n��(Wu\�Y����[�c�'xmR~���+w1j�z��vq��;������(�M��c�D�hψRi���a��2H�}�'z7qϛ�3�L���M1(���c���]�`��!C��}ha�Bc�/��i<E��^��q��P����8��\�ie�@�6=�q�ϴΨp�;�'�W4�h��U�HKu.�òeO4Q>���X?��W�r?EܙqK�_�i���m��lc��;�)��i��gnhy�Ye]<�q��+=9�:�H=5з��T��A��f�`Y:�V>�/����q�4���`�2�'�4���^���28� YϾZ�\��~l�������f9U���'�D���=ۈ+��W9����S�E�Fڈӄ��4�O�h�O鷼imݠ����쵬�����~�l�U���Կc>�u�J�f{5�)ҷ*����r�(��q��$Kk�=j��B�x�-����������g��"�@��ゑi�QmzÂ(#�����nbWl�=N�j^��W�0�f���)��l9�,c�U����\cy,�ƪ�f��x��qs�c�f*���
[�6���N�I���"�S,׾�HڎȦ�-���jM��[Lu<��g�I�0naN-k����lІ�X,�/�,���X�"��4�p�ͣ~B@���-�4�q��rj�W,~<��ڮ��Ѯc��u�ꛇ��O�ǷW�<<<���+^�KzI/iJ_���?���g�����ۿ�7����.�`��#��Q:tVpkС����V0�&fz�a,����t6+���#?;Qu|[������m!��b-i������+J������sq"��_�^�C��h7�������{p��NV�Y���
p����V��rs�ѯ��+0��\�>�;�ˊ't$v9��Hˎ@N�Gs��c~�e��[�� �VgW��C��,�4���ʢ�G��9������Q���?��7O������O}�1i��t��Jv6V}��k��v�b���<�1�jz�Fp|�8�]�nP�I��(�o�JU�z&���0u|W�d�3��j�ىU=����<T��$��'�V�Y�p�?�Q;_��T��C^�:ؕS8!fMSlלw�W��j��q�<����R��.Ҽ�|s;s�.�xX��,G���~�$�c�6���5�A�����ℏ��n`�#�Y�Sy�|k��D�C�+k��`�<���s�;�|V�����i����f�w�	�����6cM�l7u<����XP��'����)���}��,������Y��+g|�<�M�Ϟ'�Ş�M�����?U'e���R��:q.���d����m�,3���*�-�
��+�#���)�l�J��d��T�᯼�2ʲI_�~�'�h#V|N����{_u��(�/f���X�Y���'k�r��]���(m�!\�"N�k汒�raͬO4����t~~O�V�As+��up�4i����?�m��L2"-�;��_�-@d�3N�)iG�W�ͧb�]�S�+;����N��1�v����2��U7��f���Ӛ'D5�}H�g���<�&��9�8�Q�~�s�~��bo�N_[z>��qL0��v�/��T��U=x+�W�W.;���B��y��E"�\�?�s���$�]E�33��b�I�p���-�}�����Ϊ|`���u��^��_f����?���e�aU'�PC�k襼0���x2��nM���Sy�D1VY�G}��{nHƕ+�������E�Ŷ�|��
��}��Iz���W��յ�?��(�{x9^�f�L������ZOf@e=�7�s��µ��DR,̫<�т<�����,O�3�t�Ϻz�3��+}����~�����Y���{��?���������ի���^�KzI/��ײ ����կ��������s?w���_l�=ܔ[��]њ����
�Y��0����P�]��'E����C4΄����GVo�`}q@s�Z12������>� Ս꠷b��ܦP?V<G�G�?_є�*�M�\w@��9X�Oxx����|�J+��n�z �@w�K7���KKN]v^s[��N2��i�6��A������Ύ�[յr�	2�ߢ^�}֮{�}�����x��?יv�����\v.'O�� ~Z���9��v�u7ê,�QVrʲ�$�~}��W��r��������=O�d�LߐvuT�0V�Dx_�N[����u}L����f�"���}�^�Q����ˊN`vX(�����؆�d%����Q���������w����n���ƀ�6gݤ�g�cj�sNYg��ydw��+V� �!�C����2�4)Sdr`b��/��U�σ����9`fۮϣ��X�N�9�/Ǣ��7X�6=_��2w����r�m��1��Ǖ��s�9X�IC��9 ?��HW��l�Yp0��=~�	�V�+���}l��_���P��m_7,'ʟ��l��~��c:����XWۘˌ�.C÷g�p5�2����X�h�m�b��O2��̷��U�j�.��v�l�<����8�f�Gq���G�$�G�$�5�Vw��+��}��u��X2�ֿɸ�L'���~R[�� �_�K�8}?Iʺxe3�_������<� ��~Ć3fX�vN�ޟ�a?������<J��]��l��iY��yYS�Yۃ�4�����z�'o�����}��+�C}��)�]\�������k���D~�~u:�_�Cޟ��^|L�׳��y��=Y��pD��x<ӣ��vo�3�Yy���#�MiXŮ4�����]�ǎE�y'�5�7�q�y�}E}��,e�ݫ����5mu�{�'3}��q�t\O�݊�<�����_�wRR�<����.(ߥ�@��������������]�1SX>�#�<�Z�9�~���~o4��Ed�8ƽ���mf9��0m���ż����*;�)�<�cc�;�������G�ƿ��~����Wfʤ���^�KZ�����#K�o�������������|���7n��fd��@����[M�;x����xl��lm�}\.�	7���� �o,hu@����FC����VƑsN`m�$�p�B� �VO�A^v*�~>�3Ǩ��k�%�i��D�q�8�n6��@]�;|�x>O����������ғ��B��ɑ>k���s@���]�v=;�\u��l�7s�3����Ε�)X׉��)'�;�Xu�Q/���"����VbPUc��klC���1c�]r� h[�7��o��I���u�s�Zw����g��n9��UP.ց�+��U�Aa�I�Ԁ+�]�3���3]�{Q�ɓ�B�w���q/�N>F΂x���C�1����iX�(�Y;9�r�UY9p����օ3�W��3���G]�i��&�|�m�.�'m+�]C(ߩL��U^EH�1��x�?�I�nw�
��t�1v%���ۢ�S���������;��9R����h�����2Ǌg�a]�� �@�U���Y��W��O#c�}������*�u��9����>ĉ�\����*���:c���f�gQW��|���s^�����m:v�A�y�I��)�=1�竅��pp�;�w�Gy��e�����Y�>0{϶_���h?��3^���(}g���wn�`��D�������y�'y2*�=�uS&�Xk}�2���Z6�wN߷/Z.���<�a�p��U�AK��U�F޾S"�����e7��@�d�U���Ť8d��8eGiZ/���lki���Z\P����R�֨O�R3'�u~η�5x��'M:�o��4c������uݤa���}�l����_�v*-�:�t�ڦՓ|_'��8��Oe�lB�෕�w�y<e}���4�u<`��{v0�X�Gg4!/��������rm����;�W~���wQ/So�O{x��aIe�r�����oc�q[�mc�ٗ�g�U6S2����A����-���ާ_B[�^���K���1�e(c�,�(;ei�ϑV��z�s��^��t�J��X���nY^�z%�����U��+�V�A� �?a�e3bȕ~��a�Az?Xur���q��+�/=ְ-�N�z{p�fE)�$����*��u��� �D8�	��~Θ�[��prh�����K����������?���������ƿ�����|ｏ>����U�/�%�����}@�]���������-����w��GO7��x�HJ�;v�ǝ+���8��{�tg����#��b*���t�7{r�3n�?�I�Ӷ�q_w�ƨ�"G����s���vI��ժ�R��+w��ǻ��}7΄���AI,/N�j>�Ƴ���0�o޼i+�![��l�y��W ����(���I������|����U���y��P�G�e�\h�
��^���݆�e�Q�P�����t�9������5���Ϳ*_d���U�e�۵s�N�S1Ͻv�����]�ܟ�+���dd�6�,���9��i��d~С�3�Q�Z{���/��[��e҇y�Sԛl���;��ݭG¦o0t�4��lϓ8�|v�-%#�M,Y�QF7@:р�ͅǗ�[�;i�[d!@���G%?��δ@W�Az�B�;~G�< r�%�Ù��+��98˝�8����,���>�1�<���־����,0Ez�p�j�;L��R�/�Q8���rl e[��QЏ-(e�{
�u$�<��d���������Yɢ��Y�}ƾ�[>G�e���{vF�[�N���yer��ꀬ[���+������B�q���U�l��3<��� '*���*`��E��U�l����J�xV���M�1�z���oy�uj>-/�E�gۧ���ċ��ɞky��g�d	��+��FvG~���=,��u �P����|����82�]��Vu��j<���������4h ��:��s{b��=�Q��$���z��Vs���T9�����6>�&�F�g����'�<[ɏʗҜ�pH֥J���,7+H�k��J����G��6���{������c�����l��}�ԥ��2��D�#c=�m�{�c���g>�q���#x�S[�}���p�-��3�GZWx'���8��\�7��x̾'yIKă�M��><�S\o��t���`�{�x%�9f����z���11�H�m�=�i��mѱ���W��>���P@�h^�a�4a�(�z$d�<������h*�ʈ���28���[��v�؝'�)��t�sz�W�/b^��$V���P�/�\�x�;v� ��2]q�v/�#�V}N��*i(�I N�>ҏ>X�/��C{�d�2�5��}�OP�[�xR�'��=r@��(�Ǹ���coЎ�^}�^v�1	#>���,zlse��V�{[l|�<=\>|���w���O>��7޻}𩽤���^ҝ�u\P���e�|�xSv��zپ�ޕ��B���y�-(|W�E*���qe|v��n@�ZX�^Xi
v��w}\����~Lm�C�=�����M)�0bB��VqLKs����~�k��ډ���[{w��i�4�8���?�3Xܲ�»��U�'���m����Ve�S�D�ݶ\�z�hOO���Ͽ�t�����}`
���%!�:����dF��S��J��Dpg.�(uu�x�*�����e+�}���w���FO��S��u^��81�m�򶿋����o3���vG������lNT��&����'�1Ȕy9/@Q`���q�J������q yJ���Hy��V3X��y�I>c@��g�3�!�k���B�@I��Dj��Zu1jt:r:,�g��G:6Uv��:.���)E΂J�/�8�A���	�E������OL4��Q��j��o�d)��4�ȊYo����A:�Jmu��wAwAR;m��S�U}�q >i��u�����jq�W��Rv�@O�R���CǏ���gB?��Gy���g��)����p_A��[X4��8�E��<�z�*��0��O�;����Z�؅lˏ��(WW��c0U����y�Q7�YۙLIk��qAm��Bݡ�����􋁲h�'��6h�]Lec�X'�R&>�uj{ZI� �3.2c cRm�PQb��|:��E
:N#�4S��>�Y�Ǽ3o����b�N�,�O��x;i��~��������2tn�*9е�S�6��2�D��a�h�>�̳��m�y��,X��G�=c��>w;����Y�ċ��2��G;M<�f{����\v��Ǆ����&��SҴ/m���j�EY�.�wJ�j��y�È�_5�g�hAq]�+��.� -&��ƒ��&nrjS|�v��N�~[��5m䭖�em�r {��Y_f�O.�G"�BQ2��Ͷ�E(�ި�㷚�W�q���M&�>�c6�h����v�M������W#m<����7y��ƿ��+����}��D_�w�M\%��)(]y��8'D�XѬ+���E;6�RXWƵ��ɣ�͘�y�����Dlu��_�e����o6���c�X�9���C���ijK��v}��u�.�Uʲ��oS�\���'����^�N��y�)��e����׫���1�����!�P,��;��n7��?�ɝ��x��4\8}�cȏ�;�0�8����iꢍ�U_Z���qv�u��)(��/�͈���Q��|�%s{FmRvwG��E -��I^Q[��d�6���y�=QVt��jk>3�1���������8�_�G:�ܡKʠ���a�Z=�]d�r��<�!Km���Ls4k��x���X�K�e[�y���G�g��o��������Fõ���#Ns}���h���|�����R����"��^�KzI��� V�JyS.�ᦻ��{��]��dw�C(�@��2~��Tjc���I�cŔ>����r1z��kk˨�0���vE�J�n?!	�h�[[�^��<�^�ɲ�U��]5O�i�@qe�S���lK����*_��rgp��5��t�O#�� +OOW{��];�4�I����.LP'��ݙ����\��v% ���ɫ��K�nz�~^5j ЉAE�����k���:�ϵ�	�GA�k�,�S�2�h.'?�n�%ɧ4��U�9�&�V�A�؞#(��p��h'�c�g�GZ��e�ަg��p�g������f����y��·�8��<����Ǹ�'t0?�͓-��� ��߳��<I�ay��� ��F����v����e��?/���L��ޏe�#�9��:t�C�<�����e��ErZh�nJ�/U��j�t�@&�ͶiFy³|���� ���[y|��8Vc�w����i�֍��1к�� i�5�G���H\�(���D[89��R��s ��j�����i�m=�<�Kې'�r�f�5��֔&�M'����nu��Jo1\q�r���>�X1������u_�Y2O"��9�)��B�r�Y�x��������1��;l�0���޻{�h~��<�Ѿ��|�4>;�]�_NX]`�ef�=�W��h�7��8{��y�z1�FZcX[�i�	v�[�}�D'��y�^����*��������������/�b�sO|�.���f��g��ZuiY[8���<���<�侩����J����/Vz\�|#��<3�v<����g|4�g��C��ZN$��?oH�"�=R��y{���g�hRH����Kɧ�Uǝ�9����hG�����<���K���z�L�~��(+�i_���r�G\8_6��פ=O�*d�d\�q�J�ۄ�շ�m�o�y��������o��ct�;��4����\���(�C�j���u�o�%�E���N�W�OcQnu���ϐS�5�u�lÅr)�ֽ.��<���W���5��V�M��T!� ���p���xR��������a�=������8N����Ò1�2s𯒠WV1�U��v#��=v����{'dE-E&L�u�Wg�R���]!��[�2~�_��t���v���A7��2
Wݢ�m�4KI��{����V���jm3K��ذ��}�G�/��n�Qڏk�Ecb}!��������l�+̾xW�򸽽Q��񃋽�ō�7_M(_�KzI��M?� ������������������/?���C�r�o��j��߆�걩�W�Su���"���&*{�<`�v���*�AO6R�u;�<�����Z[F^w��Lw~\�8ҥ������Ѳ��Q�Da%H.�MNC��k��9U��{��H#:��>>>�|`����}������l�f*��v�':W��� &|��ߚ"��R�U~��(w¬KÙ�"�yp ��~�@���+�A��B��|yL,g���_��^0��D�w>�_;�𷗓�VC]N�7u�5��m���,<ˀ�^��~Z�uI�������(��w�o���ު�g�bm��|Tۦ+�S���e*�\�ܾ�\���Ĉ������W����x٢����%�-W9g[�˭��=;%&cm���\/(�Vm�_x�J��5�����Υq�n��$��NU8wٔ���|�wI�7�ת�;[E�{���������7�/}\�ʺ��sy�$�~�+dl	A�Ǩ;\4yΑ���m-V��NǼȫ��������J��b3g��5������۹�W}�w2i *�	���c=�]b�ħf��&v�˳��ҷ��ܖ��6�[/���D�<��~C7��!k���V���I�N�+!�36Y�m��xw��C���N��i�����⍌;Vu����&��G��W|��y�j�|��2�Zǂ��0�'�A�چ��I{7U�W���Y�5���|�Gd���Г�沨_j����=>�\�z C'�/f��y	�)��S�j��Yһp�n��cq��h;8�|��K�Uj�;=�?�A��9^q����`N�X�9���j���#W�ul�k�o�z}�]���N.jP�b������e��8R�ؓc�|��3��ֶ~u�w�K�G�B^�#��6i8�i��k�4�9Ԇ&\��)K�F���ᯍI�W�ʾ��ڜh�&�χ&�����W��R��|�I��8m�ض-��`��70���йj���a�-���b�T���m��)����	}��e|/�\��'��WRo�Y�8?U7���Y�k�����b�;}�t��_a>��b2�%g�c�צ��8&���}GQ��+��u���|�l�v������1��.��V�8i�۵�OV��ux\|���7�[,��h�[3��mf�f���^
�p�#�C�+���٬��۬�BS��b[�-���ck�����b$�n��<��M}¾���A��\>�o�G���!PAp��`�T��7*{\�p����M�& �A��ö^��}-�~}��߷����_��w��ž���Ύ�zI/�%����� �_��/��W���w��������>��w��7��K�c0F� ��*�Hщ�dC��x��mc���q�v�Ìub�+����Xڽ���3v�����i�� �� h�.Hmt��`#@#�PĿWA�G�D|H5ٽT���� g��������N7���X���m��":?��:u#�0�N������W~�rW4/ۈ�+�S�w���a]��2@#��0�i���:�V�~��e`�hyJ������Wկ�7`�dU��0hv<V΃�9���M&���[���Tw�`@^������R~�1_ �X�Ù�`4׹tRSߵ�Bp�#��'��g0BN݀b?/؀��?G]{⃷U�]9�*�e�����;KalͲ���q|#�%��"��U��ҟy���+�'2����*c�S��з��z��]��,�ݝ���J�K4h���خ4$�8�N�+Ƿ�t:���-�+L �2��ʼ��d�����u��W����;0�Й��r`�P�xL �ڲo�]�l\	3�B���u.���C4���$�	:�,ǩ�-L�(���Q�*n)$�d ��T��Lx�K���JdQ_�'TB�Bsz_7����kq�c����w��'β-]Q����)��jW�O�6���?F[j���
y	Ϝ���W<ʹ��	��K�|���IV2�(I�m>�bY�Ӟ�����k�Q����'	W��!��"�� ��k|������~���D����-�i��!˽��䬩lT~���{�������K��&X�Z���̿6s�r)�[1�P�Ӣ2��h҆U���l��J�E�He��7�-�r8�R��l�8�@��k��|Amݽ�JfeAӑ���(��Ek�T�ԅLUc)z��9�~0�4�ū=�z< �z-�R<�ٙVoE���^Pڜ��w@�(��NK/�G=�I���������6J�.���F^��)Gxf�ʛ�dE��,e�<ѥv�����~�h�(���[o����[T��VI@ǝ�.i�d�_���l���^?��}и�Ji��X�n�H�NtP�kW�2�/����r���!*�ɴfj���a澢n]c=b�h_W�L�+�'[�y<-ڝ�
r-���7�t�� o��"�Hio��g������Ǉ������V(��Ӗx�$cY��8~��|`>�9�9�oȼR�:Jdy��`������Z��w�\�*W����y4����6h^lTm�Ud��"�2�������ǵת?�� �י�޷r9�By�!�]z������?����w�]o�/���[{Y �^�Kz&�T ܔ`=������?��w���������ſ��՛�zڮ[�����k��8���@��u�v-:0u*Y�UX�6���S�	 ��+g�WҎ��﫱�p�� ��Q�������I�n���E V1rA�s9v�y�.�lx�۟m�[ ����]���d,^m��\.�ot?��
!���mIGtd����e�� r���P����N��z��,k�ʻ�tG`�F9Gy��9) ^;�,���ϦU����(S뙂ʉ�� {櫖��b��x7���񛵓�`����ǽ�ʣ\N�uRk=�B�ȓ�Р׹���rΝT�`�M�e����� _v��mo;�����J��ǕC�^M�U�� q��m[vf�?q��.�@ٱog���B��a���w+��ԫ8�cP�y�/�*��Ώ<Vyj�����[�"�Ux�Ĩ��r�w�@�P֋�ˊzw=n�s-���z>܃L�rq���R�7P���v�9d߃Y�h����޾�C�6���>c�u�3�Y�lv��;%(/*�i�X���@�ƅ�x�k����v\�/��e�)��w���_�3(?�՘c������]2��9T�������
�t�i6����K�W��,�;�]�Yo�c|3��}�)��h����&���e����oޥ�"Ƒbp�2������������,��^>=/ul�6��^�zY�ճmV}0�A�g8�9�`Ń��'m���.�Sے�Q~ur��r��#A��cN:d[�n;��U}���x�w���F�j�&����'��V�匋�V��;ښ�b|��p��Elb�k;yʶD>�)VgJ��ħk�mM�;5l��F���]Vr>P�z޸�V���sS�o�؎�lf��d�lO<�6�"����9f4�슧Y��V���uR��<�~�>b.2��L�r9O����#'Ѐ�d����#l`������YĆG���d��Ox�u��x{S�-:�}+�}����\��GsW�O퍧�u=�����՘W9e=�st�>اo!/(p��%�3�J�Kԉj?f�zF۫�-ڥ,WO�RǩO���Tn�7�e1��?Ȼ��������:�����q���}|�s���Yo ��}O>d<�v	�0긜tl+V�]}��<�����+��
G�i��m�,�YNQ���bZ�I�)ev��!�j������ �ExiIX�F�SV�WZӠ�(�k젾�bm���U���	�'��ԝ��M��i�:�B�����㐪�����a?1 b��HW�*��At>Gߏ�\�����������Q��~����7_���Я�ޫ�ˏ^]^}��7��e�KzI/��u� `_�R-��������������/�����q�}��Bj�I� *��r��S��:�� QU�#����U<��z^�ms�`N��F��DuCPD�v���(w �a�6n�#�`m���E�z����^�8�#P�k5�K��@��jIΧ�B�G�0�!�K�Z��S��y��H#,ь�ү�c"[�s��O��:A�;"�69���Q@p{yp�����e-�jԑ$�)By)a_|t�?R�3J��62�U�9訓��̼$�zR�Ӵ��<������]�k|�׎xA��صmQ6ɋ��Ҏ��y����W�:@_�}���-���<�N|��^�o|�		��~�����2�v��!�P��B��W�V�x��0�a��Q>j���,81��=_l�lϑpg3G I��<��X&���� ��F�8�N,�Z��ba�5�e8{�m�#�����}7��i��9�%�S�~�_y�yP ��@��!yo�.r����&�ɵ})�ȣ�YF�#�x�p��\�x��(�-�;vF2��<�qِ뀼Ϝoq�Y7�y,�V�¼T��/��Яu�qE��8IG��|y��@�X.�~�;I7,��8�
�$d�Ejz� ����J���:�:ʄ�����S�j�f���2B�ş6�q� ]l�I�clJۻ��ku>���,�|e��㔳�����˓b���Y. pLCz�q�zdd�Ҁ���y�َ����ȵ�N"۸�TΜ��C�C~	��A&�>�<����.�ADgB�+�]�\�KϣX�%\���2컅|�8f��x�4C���&O��i���ihDٟtFM���-�]����S���%����C��	�� r�S���6���`s�_�	��~���7���:p��k�!�~�4�W��݋'n�~Ԁ>0�ow���u��@��"0���)���e���V db����\T��/���:O0NQ}��Јϧ�؁��eYq�Q�;�q�S'���?�&�8�<�z��z����d0"߱�hoe<A��U8<.��M��G�G<-V�K���Rx���t/��;l�pkP7���Zb�(�d�M��DK�lm;�)���ƒ�mP���f*�}ి�^�"��տn�7���[|��qD�8�r��p|5L?�q��<�z����NR�1�D�	���Q�C���݀��լ�twh���>��Ou���$���;9N,�]�%`M�)�/x�}ۣ,�~Z�=� 5�>�{x`Lο9�V��Z��V����0���^��p-����~�q+�q�eg��._��63�]"8��Nkcf��gnˤ��䶃>�7드"���?��E��߯72���|u���!�K�l���+��}��<<�G���!- �s����1O������y=��ԏ&��c)�s��u+G�\�Ʌn�z�t�s�1���u\t�;�X-(<�;���q_�R��@���ۈG��ʫ���Ko��݇w�IЧ{%���Aߌ����]�XmA�_�O��)�.��·�W���a{�5c������������>��z��%����l�Z ������׿��￹n����ۭ�iV�(%x9l!&��K�x��J���0O���D�pz�C۲@��h���] `(�ƨ[�`�=�d�ۅ�} �X��� 6�P�ȩm����yE'A�
\D��㚞3g,e{��3��t�P���#��ã�4N��>A�`���D���0��@m�K���dwZ�tr\#k<�N@یaQFw$r iSP�����̬W�B�r��Ϳc�iOe�I�E�}ҫf٥3 ��Vq�� ��iwh� iu�Z�����%NX��ómt����eC[��W�lq��y�U�~�!�O�Cp���;$��U�U$`�yc Gg�Xo��s������b�S�n��;�����:�|'S���t]e�y��޽k��#�+a�+d��<�U&��c�Ά�m�����,�;�n .��cǔ��wR����1i����끻��x�M�~î�L���&��iG�n�L�����8��@�҂�m��J�F����@�y�G�Řt3�no}�w�z?R��o���	0&}�q�=R}L�
+}\��-8�2�D��;�F��xt�.p��v��6@'Eզ����4�ŷܙ��Wߏ��h+ǖ~��r�����й��_��t׍���X����Η�Q]�6/1������;b-���֓���� &��핅��h�\g���BQ�܂O�e��P�,�=@�'o��h��v��;����{�w;�����|a+�¦Ao������6��9�Y�h�3���>�a���@O/��A����T̓$��N�UMj��k��BǼlWqe<S�d�����b^���<��>������I��-@�VO:#����cƙ�yW�.��c�m1�('��v�4�"2���E��	v��7^���bI�O��c�O�b� �1���u����*���iS�Üfz���ўu,�ؤ�9ƪ�̘J�D�[�SdUi��1�]��Œ:9��Q��=Oc���A��O�:�;N��&;yeA�d3�>�bK��x�/�5�g�S�����h��3�.&��|`��$��Ϯ��O�������^�1��n��b��7�'`��,~b��8�-/P?�H\�W;+�&Sy���r#�]K�`.�2}��L_����S���-^�DWНst?f2A�slY��X�q�l���T�JӇG��K�yٙз���q!�e,:b| ���xh�jZ��e=^}����~��}�xZ�����z�탶�e�a���ƿ�{�����P���ncƉ.E�-N�S�q'O���Wy ���x�A�汻�mڼ��f���q������z�C�
����2곔7�;�u�'�I�X��/C�},�O�eQ�e��Z��L}D�I\����r���x�?�T��Oc/,���h������Ǣ_�Ǝ�M���)����4���z[���ˈ]�'�פ�坦�CU�Ԕk~�3��b�y��N��:��(k����h|�o�h��R����ظ���<]��c��Ȣl8$��f��؄�'�T#A���S��������V��כ��Q��KzI/�%���e��-�ݮ�7����϶w��^uS�=�z���5�$s��F�3n�>=��Ե�UdP��i���]���d����LF�}2v[�>yj�E;���v��97b��,t7�9@��[;�td��r���F��A�,��I,89z��a�:��l'�EМ30�82��!���2I��J,��� ���j`�N���.�y��O�?��I8�8��kj�*@��WC:s�"��Y�ӽDh��4ЋZm[<o��<P�N9�C��;!�O� un3�=]����9��e�La���_ݑ�.]����m�N��a'��W(��3�e'7�;G�'J�Ad0��
�\���M�}�/��X\����p�6_����1��K��>�VW?3��1�^��L�,�<�6�Da �H}������V�n�]H�q�@��m�?����V�ݾ
ta�;.t�������ü�6@wRd=2d���Ųl��1�L'V&$B^կ*w� �I/u	�']z[!S��_�HZQ'�7�U�&8�[�!�57ٖ@~A���ϡb�ڿQ�/F=rZ�-�{򝼍4�A���1o3ep������1���%1Y%�(��TNF� S*����q�e�?d0���	�00�/R��宦���cL�)�\B_�m*%ٽ<�����b�o�V��,bO�|X�}�'��v��Xd!���G?���(c�.��m�A�ls{�m1.��4y��1�&mW�-�~�T1ζ1%Io�Y�W��6|sݪ���sR���к�"&Rܢ'��6���x_|�~��4�_ԍ��8=#�pZ��k�R�;���{6�P?(�VY���1�u��8�)՗�q҆2�'�C���,���cRy5�S�&{?N�r��fB.(/��&8��$�GŖ�����ұ@�z�}���1����0O�c{7秶��L|���ѿB������!>�z4t�ʁ�T�$cCN������lze�O|+օ�Ģ�1�
������j劜�b���K+������"�����?m�l};0�|M�qs#>&/�N���c�Ԩk�8���!^�Q�TZT�uBs���3���p,�c̶0�N��E�A?C�At>GEܧ�S|c����_9�G>��ǁ����E��O�m��l6�#�]�ouҞ:#����c?�ݨO"�?�?�>�/��m�K��~�|����C��x��ԶQ��t�+.��[��Rwģ̣]�x'Ɖ��q	���TG�ǎ8Uy�]����xU���t1���;n��XT�'Rֹ�]c�c����:������ _1�d��,?���u]�<�g����a���E�gی�	����YNg�QǗ�B���1m0�I�j75G.$�@�^�;g=iט ��7�~|˹��'��]EGtS���\I����ďa�����N|)Q�Sq������S����8���Q1�e��q�d�%�{��v���c9<C�z�������7~`���w���sA|I/�%�$�)/ �=r��{�����?���������z��/o��յ�z��ق�ű�j'	���^�Y5������ة�nF|��l�p�eU<�'c�V���Ν���c��CylG0n��Ў	�ʕ���(�v������4<{��_fP�S3���js�j��^�zEA)Y6�x&i'�2��T���]I� f�:��C�� {�{��{4i�-��7 � @���%PK`��>��;o5 0�����_�wNr�
HqF���L~14�ϔ��,?��ѹ^ש�Gk��3����W��ۤ ��#y��7tV�)p6 �˫�s�y��JfL&ug^A����r���h߶u���6�X/��w\h�@E�:�u�rj%O���v�6Fi�I}���͓�Ǣ�w��w�c����>���lֻ�,�L7]��q��੶M����Dv}�!+^�E��	\A^�	�
��2�w����ؾ�}��}1��NA���Z%�ټK<�|�u�Q���2�9ӕ����������y_;�'�r�ye�� $���g���+uq���Y�0h�� ��� t��^V�RFmUdk�9��݃a�ͪ��7PW�L�������d Jlۇ\^50F}��a�y���+���3�<i�
��*�/���j[����X��YҠ�D��<��gg�:����S\�y���_�Y�]Yg�N�J�/>��q�yz�VP7���rV�4�1���������!m�|>?[a�8iۨr�y�βaK�x�	ˣCޚ�#��'f
��*iZɉH9.#"��uc�2N&�o�.��ϊ�ږ���}�}�1�Q�Q_�Y>���vIu]�&�����tB���?�����l�����|B_q�9�c���pT��b�џ����� ��|����g�n;e������y?�Gma���l�<�.�ԉ^�7b�n�����mL��,3V��D���=��Z��Q��a�4V�1�O���:�b?F}
;0��V���x.��6��T�a]t�y�ߵOԧ�����p���yb�6�;xР�	�N}�o^�6OY�����>�pB���<�0�������`��<V �ߔ�.Vw�{V��xg����C���z�'ŉeo��žu��A̶a��UZ��:mE�t�Rw��vͱ��t�
}�'�r4�M�$'[&2b�������4N� ʇ�5p*t�UG����̸��HkD��x͌YXϽX�y��:C7D����b
]G�!kk;��us�Iq�r}�c|P7��P�����F�F
Տ��C�X����rl���7�&F1���t^ �q��9ڧ��y��煾*�M/�����@����m�|&M����}p����S��. ������mj�v_T�6��݋�FA��^�����~_Č�/J?U}��<N�l���#{�b��w���l5.b���b�Q~���1q�Օ�����r)����_�������~���W^}��޾��}��h������^�I�:N �����������_��[����{��c�n_^���#>��_���6��FL��ѱ\W�臦�uW����+�cׅ7�(����@���(Z`es �T������ҏ�yu��[������)n���d�]Z�#к?tPeO��f�/}��Nu~б;(0R��~ހ9�޶|LU+Սh_m��p�
���jĸ̽='�1:w	��;�c�F7��*t��$[N|1��z;��(��]�1:$<���N^Nh�m� ���M�C ��]�k��A�)t��]-+\�w���Q���a������&�'8�_���)H��D����Dڋ�I�jN�qI�~ ̀��H��:��p�}��>�-���w���.N��c�t�/�K����O�����뫗�A]��'�;��A��5��{���1�~���r�������ْ�����O�Qe�]	1z<ۍ�H(�s�����?c��T`w�o�17F=�E���Y����q��瘸^��[L�@��UC�����g}���wX��y ��`<�a�뼟ː��a���u��ɢ����З��^f>�3�*�*7:�^Q�R7�W�A�k����
��$����0��qglg>�������ܬ�=�A��.�~�3..@�w�h�N��Ѧ�M6<�����>A�G\�Z ֏߶6���׻�I�W ,�CNf�o�ڞ�Х���P��3�֮=oX��I{�r�k��r�}z�n�#�X�g�����;�7ȶ� ��B�Ѕh�p2�d4���`ż>�����ȇ#�{=�n󾰫��!�Y����6�D��~����+�%s�q��>7绖�:J�.�H��L�qn�e��թ�^w���H��ԧ�q�Z �����c}�}�A�L���ú��q]t�zF�d?P��R]�2>�|\�h+C�J�[�N}Ⱥ�g�emy�alo�Q����Eہ�[�����m�W[�����U�F�a���'�tr�r"��c�-& #&t�(�j�8F�����\�D��ō3��c��̋m��1��耀/�S[Lp��mvlT��T�x����6^��j[a��P.����N��2&[��Æ8�]Qq�;o�/eWi;��΃����ܺ�62�s"��2v<c���Za����j�Z��kt�qvm>Q�u���;�Y�d������0�#�4�K�`�ec�Z}�'a�vі ��!/�O}#��+*C_�D�>�㷐��9's|(v�CN����v�|�o���G��XB�t<�����c�}�1�O-C�b�p�	�ѝ����ǂJ�
��\6�w�gq�Ȥ+|���\T���b��U�]˵���c�R�{����U�C�[�?:�f�/��g��s�vie;��1A�����$�T�Xe�p���4
`�vNDNq��Ӯ�;�:tЦ�t#�X�Sz�:�7�.h�t ����t�#aE�/��z"�n���������Xx{	'���`̈́C������ob�'�N�bI��Xļ#]|7�1��2n����c����XAu�MtG�#<;lL��y��ʏ��J(/b�lS�q5��WM|/��c~���>0@9��2\nm}ẉ�d\��({\=������:t���e��f~ň�(�c�,��xb�2ڴCa�NB�e��}�*��������ƵR�1�٧�?~�7���o��_��?��?�g?������>�/�%������������������������iܫE�]���2v���Q�8:�t��"�6	��㔯⫴�g2��;��9�g�ňG#� �H��m��(��޷͕4{<�|�.�6��8�p�c�-��:ũ|.#���}BԱ	�h8�ٖ_V*xPЅo2���d�d��ͽ|c�@{t�J�ߝ�Mg1:q=��v`�5&���2�Oޅ�W@�`�yb� ʇ#��L��4��:��:��t��e&aW�;Z���w�[���N2���}�v�C�� e
�"?sy��Fw(�YLuz�'��9P�� �u��)�T �r���S������h��*��i��?�� �i���<+�=˓��v��.�%<+����g^ю�N�IA���Kl������@0�XgrE���s�no��P/V�_��8!͠����?9� ~�X�y,|�z��1��ΘX���]�+^��(�Y�~⤕�:3���?�d&�����|�?��c�6	~(?U�O#'Pws8E��6��o9�����Vb�ȳطh��S�G��E �N�+?�G� �}l?l;N)��C9J7�¿e��:�qeRouG���.s�q"���T��O��v=�M�E�('�Vd��n]�����W��s�+�$�C`n%S�~ա۠�h���7��:)!���� P���>�(/Z���k2���Xj�源��+�K_ev���.�Xhrq���^:�K����'�q"���˟%�d��l.�+����y�::�gm�_||q��$|˓��B�8��y#NT��e4�g�O]��]�[���.{���۳���#�;�Z�HYq�jL��X7ڪG���0�8�Ƃ@���]]�o��G���C}*��7f�QW_wpת�.?����;k���B]���s�}hy�|�����M������w]��O=C^G�>�kL��G�W8�A���o��
Q\
\勋����q`�a9F;0��츌uV���i�c
�d��h�M�I}��կԀ�RƖ���<������F�>]��_���.�Ӄt႞|����<S�/�	�.ʳ����NS�ßp�GT[N�+�)���3{�H_�rtlF�i�R����D�S���G��7���c�OؤҦl@��!���.al�=�^��S��,F�a?GlI�5q+؉N�LB��i`��� ��^_����4,���u���"{3���.��cQm���̝gɆ6�d�b䕑�1Ϻu῾�,��rY�aW~;h\�(��D���	u�F5�.AWƱ�]O��VK|���[^t@[�����j�ո$n�ZG���tv�M�����a����X�c�],�q_�]��d׷�ڄ�~���#�~�l�"G�B��ϝ�����qi��"���ݴ�(��.�@�ƍ�lԨ�;��y�;��n\��n?l�����W�>~���ɛ���jb�KzI/�%���� ����f�^�R�z_8��]�c�;E�+����N�n��S �8�FЧ,��WxA�:��<U�P����]_���^v�m4t�oۍ�O���>��q��z��r�~km6��57@Ѱh�%c��!@���6i���-��h<�E����� �d��һ�O%����E��9N��Ru��}4�抉��l����s>F��g��6է�I�� �}�'����,j��?ޭ�+�ͰB*�Sm�_m+wأ?��������n �ar���6�e�=#[D0�~���00O>R5���4�$b������$x�w@[h�Y�@��Q��0�E��wg������,ٌ�2������q�/�� ��uG��ݍC��-�T�B�(�{*��~�g{�XdЦ����+~���pL�q���^G<���:.�1�P�jr-ta�3+Zfܭ���������ڶ�s���T��PwEZMdb���J7A�P6j[�}�1�Uǈ�c�2��=8���V�z���;�l�]Zd���5��J�����%S]=M���Ne��2��Ad\���*1Л�D��vu�K�Jq���5O�!p�զ�#ފ��$*��G��]Ӯ��Ol�UU��+$� gbj��V2" ��|�n!oO��ڂ�}*���,�>~@��ؘ���^E���I�{��dO��Z/�Z	5y�2��^�Ũ����;��^�+i��4P��k�/�2r��f����3ި,�t�Y�T�gx6c���0&�ޙ!�W�O�0���BsG�'R(���#}�	?qOs�{�W�;�nn�g���o�7W�4)/��趾����*���A��+�<�Hߙi�`-]��=v�>/��E��������*��Y�	I���<t�e��*x�r]�)<�l�UTo�oR���+�!ڍA�Pa�`kXn��ksٖ�q5���.�Y���(׹>�+��S���G���'�.}�ܵV��(��4�������fÉj"3��xl�ՏnR�l�&?B�vD=Υh�6gE��qe��)g�=��Xw5��2���yD�'�\3/��ա�6�8�Ƹ%^N�;/�����L麠"�v�'jY��j�<tyײ�)�L�wl�Xp#�J�b�qW�@(~��$9��2��6b�b����2�:!s��f���h����y�OO]�1>��I�t�	�OĢ�dH����G�/�����u#O�z����1���]O�y��D�um�͊�V8�)#�lʯs<��^���9��1���O�v����S?e�o�/��:�.��m��/�3��QH_�K�-[������aӳ^�\�o��ϯ7}SZ�k��ۏM�����^|{}�w79���c#[��rlpx�o�,���X�e\��4�UŻ`�pGfJ�K���0���r���ȣ~��6�@��/�b�������G�����^Y��{��	_�KzI/I�ױ `����������o���>���/�X��`���G�7�<��*Pt#��;��u��(k�G�!XPVo@�a���9�ר!8N�;���A�V�������n�>�~<̱���>�~#�xS�e� �/L8��'�\�3J~E�nΣ����P��Ƴ�2�i�fv'��:�U��/1�E�{@ДA�1��%�9$��I��v+8T�@1[�4*���39*ո�����PF�@�a�b=�KA����^$��~��(�j�(��SJ�_�O�Ѐ '�������{�㴌�y<Z�J�,KO��!�I� ����с���x8z������:`w��I�So�n"OY�Ӎ���>�T6�{��Q6�ü�>�������q�΅�;}ّ0/�H^����ۈ�W�K1�\w��:�:�q�"[T�qG��q�Cݫ�N�yb}��ח�AW����͔��
���G�¶́��L�G��J{,#*9��ڻ,�m7�Y!�]�����m�c��g��R���w�'s $�4�ƚ]��69�|��/��N*u
�g|y��.�%�[�X�Wi�9X�O�e���'n��u;I*A>��F�kM ���1Q�� fƈ`��Il��.�M�#ݽ6���[�-��b�Q����\Z�]4�D? �;g�B��[[__F�t%�P�����u2Od��D9��Kۖ��z�J���2���g���m��C'�������,l2-~���M:.VX=^muZ�'���ԧ���x��qa͙m�;���x�}��+���!㽙���m���2���G�oy"ӗ�>�4�:W�9�M��,��ۀ\�������z���Ś�L�b��7.\��o�/��㣬��� �q���i;e��(;��;��a�U����0#�bi�T?D"Xz�s��WK��:e�i�`h��L�t&%˿Q��=<ǘg_�QN'xV��{�T�Q^ۿ�b't`����}<T)(�4�O�jK��v�|V�+�n����C>��ݹ-�Н�\��M[��`=�.�_���x��h�:|����q�Q}��#�IW����z���<Lv�F�����?�_#n�Mi�<����}!��?�y�X�m�J��|J
��)�%�65~�<�+w�'Jhw�=O�Wi�6�7.X�6���nש}>�J_tԴo��1�y�D�3�5�)�,q�b��
1k�z� lQX�6gU/�)�|]�'�#b�9~��1'�j�g?�a����Z`�})�Tw|�rV�K�G�]��g��̇N��"��/ケ9��Y�!U~����R��G�`Y��f%Б�'ڒ�߀~d,�c._�6�}�,	���{��͆���,9�u�1����aOM�B�AT7%Y:��O-�mgi4�6b̆�	��������^��e�{�'���v9�g��Ug�ַ����&�>���!7�^�����==}f��K+��#�.cΨ�?�t���5�+��+���1�QO:744���4���1�u��g��j&���:ҁ�.���}fo���'������>��{��@�����^RH?� �������S�?���_������=�}���ײ����#��~7�ف��2����F�+��J�8Z�: [?r�2d�bt6��<��\l?�����k�����ό��`�P���_~����o��}�Xe��ɶ77��ۛ�`������]x��*�FB>ͻ��s�rW��� r����l�o����S�<�>Ob*��$�g�w��c� P E��#�p�3�Ř��4ѠG�+-h�N���l�J�>���u7\�ۭ�|��ǎ������c�B�TZ��O����G��<�A|^�G�aQ�^��o�/�� ��:)G^p�h@��W1��6��C���#�y�qV����x���gI=Mr�r=�,��,��|w�宧��b��!_N����Bp���cU}��>�GҟM�k���R0s�5(�g�m� ��Sy�cW����W>�#'��S�;��1�Z��=U�����o�5�>�zn���l�(����Nd�C��e�v��!ǳ�m��U��*q'��]�+�`M���9�·^�1q����Thwq�,wԍ�V���x�|d�-�T��=��軩]���������|E�bL�U	b�V)'���il]ӣ�����o:�Z�2�rHVpL�i5��i�d��%�܂�/ �W�bv��S�����^�]D�l����p�}?��U �_V)��xs<i ��Ǐb���]3�c>�7`M��C�\�S�_,����o8v�R%�5c���6l��NSY�wA�+5�]d2�a֣m��L�!�,�#���+�c�٧z�6�_��z=ʉO@���K���j��e��^�������P.3����O>]i���x6Z�z1��z~4c����\��0���^,�վ�B��D[KYC=z$��7�	�yi6tg;�6�iv:Θ�`/����t�^O�]��(:���Xw� S��U�ˋ�4�����Hy�|��3�Q,�z��
A{����Z�_�^�]r2��u����C���W�D>��7֋c��#]�}�7�R=]W_$��Eֻ`�!��olT���IK�^������aRWh�q®���nb�ܦ��ĵ]�#�S&��k��x+�X�������ᛣ���]�v���zF8��R��)�h�	=��l����ا��.z�5��x _�)��DO:�0�{�{|������B�c�c7nfR+L�n���hy����+��.��m�f��^l�n�XO�"nHc_N�Du�1�1.��<��B:��X��xZ;"{���ܯ���Zj�}u
(dR�wl/���l�'��k��b�2ɪ��TE;e^��2��Qΰ���'KQ��v�8�m�F\��0��ZbΩ3���B��h�n�;
<+q�YŉL�}�%����5����'lk��h^Kio��̣�1"�b��u;`�'5�=��KI��=�G�~˼��α�K��������ǜ�/|~�Ҿ����|y�O������������ګ�޳w߸�\�­�ɰ�`�mY?�R���{�&g��@�|������4�%s9܏��k?�)�D뎛�,�ul`z���t�+{��}`_�/������k���o޼�����^�KzI'��8�������#�����7�������KO[�������X���Ǩ���������� .���9����T3�'�Z����x8�~O�0\�i4w�7,��A��/}��>�k�/7�����g��={���~���؏�����|�^�y�_��/����r3�����A_��\&��.�Ы�&�5����#�ꢚaO���߂��S�F���aƏ��ȼW���w��0��=��E���x��o��mS�hT*��而����ۏ#�@{��Y�WW*��$h��j,*Xv^���u�+���4�1�uڲ���)�����'�f��oչ�$�:z6%��=;psP#ʚJo�r�w��|��馝����w)g�k+x��yU�*� ��mнU���$��_b#�=U��|����� ���4�X�D�k��t>&�*��08�UN�擽��ч�*a�c��:UV�x�� ������:fb@J'H��p�����84�S�t댺��e�)�,ԋ��|t6��=�	��GY����@V��ŉ��P�\�(�pB�8�6>��_�}��̢?����cb��uEh�9����i;�t� 8����@�����&��V=�,�2�^��9ߺ���M26��v�*�*c�w	��h�4㢁"?�Lƚ��
��������uI�g�{����̙/{�q��8q�b�@���E���	$��5 �dq�\ �
"�(R��|�P��#��g��x��s��Z�i��U��_U?k�1��M��>�ߵV?����U�������uEk����2_[Pe uAn�$@/-�%��0���gՅ�l���岥�ăU6~�}���P�����Q�.��VM��S.9h�cR~�'�Syx��̗�S-�w/�@�j�菾Ϲʋ����P���w�L��9n�=ǰ;��sP��|��
����ό�0MZs�6m���w���GC�v{����_H��|͐����]l�;!Z5ۘGh����Ӣ/�''"ш�Pﰵ��-�R�2|M�ɰto�ǇmA
��<q��w-�Jǂ�q �� /ZV߆���-prC�:��~H}��8�&/hD=�����ڇ%�}2�\���V<ϲ�#F�p��F�0��;b�$���.��ϋ�q.��I�U,"��(�gG���}΋�	�}���RN��c�:;�7K*��&c�:.�W�GS�f֛c��$0��M�����!/|���Ⱥ��,X�g{�x����|�r�!�����m��� ���:�7�I�D��+cH�wp~Q"cl6�|����Y�%,�c�q���3-^��e��.2��\&�Y�A9����>��~�xI�ܸ��a��%�͘{��>�+�����}���~B��2�7��<WЛ���\Ƣ����s�I�`y� ^�c���-��L��.�t�����`<�Qd?���x��q�K�ߥ������Z�k;lw�I�ϧ�����(.��P�=�G1��u]x���	v��WM6>)1����o������m��:�ev��{l��/�J�S����_���O������W���#y�����~%�*����f����^�X�d�|.�f��}!ַ�Қ��4�{��K��&�����a,�[\N49,�
�@��i�,r���;y������_��_����Z{�ʣGO�n��������P �J�����ӏ�gw���~�_������/=�.�g�m�b��� �]A��.\�k\YV�{�h�%��yDA(�N @��vD� �f��"e�k�{��q��Z�����u��뻓<|�-Y>�����|���[o�._}����'��ᵅS�s8���J�><"rX�0�bv�¶�/m����˺r0>�/;b�S��e*P�E�>ŝ�
���������f�0�,��<�c����q3(�n.W�G�c���Q�L+�_��G?�3����^��S�cZ��s�8�}�>в�1XJ٠sJ&�z�j}}�k�*�s�Q~�M���j���,�X�\�+��<�� s2U�_�}�3�IR%�S8S�L�������Y�r��'5��9J2�L��ݐ9Ҷ��ѫl����g�Q7���\� ��``�p��q�a���݈Z�������<׏v\��(�}�6r�y���A�ߋ��4�zܮ�=�gq�?���x�B�I����;�"`�� �VLD�[�&��G�P�q�2�ﭗ����j�ys��4f��f=<D�^��VlO�cg�����sh���@~&���e��4g[[��V�e^U˱�
�(��)�E!kQ.c)�`Q��_����Sn̩;�Wi�i:F�.�ܧ���g�Ǹ�����B6ϧ��x��t�-��u�]|����̟�àK16ܟ�G�.˱X�m�_��5�^q]Ɗ���%d\�Ȏ?օ�9IR��ɑG~��3��e�h�m�SO��z*���Z��:�7Ȉ���Y�uU�	HR�w7�NX`���cMW�������G�:�����ɰ=Ѣ�A;�'��0�ɦc����wF�>oӒ�Fpx�lA?�z�aw��Cv4�|�Hu�b��+��"k��[p;���,�<�M��H���������&�U�Er^���;�zD���MB��
��Sw����~3���8�Ez�م��������;^i6�� ��4���h�]�3�i�mCB4��)	� :���xZ����d��M�]o�1[�����d�Q�Ӑ�zHc2f����?�X�*#������!�y�U��iي�T��=�\R����y<_�"�8���{�7�a}󿱨x�8�㎞q��?z���4���I�-mjlt��mT�g�	�1��?���z���7N��o��񃮗���3�̼��d���S=1�Q��!��H��	��e�жq!� �+h>��8�9�����a���i<���#a:�h�!��XI���5�Ge�z����O�6Gc��<��¤�鴈#yJ���w�=:��]��$��哒������-����pn!�*�'Z�M(�������t;����K���o�?���K��Gr9]�k�J�lc���]�[��#%|j�����ɋ�>Ɔ!���Sk��_��:�4��N���������}���W~��U^��_����o~����w���G�_����������	 {��~~��;�|���}�����G��m�<ﶖ�A���7@�"B�Q®枌"���U
��Ѩچ�ہ�F���0xd�<p2l�չ���G��g�B^��ଋ���&���q{"_~�]y�����ݝ|���_";0hˀ���p��08�u# LG��R��, ./{ؑc�fG,�1G��9�O;�G~�?ح;��7Q&�tԛr_�K�����#����J�3����*�\�ag>3@ʠ�eg2��}��@Mė1� 4;Y�� ���gHګ��ՙ<^T;�9m8�r�o-�;Q��q�0r�G��:3�v���E�&_A�U8<z�J�\��D�4�>N���0�O	D����<�EZ�U 8��v8�y�����	p��j8�U��fOi�;j�����3;= �/Ƭ��q�Ņ<�����m�ys�s}Ѷ�rD{��U_{�������"�	��9a!���VI:��S���Y2�u����g_��$�,���тa���9�Gց�|Ic�����/ ,�M�Mt8�����$?�?���t�N�c}q���"qB��,��>r�5���Y�7�Jy����r@LI4U�Q�z���b�\x���"��l0o�~[�n��K�S�懏�<��c���;�H7��Ϣ����$��ޥ춍��k�������x̛�=n%�fl�r;[�w[� v��y�>����Xⴒ*��&��$��o<��cz��Y�y��Ω#LX�Q�X&�������.��T�%���ǈ��~,��*�@S�.'Y���`l�o'{C��w.ռ�e�D���G噆�7^�~�i�;��ec\S���f����-�����`̡��7&t���]E�_%�u>m�N��3�%�'���Z�]\��(�;_�u�"\�q�.tU����3�	U�����ć��
Ǻ#�N��¼`W㕒�H�~d���vp�Oa���8�,�7N���P�P$�5}S�V�
�[b]l˓�	��~g���>J��]l'a7s�[ON���y<����V�>��t�B��;Z0���SV�Οk[���� ن��ݫ��(��q�Ż�������H���/�لO�Z(_�}$C�1Ʊ�b����)m�N��#y�{x'Q*,�Ӽ/�>�1�9�4��(�1M���e&\1j��qj#�L�c���))�������D���R&tNđ�6�>��I	�k�C�,��"�ƌŃ��]��=�׬k����n����ס?�������c�Ŧ���%�&���>!|��'�C;�C���1k���V���+�����/K{���_������&��E�%��W�v�����>�˽[��V�m������lW��lN(�f}g�"('�r�ZX@ƭ�w�}���IC�:޸��ʃ�/wO�z��ѣ������O���كu��?��?�Ϗ�
 ��U!���>���O�\�/^l���N��3xa�"
�`E�GQ��~��i�́njx���ۻe,��Z��f� w�dP�]N��������f�JSpDFP� �^�h�|���N$�#@�K�gY��y������_�G�C���W��Ͻ~��*��ַ��Q�h�qk�q贛I� �Zv��C�GojU�^����{���gg��$�F������v��m�;�P.��@���A�hr�m�A�!��G�U OX��EW��m���{�Wu6ىi�v�Z1jF@!�:���=՗��ӓ,���9*�Mq��W�8rٹe��_;rZ�ہ��Sf^t����:�6���dz(S�t�Nɖ�N�}�2������V�cG6c��N�/0C�z����4���X��cw���K��h]�A���1��'�������<�����8}��Qv]y�p�0�F��t��sO�֌yq��>ο�i���^�t�pHK0�����b]�N�S�G�7ϓi�u�fЊ{�36�Mb�[���#�ʎ�A��	"U���+�q��b�n�|^H~��B�]O����[�'�����<;f�2���}<�B��ؽ4�W���4�ضƉaKX^����z�� ��}������H#[��_BG�� ~�Mb<��F��S%�w9���w�}�u�)/����Om?���� Y�y�6��z�V�z����8,�R#N^���1lJ,F�E��x~fZ�{Y���K�>�u�-B����T��e]���L��2�v>�-*�dK��SY���.�9�!��g�T��s�O�֞����m���b3���(�dy��n�����X�f'}���Ao��4I�e����Ty��o�#mԅА��Α��b;۵}Fڰ/�*��ˑ�O}�z�'��y�^�r�w�?b���a�Y�#�<[ʜLש@w}��4��(�_e��B�g=c²��g�p�+l*�j�+���"IY����'F���x�)t^������5��cR���]<α�P}��dY1_�e��@��|�]Ú���\a�<H�zYGT��<���݈߻�ʌ��u�31z���P�
���q
JO�wu3��߅��H?�oy`;0ٯ�1�Z��%�w4�u<�ߨ������H���ֱ���,�5�c�ə�kߏ�$��]g��.k�F4̶;
f��S�ԙ��ʺc��Yo�X��a]�b��O��_�uAc�Ͼ|�<��&�}G����~��d�;�%Ni�?�7�5��ޏ��I,�d~�HF�N��3ԈK��'U�xB�L��2�p!c�9N04M�+���z`���Yλ�u<v�^�	䱯����`rtv#0K�E��}A?���}h~���Ѳ~�׈ĵ0���֟_�K�$�=���o�ǯvy�_�����]'�E4�`�b��� �v\�[�>�v����Q���I���5�d�f��S��-��B}�0 ۳��s�t�|��d��}`����T������޻~���v����s��?�O<?���Bj���w��g_�_��������g��8������ZNwK�7�8�ÊQҮ��Q��2�/�n/�^Ϣ�s,�o0��vG@i�s�D0@�
�X
���݀�1;�M?�.�v�0�W����<����^����7�g������ץ��"��}y��( w��q5f�v��g�����s��;I�ۘ@ @kt����z���߸��٥)@~�!��dP�����v���QYuX�X� ��#�����1��
���
�{���N��{t��r]��*0�;��Y	��,HqHL�C����X��|����[�G����9$	ѐ��o)8�x:���3��R���,�n�(�"�s�Y��jߕN
f5|�e����hu�H^�^��q͋45�(����> W��.�>��]Np8rta�P�2�7�9��3�ǡ֩��>Ţ}�:*�����˹��"�Z�\�v�<�;t�xς?���Q��g]T�x%��@F�{##���Bu�)������.��1	x�EׂWj����3���7�%�y|�v0s"U��Gw;�_��l�z���7��`^&^Ă;�REP<���<F�|'k֥q#�~l�ܩ�K��n��@���5/����:(���A���~�
7�tvZ�f���ݎh�<�`b��c�J�Mf��e*�3iw�"���6����g��K�1�J��PM�2�����Vy��]em"� mt/c�9�(��>j�ë�[�cU�2A���K��<<J&���v7�M$��w��i��EO��1m<V���-[�1�Ʃ�wb��{�fۉ~d=�zf
A[NXe�
}]e���,�"��^D�Yq�
��t�i汀�����/e��c!�!H�X������/T���h<�~�RIOw�/��o �0��/tڽ��n�~P����s"G�R��)I��ϑ�㫥�l�)$}d��>h���*v�˨ͼl\���+��ZW��� .Z+'����r�<�3zP�S�y��g��,cUe_�uK"̶i�xb��Fr���\�x�Lk���3%(�/�a!Zʹ}W0�p�A���'�#H@�-�|cy����VҼp���v ���E�ɡ,����O;�kɰ����Y�Y_׾V������.��XȺ�i�lW�K�8���^���l��Hj�1�Q<#q$�vd��v/�k�Y���2�y�$|�~��<�?��7����������[�~����q�#��1fC�B=Q�>G� �� �[_;?|\�w��3�gb ���(Z���b�<��>[{�Ҩ�i�^ǟq�.���>9.�-�l�xN3�m�x<ꥮ�+�	��s?�eK����sT]�so�[Zkat�~�S$α<-U��^��-0��E��j���YY[sw�_uʟ��Z���ן~ ���>��:6�]�}�_FG��\�%8�v���#�}sz�H���_l�(�ԤY��&0b~J׵$������:� ���ߘ�a'yNb��:$M|g#7�]WY�͟�u�S;_������O�y����~�^��P� �>	���>?� �ϯ����7~�����ɏ_���=\�.}���emJ�.0#;$ (��ƽ��p�.�,��;;��]��&�h��~t ~�O�������P;�rT�j�������\����S_���o���?u��|������z7�Մ�s���+gt��և�T:fp���te�f�@o�I�cs����?�mbY�z8VM�`r�V����d�]�D�{ٳ�k�i|y��/}���&2� ��c|�,=��{ �(�Oى́��c����w�X��c��A���i��e߿��[4�u�o~�`4��<�A��+��C�u0�d�k��VU~�O���yuL�ܯ�w.;�+-tͿ���>��tm��^���.��N��Z��G�6��C���gy�c4� ����$�(�}�z8��Hǰ.� $�f��y�rT����A�j"P^�`ǈ��Ov`R���Q_�G�΃�vsf���<�LI�����O�����ﺧvn����n�a�V�)d1/�̶��ޭ����6�.���"�}'�c�B?j_o�z�?��G�sGv,�5�}�����fd�.ާ�>��l���ۘ"/�F��ʇ�~h�w��;1'��=�hgz��`�_���5ԫt�\9
�QM�F������gO�+�Y�;��8E��g������\΋�G|}�wG�i���G����U�X�X�F�/_�Sig�m�J������Qv,���(1+���S�,�X��^��u�﹞c�Y��^2�i��xW��}�;�=l��e|W���|IK�\��Lk�+�\g�fZ��������ti;��*�Wa�PmY�=x���������Mu�3c��ˑ���(����$Ӗ1�6��4dѴ�E���<���4������4����v߭c\���W�E�7MhO��A=��{��� ��=���m���-�i�|�i���Q/�r�;��1'�\�D?��Ymd|��C��+����l��n�����q��x��o��Lry�0m(��oq�KP���~���N �b�G���|�H�����{?k�b�s�1Nῂ6�o~��2��2a��W�շ>��7�[xQ�F��b�Y��Ĳ���K���C����L�� ���۳��I�4��O�dL�g�td+�qq�;۔J��C�z_�!�N�=�}+I�Xn�@=��{,W�M$���Q��q�_T�j�e2����1��o͙2��1�[0.h�w�1^�Z�2�O<ޚ.�������Q�cq�_�s?'�_y./O_�r^.��266J3=�_y�t�||'�����ظ4��B�^)D�{���XG���F�����`c��l�hM�&�:]��d�X�l�g�Os��������廯������_�w�滿�K��H���g�����y��CM �T�O������Ǟ�տz�l��������ΎJ��,���>���8Fr��f�[�v1�F��9e&�7;�  �F=�f�+>ϋMǠ������� ��l��*��{,�g�=X�|w���<��~������Ļ?.�J�G��X�q��f��)o�z�T;aᆱ����G���L���~�9��y���k�r�~���NDS�k�G��֝ �#en7>����J~��ĻP���<e�h�����}I}f��,����F�>��/�N�9l#�3�2q�^u���UA��[�Ʊ��:�e��F��~�!�Wz�ȋ����7��G�Z�^����쨂��V��z",2�y���u�K������E���<�� O,�7�UG��s�9�Ϻ/;kz��b�N�#��Wg�s�B&Zr!�*�`KC��w5Ƙd�߳�\�;z�p�,<C��[�-u��wo1�a�C&ў~�Ȭ;�|��W]�L��Ϻ�͓�R?Av�׫����5b�ћ��I$��ʋ:���P�ѿl�C�A<<vu��L?�7�rBt���^��i�8�Ӎ�*����I�G:8��j��9��O�Ų��s�9_�n��Tp��r[�Ή�5�F�a|��t�<G��?�c;�����o�1̓����/�;���M<yL'�Ԇ��N��9s�Y��^`��1��qU�������'��s������un��i��x����h)����|�w/��1W"�ǲ�z9�:8`�io�}*���
u��y��(9+���Ƒ^�%٪�q��ӒO,�]�(ú%�W��>�}��i��J���Վ'11n@���y]<�Cɸ_��pw��ZZ��яTk��;ckq���gC�],|��5�X�e]>����+X��c��k��3�z}��+����lG�7����Ҿ�WA����G��Le=�%��?���^�S�M�qQ�KΧrZD�|�-c��1B.��z�I�nNUW{���f����El��N�B[ty�y��I3�C�n�G�C�9�_��[�"x��Iq*]�C��Đ����]�1��9��ǀg[d%�YV1�[�s>Qm�~�/Y��+�X��ҥr���	�?��[���_����FYI�33���<��6o��������\�#��'k}�^ԗ�UF�W�3d�9��)�"����8J��v������(�]��s��_��>��9�OŃLG�1�ڤ��0�9����^�^[�N����k�u_ȸ�t���m9ˏ����W�������"Ϯ�9�M�M��z5�5����X;2OF!�s�7.>��±��>��I�]2>9R0>�]OB��
%�/٧E�r�gP�>����yv��=}u{���?x��;����}띷~��~��o��' \��������8`�G���Wo���|y�����WK���m����A��s�AM,`e��߶��# ND
� ߳�w�2w?b��Q�v瀄x��~(mK#p��o8Z��h[�[?+�{�$�%�?�D���������<�|�{�z��ӵ��j���e�
_kka���������$�7�I����T^���r:�O7���;�റᮠ��:��Hxǝ�^���#;�P�I�Q��
�=@������
��-�l ���;�����l@�Ve&9z�7x��0�y���ǂ�Z8�$T~�CN}�Iۦ�s +�Ч���`����c>^�����|�c����<�{��<`�j��Wݝ5��`�e�:�����/$`Vc^98ƽ�T8}���$���,��U��  �@��<3�tc�c�� 
G&��`w�8;�G�}�o��r���8����N
�0�<r��z�9���[��hA>]A��e���8`�����9�[��Xo�钌2���׻�sд�x��]T4�[��p�~Z�q
RI�i��G�=�0�:�Ok�^��v�G��Б��?̛}���i�y�5}�54�:� �m�������,�i�<�Ebn�{�nnӃ�?�9�*�,ky�N�y����j��6//�xaԛ�v:��2>u���g<�'P�ѧx�uJ֋����;�4�2F��'�f]��o�Oyr"�]�~�}B��mՑ]���߂�\?�T"��2���,{�Q�~�_&��G�]S�ߣ�?�7�Ɗ����q��i�Sq��G�os?籛�m��l�v{FC��L���ȴ�#���&|�P�c�/'ʡ�V����z@i����u���w"�//����>�.�~M_J��I�U�-�D�9�qRR�=/0�*�q�w��ǫ&�q[���|�B��B'�k�W���$xQ�U�9��5�Y-���Y�ui,Wb|�b/٘.O��.?�CY�F��H~t�
�m�y1�_�4F��Ƒy;�*�f�c��t��@����W־T�?��|��۲��^������5PqLՅ2�ǹw`���;I�Z���B���#���d�#{�F�繚eF�E>�N�\�y<���d��'�cYˢ��rr�ˋZLGԟ�'t�,/����RջG�>ы�Y�r��qD]���uF&�����r���SU�����B�k����S��y\�������������~>��8Gx	�����
����,G�3��.�|`�'����̂���yQ=�����+����*�"��,ؔ�r^���Z������/���	� ��Y�[�.;�����v��Z|m���y�g~\>z�"�>��w�z�IԱc��+S���:�Xjsw���&ۓ�f��;ͫ��)f�����ֻ_�܄lނ��4 ���ps�4����@/��Ih��.�w�~~�>{p~���������?z��g~����O������%�;`h�7�|؆����^5�nw���B�^hDTE�U�_�j���XDCYPj���Ѳ�71;�ǿn�x�C�����L.���u�b�E�Iׯ.~��qpدF�����{(�=�D�����7�(o}�-Y�E>�㏮�^�|Z�	ّ���9ua���_�����
f%}汉1�f5�czr�������;��@u���u�]tAb��|t��H@�3,Q6��!��rh �
���B�Q�2>��Äw1 �Ak̫�m��T8u���d�������Tf>��8�G���i ��9�<�C�e���HN�[.�<�:��y�a�~YBNQ6_U���8��-h��H�9r���A�z�]�.[����0o���؆�q�I���Z�-��e*�0�?d
��}ʺI1��ks"G�����fG%�[���m  ��IDAT��뫲8�z�\�9�	{|o'?�}�C#C�"�p���5�ak��G��F'�6���5�h��ا��;l4���@Y
ƴx�� Yno�ˮєk�`A,(S~���&�y�o�fd�F)㏾��������&NZ eogQ/�lg>������|�z�u���(MAw��T�i�����(0�v���ɟ��H�W֓N��~r�3)�%���>�\O�oa����[���^��2��os�p����:&�DBQ/|��骺H>�����<���иn�_���â�F6e�?<6�ޑ=f�˼b:�Tc���@��ir9����2�2W���N�gg�0�{��-����z��z8�zTŲ�\|��o���ԅ��}��"�L�k|U��z��{��d]0�&�Yb�s�Z�/PUY Ƌ��#=�j}��0�9�)ݒ�<�C���s�w��V��c�1�����IF,/�����ß�&� �n����=���{Ǻ��q�u�V�wTmG�f����E/擎�~�g��g?\�8�>0_G���z	E������xƼ<�1ϼ0���5��!1��IY����y���y�A�Ce+�|��^a����d��}蓰��޸�!���� �m,hg[����6����<����/��)?�C�	m�5H�����_>YBq�&i�o\�'6b,yl�/�,̲Q��3Y�������q��$LX7�:0F'�s$��(�d��[�H<W�8R�S~�ފ�D�|j���f��z�1^�X��X#.c=�;����^_��r�_��l�j\!�	�U�2c�e���~���	�="X?by�#�D��#hl7NP�~،������ �_���o�c�<�4�߰��|a:���i�ھm���o>܏��������������陼X���_��y_ߐ56z4���q�h1|��~�R�w¿ظ�c��?|<J4��9Ħ��J�e���b�H}ۦx��$��Ϯkm��ņF�к�%?�ض������Y�z�-������A��	 �k_�Z���My�O�_Aͳ�1���P`�,
�H� H8ѱ�|��I� �o�؏�r���q�q��0hgP c)��:-���#}����_��q��6�����r��7壯O<�c���$�?zU�����󾼲�r}����-����I��l���H
>� 4?���}�/�1�r�sp�M<�l8����X3=z* ��@����lኌ=g�k?bg+x��;��؁c2n���r�|)�yѾ-\�~W���ǇS���L ~v`�\�{�i��+_��?,�r9�1��?�G�H�m������X����"�I�wD���� 8�TerP8�v'&q"�;����C�����޸�0���C�2?�����Y�z���u�͚u����6�D��G�G8Wu�}^��r|���U��N�^��h��H��p�+���ˍ�����w�]�9�*>.����g�{�7��<n�8۸G�҇�W�p����a�Xa����;Öoq��^_ׅ�j��.!�ps�|l�}_(��� ���r�ą�Ti���N&cѻ'*0#���n^R�JSf�T�~٨�b���]{D�n�O���X2D
_�7?үi'��i���=�t����L����
�͓��&�${-�)֍��eFm�`8h$۵8��|^`��&���V%N�b[����3��T��:+'&I�10�$��w�u���̶�mP�Q?^$�`b,ư�b����v��?Jb:Z�f����4�9����sf}=��uh��x$㤺�4�����v~�����q�|Gx�yu��������ZņYVo-�c���V�/�UV�*�/������B�}�:_f�ݫ�~B��.�8F=�B�1�Q�U�<�xz�錉���D�@�xh�-/^a��!3�'O��u���9��ʛ��M�����������4h�e���^ a��\]-��d܊~���3��K/��q�;�6c���L�������!�����
M�^��9�l��]Ř;<G��X$���!�17j�?�*뺐��(�ʣ��s��8��jOf��S��k^��'U�bn�S�@!��߱���BzTl�I�A��p���u֓�o��u�c��/�qý�A�2t�%��Uz����g}��8e�O�T��˳��|`�2V���&UW2�`ț&Z㺃���Ԥ�j;B�tA֩9>?��l_�>�7\�1w	�;ۄ�yy��b���~>U`�g��gb����8ym�	z��8~��*�OAYN�T��2ϲM'�ɔ,�3MqȬ��o�;o����H'ez�8Oع,��pU�`=���s;�y��w�یw��_17�{G��l�lѺ�M^lg��?�u�3����g����y�\d[0�� ��ݟ��3lq7	�6|������� l^=-�����5d�t�1���� vk*N�R�P����sl��yV�y��1x��6�ƣ��<x�����;�Q�R�ɯ�L�5Y�����䇟 �+������W��{������������K�ڶ>�;U�Q��G��w��pV���j.r�/�m�ߡB�c�JF$��uu<#1 ��rp1@Ú@�.��q���0��O �mm�������H����{��ޑ��}���oʿ��??����@|��c�z@��S��C�O��gP�<��'�H
��S���q�ٹ�:�p��	� 8��9�3����k"ӑ�l�9���2�y�Jԓ����hˁ�<����#�|��1�*t�#���.�g3��d�]�8v4�� ./К�(�F 嘞8d���,g��;
bw=g������*�|��- ����F�0�c8f�+�8bZ���bٿ�c|��b�ܰ{�s��UZk��I����в��ߙa\瀃9�ża�#�� �G�d��w���G���ms�-v����S����>nS���,h�+��5��)�O3�d3y���#�l1�%� t>^��:Ga�d0�wz�l���=��&�u����P0���U:4 ��������췣�ȭ؎%Z����A�+{	�w�eY'�b#;&,����sR��Fre���I��5JB�_�Q�̽�007�e���@��ů%���k+2��*��	�>�M����E2�S[�)����o�o�����ؘ��0�ɲ�t�]�5x��Lo
�&<�������� �����G�ylؾ�1c���8�%~d�w�������#�1~ûÏX��.��E����;p �ڪ�2v�6�w"ׅ�F�e��s����ʟ\o�}Κ֦v�/k�eX1� ����'Ǎm���Q����w�ߌ9�1x���e��_�����JQG�kyAA礩�����3�����s4�rg����n���3M�����/�T�kt�c�~>&�����8&�%��i�>�J����9�_�����]�!#�7`�|p�u�cKlWlR��/��t���Q>��>�0�j7���ј'ۙ� ���]�}{��X�yl�4��s_�����SW�MY���y�B�10�~�n�x����|��2|���)r�r�;���&��]��`�D�:'3�0�$0<x�d�&ZKr�§䡽%��$�18Y:����|�*��@�Y�����<�bc�n����&�a^����m��~t"&�����ݹ�骏�/z��
,����h��5�0�2���x�,�����-Z*�{(]�n+�HF�+&�b�mU�����X�����3��<B��Q���H�G>u�N��[�or4'��Rr��9�R�v���,Cse|�ʻ��ҕϰ��d���:�/�شz���ٕ���3���W�_ޗ׏�������nz�1�z�
�yغIÖ����b��j�}���N:�GiW�ͻ���ܘ��ރ���@҄ͳ�ŵJ砱q~s\GcC^��K����<]^�k�������������Ǘ��������Ϗ�������_����G���_������?�髽�+�m�l/rZס�p�\ ���� .u��! �-.!�w��7���o���>���HC����M8��"�����A��XD��@�v�E�����i;ˣ��#���D��o���?�����o����7���'�c=	$�Gsi�^@�� 8y��WŃ�#�{p�m.{�]�ؖ�|�3�1���ΙWLt��-��o��x
 @B;o�y��c@��E��t�'����J����ى��!�����[�m����r?��|V�n��g�w��%�:o���[����d�t��p�-�x��D{�^����$���yGo�g�_O�KB�5�ɼU�(���d��ܷ�d��g�s6\�v�7���5m�9+5`$47X�@i,xE��/7o�@���4C��v���}:�l���s�y���<�/�euh��@h��n�-v�Sž���z�c��]�8���v�ј�t�m�5�1%R��F�&���c���z�>�¯- ~
��M�^(}j�
ؘ3O����$v�m���T�v �.�q}'�V���wm���9*D>��4=�EY�OjU����d
�,�o���K��Իf�},llq=Ej�:��m��[.}��X��'>H`�[��bf�$D��~�6��;�����lC2�YwW��g|R1}�D2>GyJrP���d};��˞[cU븍���l�����w�RgK~��}wT&��v�ý��S�C��ۭ1үcWn^�z�iWq+F��`���<�$����k��3x�Y�7d|>Ƌ�SxM�'-�
H��m�){�"�pg�t�/溁iX��>m��k�r\'�o�Ⱦ�օ]�G������ѫ��YO!˼�)�v�8A���#�{$�Q�F0�N��|���T��yM�l9�䘐�*��<����߅�wx��������4�c܏dv>Y ���e=�ؚ�!�2��i�	��ݬ�����А���ua+|&�D1���B����<,����M@�m��)��>�'܆�q�z��v��V�?B��M"��d��1��E��o��c�C?��#��}��a�s�)lK�?��S=��*d������e��G�[�v�km���m*�U�<���'y��N*	�y���_�l��e3���@��zƶ@cl�����}�?��:�I6G����qE��@o}�(A	>(l|����D������$�q9��>o@��;3�d`�e$��_�o~\��rsz��w������C��5�����u��_�W��מ��?ٳ�������r|�^H_�V,��;����Y��Q����V�����9We����=&5� \�m���z� �N��6i�#���3��
v2��C�o��6�(���ݳӋ��?���o<|���e���W_}"/3����s��?�CN �*��+����tY~����������s[��P϶�@�(�3 f%;Y�Z�|�TE�;�����) N���JƠ����F]�������f�q��2-v�����Q��W`sm�鵿�~�Uy��S���[��ܯȏ?}&Ϟ_��S=�~��w��j���`�i� +���l���pQŌ�,��v���΃V�Y�|�A:��&P$��3�C�zq��D���ӌEN���ZG�m̶���M��������wGgp��)��* �k��l1\s��FG�X��x�w[�'�x�Tb>1�:+�~�\�Q�y,�� @�1h�u��4��/t���g~�Y�����t��h�Duv��@�Y%�i�> ���o�,9G�g�c^��ώg��l�r|�
խ��U%([u��jN�}�F}����7�-,���������C1o/��Ω��yЉ慟Z����3W��q��Ŏ��ߛ���^��uqg
��=��r��4���8���6�o��x�_`���K�Y�Ϯ����4����+!�k}d�5�^6��^Z%%��ƽq>��.���F\��Wu�̏2[8����˫xAV]���xL�r�m����9�MG��6ʸ(w!R�}x���t��� ��v_Y��7�x�$�L}c��A�.����/���[�
;�@�,\��0��r(���z׎�=��m{��Y����aWPqOv�!,��$A�l$N ��\['[ie88�]�+��T���1�������`sm�["�x��9�o����`��9����o,�$ygai�d��"�)�;�x7�.�Y3�N@��p�����d'ޏ��pjn���v�仳���y��u�(������(�[��c�<+�F�K�P�}�s��h3a�EW�-� ���G�z�%)v	�ں�"2��؜����NL�%��PZP7N �9���e����4oZc^ŷ��!T�_նbn��Nc�e�����.-�we�dIm��h�W\p�.��L� Y��l�HF[�b�Cہݽl`�L5������v%;�/����I(3��ق>ֈ�{��^��^������u�q��׆Ѭ5p��1����I�mW��8`�v���3���b�X�v!��'��ak���uQ(����`��N��/��1���`I��4,�#�"��{�����C�K\��c�Ř��I��)V� 9��9q3x�k�Ȅ�~�.U^�����C�oB�waL�t$_��K������]���:�I�^�oҗ�v���G�����H^�.�t:(P򻛤n�k/��e��M�0���~�9�6M�Nrk{�y1���a�t��D�1a���7A_!]��K����G�s���Fɒǹ�⇍�'���q�l���Z&�-�R���e��bAR��D�y�����>i��c�6Y�����*��c��e},���N�[���Xg���2��׀�ϝ�<ʲ�s����O��Md
�H8>q��Q�ස�Nr�DE����̰��m�jk_O�,����F$�c��\�O��Q�/<�����I�u��t��d��Q���D5��w1}
�!_5::���'��&	}�y��d+̶�M�1vrG>����x��/L�4O!���5���\��^���۟��_���O����}z-~�������>��Q�  o����'O�|��+�|�j��صݛ4]7 ��N��+��=�h'�dN�ş�;-!� ,�N��(#jR�pI�3+r:��7���ی��T! �x#v�����WG��ۓ�\~��l��������_�)y��#����H"p��`�`#��t�X\�}���&`L��0|~gsϿ;0ΝƯ��� OC�*4��l4-`oY��������)�ßy֟�>� �p��0�y��;i���"(�|țQ�d��O�bS���� Av�QD!�ㅿ[}mv��MYie������?	;,\&��&^������"���~懸���$�I6��>���|�b=�S��b�	s�r�I0AW������x�l�;��C�m.K�/oõx�ym��`{����y�^�Qd�6���0�g�]ڱ�zχ����DV/t�:���h!��I'�t��# K2���������b�A�0�`/��c�f�e��E���k��b�U4���z��^��4�����:^'�7O�Z,Ѓ�."�A�C�`����Q"i�]/����'����Y����6��m�0p�b|�CT�� ��B��<�$
A��d�
�:�`����@7�=]��_�R�H��D�Œh�'���(߳_l�b����_���̾3�7>R�`3+��_Nӊ����J��疨�XE^�qy!��@����7�.�g��i���=�n���՟n���X��8⏨��Knc�zݕP�>v��͏7�j�[�ǋ�$�5M�iPu�����=�)XT�4�\�f�j�g���Ǯ�%��Z|���&�Irӽ��������ǿQ_�#�N�@=�7���~^��#������!�M��ń��Lk�o����LAw\��h'����6�m|ᾜ�"�����#���A�0S"�}��hQJ�E�ѻ���O���>�vN���g��si>����d�ޤ��b8F��cC�P�<3�W_�[�cK,N��@>�����y'y�c�m� l#�,�Ki�&��qr��G��Gu⭕i��Im;�"�@OJ�J#I�Q�xW�߱y���c<MEb'���d��E[�6!?�?&��4O��H�ޕX�� c6��Øױ8b�B����I����m�g�װU��c��&����vBdفߦ�u��i���.u�΋66�c�}l��_�'�i��2��k�l�6�tŇ�EM��b���:��5��E_���z����N�]:��r���d�d�����!��k�v�l���;��b���#ĺ�S/��Ɛz����67��X&Q�˙�T ��u=h��Q���B�徃�v���'��������E��۲Mq�{?c������vNt�z�VƧȈ�S�3Nv��C<��W�o���S��0�<�t0-�^����ИDs�@�W�8zj����<�Q���}�W�k���mؼ�u�N�3Z�[��H;�E�+�H�٥��2�es��f#����}���[O�$�z��[a�[�����B惿o
7��d���o	}�'�H#�_��Aw}��Qq��6�=��SW��_}W���_����?yt����2��tv�6��5�c�V�S�ߝ	��}t��,{��\J�q|�U��-�����~�Oև�p���:W>d�w�'|
���uٌӚ���<�������O�i}O����vB@$���s��?���$ | �O�����?z�Iqz�/m;_���������O�^�]ȍ:���%\F�k�^b8�n<[?ِ�`0-�i�m�ҪA��-��	��s �U�i��(>�����;�x{&�������]���������MH8F���E�}1�}GL&� ��r�@�j�:�a�%L|O����� R�m���ae--���Ǿ�0�}q� m<�;�5f�}��3e��� �2'B��*�C3S�}����Y���ü���pقP��.A�D/�d���8f��r����(�Xׅt����|�	\o}*�,��@�����K��
d�B-���R�Z����݁��ăf�n3�6����^v����[zd�Ñ�m�"��J�Ώ���|Q��G�x����3����KRD�@s�5���V�IX�ku��:��^������n���ӝ��z�wl��W4�J>�O�Y)p�Ҝ�Pt�%dk��U�D�cC#i,Vo�r�
^�(��`���sX�=�1XA�{q�u�+&���ve}��bQ	g���#�:� j�vܥ��I,�-��l�F��e�CA���/Q�/�GmL�N��/֨�k.�ɵ�b�e+p�����f��}Li땘<�w7+�.�q2 t$��d!�(�ĮO����AztY����Y|G���v�K,��$�� PƱV)x�0&i>�8���^�k�X濯ȷ6S�K� ��n�o-�|����SW�ic@������Xk1'Ku]�QC�	M����5���r>.�l��c�ΈCb�}ƫ�;k���V8
�F�5���h��]c®�6CO�6���/�N<
����}:�9/ߧ�V�[�z��U�������m>(�y?��yf_����n�[������^[����.�P���OH���c���y�Mݰ�60�X/o��>uN*t�G�����.�����l#�������%p�/��ٿ�B��1���5a,�a�zg�O�ӾS|�4�Nr[^��Sp��Ԯ2fu�G�%�.���
�'�+_��(qc �1b�Pi�{��T%'&d�Ƽ����M�8wg�����v #��Iӡ/ݎ�Bkgik�)��6T��WY@Y����z��_I�x	�%������)1[�bD<�/���%CS2��>4�,�P�*���Փ��&�dz���|R��7p�*z,���hv_���]6�֣g�6�z=�����N�60>��1�"_;����6�XFz2�@�C"�a��5���-�=�;-�Up~������H�ŤcA'=�}����Hk-�K�i���J$[T��[\�H�/���c���n�5��K�x�ْކ�j�_����r�wrgr�����	�6��ۙ��v�g�|�e����[q2A�nS��tois�R��kn�ukMe��?���������L$�V�AL�E�[X<_�D���?���s�u~D#�	䭥~:<Ϭ������t��:��k�ׇw����[���^[�E��U��'��A��������u
d��*"{�6@�?��8	>G��D��N�A���u<���A��K�˰A�ِ�욊���Q8)�;{4�f�<��&O//N�����E^��Ń���R%���s��?���$ ��wZ��飿���7�?^�=|�.˃�S{��	p;@t���/�"�G�V`$�=��9@�0�v�#�B�G@������Ֆv�T:��^���� �}�[>R[�z7ݶ`�� �r�ɋ+?Oo^�y���y���x�^lr��^A8h�'gx?&/���Q>�X�����Д�JM�������`�!�ᵹq7� 0���2�-XMc���ù������F�j���i oMp\_����n���N�.�wH8�|:[T�?p҈8��^��{ k�{�Y:�M�I��A��h�HԨ�i(V���A@`O�Ի����Nm��N�儅1O}w{p�H��s��I��w���+�`nu��ɭw��:$&|QWtGM�9��]\Zn���Z�rcv:��>�.쀅�w�^T$�]�kő�8���v���{��,���k����#?�r-�ۭ���YfH9�ϓ.��T�q1���H~�۪��g\�U=�Gڊ���ee�-��|G���Ny�����^��T�	�mzr/�p�����������v�^���:���C��:l���1����=�A��.3㷫�l�ݽ�.M��v������֛�9t���w�_%YO�gbj��gq�K;��ܰs�މ�sH��EC��h��q_-���i����7N�ۙH��]@�t}WHwZ�`��c^(O��t�k�t��b��r���_?�����]6�P����j_�����k�����lG�U���o51�a`0�u�2���1��<0����3N�0�@I���o��@�_V���\�y�Nn��2�b<�b�c{2�Xx��=u��G���0�[�c��9��]���>�Eu������D���-b<�n	 ��c3j0s����5B��9��x���(��ʾ�[3������|bc�>�#|�>�b��O�ĮP��������|��d ��+�'��S҉D遗".���7ē=��9��n}Hw�{��{�c�����K��2O���^��+1���h��+9|�J_���=��㰴ܯ�PՑ(������6�Ls���7�o.{��b�I2~�*v�7ko������]7���2x�b��c98-%��Ƹ���.t�"��~U�&|$�_�A4�.�'�1�u�r�����byg�����|�E�ۅl�^l5����j��H?�d�ci���Y��l<�Z����C.:���D�s	>��Mss%{�zfM�@;Z��봄�����,h��o�=Q��ʘ��Y��ݝ���l���Q_���V�ۗm��},�F���Z��Z��}����Hz��6F!�8	�����?˦�{ԗ�St���5�����1�n�%�b1q���}���}s��ǼC����lI	�]X�ɺ�4:O|��ck�_e��������m���j������^l>^k�w�u>� �8e�t�f��g�{66	zN,^�|m�l�R�:R�n��q�Q$/HG�	���p�����7�=t���1&�yA|�xc2ϛ/�.�)�3 �h�u ��o����4�>9��<B�:wq%B�����V��Y�NsI���)D5i�ƉY��I�[��m���Э��s/�r\���1�/<���N~���7���s9���Q�hy�<���b}@/��_R=�@���8q�7v�$�6y��Uy��#�g��P�<�ȧ���ݢ	\�����]l]��<1�6�qh`K���������D�c�x��;"�$?�''ՙ�Қi	�� �3(v0�(����o��<i��W�o��������{���^�ȼ����9x~�	 ]�w;?8?�/��_���y������˛��קϟ4y�D&����Ď�8(��`��F�[3E�@��3�2��H,� c�� ��9�ҝ���@O���2��؉h���%�$�&�w�\.v�� u,�]���p��p~�$=}&����ލ�_��DG����|��Y}[_���8�"��rp���/��ã��G� �:�|6;{,#�i�I�1��C�(�h�����`Z�<�p��� ���z �e��� ���k��7���>���!�}|������uu���R�́��=_g ��ߝ�An�(�}��(�Ծ���黐|����N����4�_����˱�$�1���,`q��q�?S��Ա]�/���{`"tV~x^����=p�tZ��� �^��`��N�b~B�/W�x��|w������q{��[G�*�8�w�l
nnqT(�sR����G�-t�˦�	Y�<�1~W��%�@<�������;��4�r�
;w+%C��}䄳������=�w����ٝSJ�`�Ag>xpJ��1@p��GP@��ݺ����^�+׻��B�u���XX�N��ao�����hQ2wz'�b��F�	
c^�cbN+���� 9ñ�Mt��k��w�["���1���9o�&R���.�f�/<vK����,|���^��{��N5�_���?��
v�bn�\�����5�VvZ�D���}<O�޽*���kƇ����o��<��Z�b�k�u�q�ڝw>���E�Wkg@�]�����-B��$�qҨֹ�p����B��FD�>�����4����M����YZ�Ӡu岡�8��r�ZЃ���r��&A�Nڶx�'1��{��a�V���g��yO�%��y��T��-��/x�34�-�M��*c��e�&�/t�S�0�G�h���^`�(ρ�H.U\U�$pt��jhay���2S�����>pY�x�a�T����Z�mY�8�}����Y�9�ǵ4����>to��^��r�/������h���<coK��7���m��"��-�\h�5t|-�<;9V	�g�:�xV�K���v���߁��+~#�k	w�<YƷmI�O:��a���>�k<���e:v�^����Q�G�����|�#y6����+WW�n�i�������]m�y�����Ӝ`���,YG����|�+/����Yc(��6��� ��^n>����c�������t��Fw�.c��8�R��U���/���}O\�vw|���6+?Ow��з��1&��#Ip��c�����vd��y����q	��E�'-!��)���IM,�P$��۱t����;�c,X��Oɯ�5>���8�\}������׼҄vQv����"�[���z[�(pv���S�ٔGЃ��!��U�oa)�� g��!9H�ޚ��WD�g������W耰��u�>T�7ǝ"q��a�<c�~�7�ٰmn�q���1�t�Qۼ�:�S�D��̧�&�m�I���l�	VC����g-��k��Lw���5!A��e,-l�|�cv���߬��	;	~�GO�h�]Ǧ��ws�9_�m-I�p�%6�HyX�E,\e:�g�1�/�x�2(c��ґ<h��j�n���wߐ��'�s��t,<��Z�yӓKF�Y__�Nv�)�F	L�[�q�3š�|F<�ǟ�`$�4y��C�F���䉩I�z�b>�I����*��K��[L41={�7gT�����<z���?��������_�����۶�~}v�~�p��?����Gq@����跿�{��7�?������e�'= Z�l���=�
�b�F��^�߻��}(m5 y�r��.�uJ�W���C��!�N6��/;��<t�����ы��������:xX6y��j�޾~~��2��#�Ǳ�z�[�X*T��&nXz@��m �O�/|r�>#@Z�V_�	f�_\t����n��e7�]�F���v��3|��`���V ��{��] 0�Φ#�4�I+��Ƿa�'���E�XLfG��� 8n��N�[NH�qI�.��5͎]����fs爖��ߔ�`GM��yACn_�oV�3F����>
��Qw��7-��6������qۓ�:dR�����eӝ�FA�� ��Ülc@x�
��E�+ߑ����b(R:�6\=~��9���Y#uA�ٝ�2����dp|��n�//��{��P��qG;����=���'���-�+�t\�$��N���U�O_!�$C�_w����-ڑf�S�w��9#��lw����c�����1~4&j�1	g��v+�r��$�G$�@v�[���2=����{]�@��c�u19�eF����c�u'����`ug��G``�u�ރ`E��|���c�;Q-h�s_aX�aG�����������m�1��������.n7�3��ݝ������ی���;�a�����t5.� �7�u�Б������Sծ���r�ͺD���%�H��F�k�#�{�7?#�`�|(���UƮ_���G�WŎ�b��-�,#�4_�X�i7��J� t���:u�Ê���������Q��d�P���1E���3��1�1}��I#�#nAv�[�NȊ ����M�@k��J���HR�����`$p$��1D��"%�+Eٿ��U�g�'c���ٟʼ	Zlt\�v�;|�����	?*#�K������^AW�b-�7�%�ӟ���H$z��b1{�I���qh��䞇�d6����JZ��|Ȃ���A̗��|!L�]���B@�-JPn���O5��Yv� S�aӮ�.�����]Bgm��%����'Wypw�B#��0Ps�rMmc�11��co>����'�x�Og�������l�ONhN%�b7�Lћ_O��J1�e������N��k$�����d�ԨKl^��.��E����Ĝ��IB1�F6
8'���Y/�1��|ȍ���Zr���O�
Ɋ���g��k �Gҏ�#��6	�v;ݚ��2X�_}we�PKsG��z5|ei��I�����	�>zBϲ�x������O�t�K�M�#���� l��y�B��@����w�-����b���&�����>�y!a�7K��IK���Ft���|l"���qeSo�n7�n?�,%����c��������<rq
��xԟx��vTw�}�O��|7�W|�h�v<�'Gle��NpOu�i�"k��&P�:���7�R�e,��g����F/���([cx�7��1r���q8��� 6�0��zZg�y=|s�8
�+}'��R�-��'>	��W��1D]|�Ю�F��1M�A�%�o��Y�t��6eus��e�O�/�{�XY��$�bs�j�7ۅ�;!���k�)6AH� �ʰ��`�~B��ih�	-�s���^�H8�r���8!#��&�Ի�)ch˝@��D�|�W��c���mO�8A�dR^�u�O�*�\�������z����TT�#h�%���8���)ؗ!�K��a_î���_��'��I.uJ�`�^�nj9ۈ�B���]�_*Zh?p�yb�eBr����	��*�h�����+������7��[��o��W������O��?o���?���s���H X~�[_�{�<��<t����U[��`��Zʦ�X8��"1�_he�G�5�Jia����������Wܰ���*vh�.ּk���#S��w3�<�-h��^����-���>ퟯx}�jt_������A��Q8o[�a���M��A�u�ܔdQ��j��:�y7�k��N��98�w�p.��&Ծ�i��Ƭ.�ᣡ� �������iGM��̯����v��f��,7rp-�<9�P�I'���|?Y�a�/�.����g�RY��xW0�h��>;/�Ct�·�`����h��I������u��"�9;�;�G�g�E�	2��G���C�����)c��X0�cR�o8�p�.����s��v^/�䌿߿�}���uq�p�^�D�:Q�'��o�C��g$�;)bN�Lw��q��Bৼ�E�юi�9
��{�?7�M.x_/Q� �:�#d�?�^mh��Y�(t�B7�]��#~o�����,ڏ��T��ܻ'4[$|_[S��@�i���Ӆv�وx@g���p�6+!Gn<��s_��G?�i���L#�z�+�&;�I�fg��wϩw��7�C��N=���+7(��z�<��;�Ŏz���7�*.]��%�\%���Q���,&��v?���p���QG#����Xp7۴���w���S����mg�3yӺE��[Ý�}���ee�@<����C�w�ݓԻn�/��%,h��#�&.��#"��h���Ni���$k:���X�dD��f�[�~��Zr������x,@?WJN��1��C����xP�:���n�A��m��Ⲵ5t'P��]���l�wL�؃>QN�a%�Z-du,�,.)]&]���� ����B��_,�:<�W�V\��w#{ X��Hތ��WO�A���Td��&�~|�&Lq�Әw�����K�p��w-��1����mо���8Į�q��?�E+� ~����K�/Tu9�)'zF�Smm�,Zx�!���l�^���JA`6`��i��O;�V����td�)��r�9�h����i5��y৊D�a������za�;N�3��	���ZO����%Ͷ���	0���o���}aWR��l	�5$���c��5�/��s��a.t�'�'�A~����d4Ģ��X��Z��$T���qĬ���I���?�^��,��k��(>�1J��%�?�7�\�~�Ӑ}[�&:����W�NU����Bov2�O�'/\o=v���8�-t�;�,Vz]Du�Jǻ9����&�|g� �܋y����2vS���ol���k,f��
��_ �%�U���9�F�|��Ʀ,~$�vQ;�����9�~��h�Oq�1�r�Y�GLO>�\R:��y��4��z}��d�5p������>F��sm��U���� ?z�`o���`��ڥ��f@�����<�#ց1\���و�vX�6�C0��ؙ�Qw<t��K�sNc��֐�_6����pU��푸f�:����~ޘ�1#�.�-Ie����bn�[c[|��gŊ�o��cbuG�>9�e��Is�O2�ej�lI�cl�	�81o�S<�Vl�H�����De
�`��K$ь��%�4_;-Oы�vW��1���}�}ج�r`���d#��g�䍾0��8�f6z,�Z�V{��R�2:M�� C��>�ڂ��uhg��G��M<�>t�N�C�o��=��� �Lp���>�ˋ;є�8}mW"[3�H:3p=�VF��px��� H:�pi�!�����>c=���Ir�׵�ez��I2¢H:MX��ƹ_"�&{�Ꙭ����]+}��d9߽���w�=?�<<������Ǟv��`�������w�<|����a��r��Oq�g�������6��eIzP���9��|Y�YU]��ݭ��e	a�@l�{Ĉ)c$�	H$O�y`D#����@H �Q�E,�e�iWwuu�dfe�w�9{��^����2+WI���^�{����'V���T�me(T&�����V�wi�(��<R|�����9Fqf����,@!f�ЀO�Q>� ��/� 7 P����٠��>��ZN��͸�]v�q��;�45 �a��3� g@I\9Kƹ���뽿�z%�GRv����?���I9*�#��/ �!Ï��8�4b��X��p<dŞF����w0�~��s�P�� ��[i���7���372���>� ;ّ�Ȉ�{��Pr�7���?s4T��L)X�;��cOY-��#���2��^��!�E` ��WJ<�@���2�ٞ�c��5{�π=�3�K?�qރ�/�(��&�G��fo��,JH�kA`����?�co��}l���g�B�	ܷ6�W>����O�0<DU���o�,���r-e��a`kp�&c"���>�I�5RV{&��s'� >�?��i-¸��NFx��.1��dx��0L��\�}�]ZTٿҷd�����u��b��ʗ˽��!�;�CL�UܒC��F��Z��s*,����~�S��Zr��`\`�4���m�\���4����#�B�I��3�^/*�4`7��_��ú�R�!;�!�:{��;�ml9rm`AFٌ��U'�����(��D��)��j����:܋������A	���H�K��p7�h�޿�,C���O)֘gy���^�6o�F]��}yK��G3�1i��G�x>3z���R�6,a�4½��K��0#Ui�>�2Թ(o	����g1?�i�`����m��mZ!���;��������*��� ��!D�8~�� k�d	�a|�a�r�\w\h��gQ:o1��:�(����(������bs��g�0`������S*��N\���&�UF�_�$������
�!aB���#9s��������r��E8�:,A�Of#����8V��K8�X��QItt��n�-�:ݖ�Η}�&0x���m�M�e��;u$���	�9���x
t�Qq�G���� 훌��_hKS��������6��.<n2�3�'�f��5�(8:2o8u�-A�6$ĉ0f:=�w&�q����z���ˬw����9h'�|�Ñ��y�@(o-Sī�P�P��cb�]�������y��.0�C��d���=a�R�^�	�{��}�v}:�F9j�u���_�=�.[,S�����<�vK��s=�������,)��֓�T��9�
<+���쒪H��-�@s&K8��x0����D�c���9xt��u�z�0�u	��v�U�:�gMwdb	TЪ%��Q�΂^�*��-Kg�a@�D�b'!�k���-����z1'���y�vG��2�a:��Y���K��-�ݫcx]������L�,%YV�� �Jm&����w�^=���x��r�d%�N�5鐥Ȁ5�;�P�̃V�Ϟ��jg�'<F,�����\�:?�q.)[gŌk7�?�(��^׺�+���s����`����|�����eņh+/����$��up,V`8�o��F<��i����x����{��H+�w��;8�*�7z0�q/K�TL't��H�/
X��.���%2�ȸ�����'�['n��)�E~�=c��c����n_{
�9ܾ��q�bɧp߭>���?u����6�c+7�aq��I-���'���l')���i���vvr��nI�(��ϱz��Ed��F���W��F:����E�-��n��3<y�U����8���Ħ�O8�v<�Q�"˔O�}-���g\"���O{8�I�8�gG{,����f��gO�������Y����K��O�l=aFB�{�<�E�
MG]�H�l�����y6��Sco�F�5��ēψ'8�K|'�`�Kq?�7l�x.F-��A��wv<X��Q��o,��d-�B��z����˯�t �r�_��~q���{����o���)2d�r�TNTY���\d�$�L��x�IsͥDɼsߪ[3�hB�� F��φWdO.RD�`��c�2h�ح���6 d� ZdO���4�_���gr�����ң�V�<�������(�$�@'5������87І�C�N��S�s��ؗ����?���r�� U�8?�,�$�i?
ҰR�٤$yg[I����`�O�6��i)�8]�]k� �Yޭ�Qf�}�^8���b����w�y���Ur���I�#+*Y)�9��ww/�>��1�ر|Y8]n�>*����sI��~�N�a=��mPKk��-�9�CDN��0��Ʈ(���[�~�s<�F��D2
��
J��^��\��l�=$����9��9�F�Gor�'f��lb�]C1�q���J�\�c�,���N����Z�6��L����4*Lc�<+�,J)F�QPeI?�n��!�.j�X��p6/U)�l-�׃�u�6���ge��L���J��j�zqey��eIQ��X�.L��y=��v����|�Af�K�be��N���I6�:����`f�	"E�u0�����y�t��í2J�������^��)���c���lo���t'�.��a�T>I3��H�]��B��wA�@:��j�cYc��]se.�n+I�5��"f�j����Y@�IOD2J�A0ž�"
����k�S�N�o�Z�i�H2�`5���0Η�~�z�y.!̱�+�?�_�>��se���H�4$�����y��I; ������*Q��!��5|�Q�֝��06M�oN��i,8J.�
�Q5��g�o��7���<bNH�2�ɸ�!K�y⬍�89�t�1c��f�{+��
�A'h��<@05P��`M��Y�R��Y �>e�Mk'��	Z��	�8'B�)�7"#��M� �"Ͼϧ��k������v֤�u����f eH�m��t���y����(=\��<e��Gn�a��M����G}�1v��8o��J�r�n����I���A����L�����^��'��1���[�۷h��1	�C��N�$3�[��0y̙���S�WB��œ�i��f����d�A'�k�D�_1�S,8��ط���&"~������>̡�;�c�v���}�cC23�Lg��i-�Y�X,�P�<�]V1ہ���8��ڍ����-���9E]��b�`�9�[�,[I�O붵����K�vH���vN|����ʀN~�[61���?*C�^̀���ddS�Y�E�ƈgr5�j,�Ҍ��=�ɯ������{-9��(O%�R.�gw�5q�V/� �Z8G&f�uǚ�~R7p��u�n{O�1]�8K+tB�#ճEP�}U<�P�K��1��^C�����̯dD����ƞԃ�ժk��@������R�-�8�a� ?d��e�q�N�r�rn^�M��������u��k�f��V~2C�W���<�e$��N{:�F�1�l'�Rd�Ft�h�j=gG^��Db�fm�x&)���l���Ni�v��,����<�����(��"!sI�c0�AI��xZ��z��5�g�w��a<�$�i"��=㖘xO�٠�4��9�=J�G5L�����쥨.�s�������8�)U���u8#�?J �S����-��}_���S���l���A��s��俟��	�N�g�5q7mwԡ��ߎ����f}�����6#Հ����ҡn�8�:�3£���Py�:���*��� wؖ����*�'B׹]w_k���I����%�Ε�� טT��dcq?B���sY<h���L�}�����**��W7a%�e��-���6�y�VR�ay�z���+r����+���m���� ��2�y�H�?G;��&�}R��+I�`�Aa��R��O���7��P�~;�5Cg���ά��o���K?�G/�^���t:MCY/������������`,�W����S������|��ʵ|��mJ�~ECq���U�(�P` ��, a��Ư��	�e�B�T���"��WQ,�~۟ݳs�(��00��(8
i���)�X�e�]#S���~�}骸LQ��'���A>~� �1�hx�������
���P⊗���ѹ��@G�(���Ʌc�{po|o���b�/B�c/"��G�>����`dㄌ'�&���^`�`$sA_G�ԥ�g��@'�o
�pU�a_a��f̘��������t�w�/����//�=�efR_��_�v��ɓ <n��؏4����\�i,�hl#`!Mn[ݢd��ΚD)у2U���Nq:Pm�~�H/�� ��q�$�2q�ol��k�l-��w �)k??`U,���)ü7�,���5�)��۽�k� P�9<5C�z��,�v��ayf���~~��^�T��?Q�ކ�'f1S~1{D�r�����GE�Va�[e�o��Z�wO���,�}��H޳t�Q�͔}�r����A��-��~f�bIxN�N��Dl��cu����EE���`�8���Rka%-�J�ީ��X����cS^Q��a�:WC?�_86��L1*e�!��K�|0�ݍ����1�u`�X��RX��(�$))���������,z6` ���q�c����{��A%ο{����#�G�7��<����܊
-O]_;�xU�m�|�C1]�5vV������<P#����D���7fo�	�� Th�������Y�ĺ�|�l�3E*��#�|���$p��Y�a�փ��v��A�u-|�buDm�Z�j�>th��Tθ�\܉�����7-�QD��0��uw��a��(@#���3,�z�$�*�ޫu���YT��uo^�;K0M]��yN��l�u�����0,g���W=жw`��������Q6�\�2�V}O��e
X�M����i>^Av�g��L)֥�Y��"�?� F-shnB����� '"�`b����y�
�=�~����y�U^�/���N�}���cyt8h���6���;���ʗKd,p̴�_�EJ���+��ndϘ��.��|/����l�`9�#�O6Fw|6�algck�20��f�����f��Y�Ǭ����6m�5}{VT�qU<2;+X���4�<<�g�]����<���}f2�j_�b�>��gU��h�y���y��l"��O�d����4XPe���r��3Ur���i�sZq_��5h�LΦ!(D�p��3x�|��Bv8�`�q��"|M��,��9��$z���>����A:Y�%�΁G̦; c@S��u�w\g����tN:R�e��� ����"�pDo�E<Z�Au�4\#.����e�$�;��t��� �����m�msݗ�+�-�P��瞁\: -�<U�8���2U{w�����+�7�V=�fY��1u�� (8a|�4��V���s�&P+�[��Nؒ~|O���Ǩ���@>#�g��#�����)��j`�m�h�X�+�I�4#�>R��09�!����J�+��q�k+�c�Op�����z��?���H<O��<g�߃g��d�� -���>�X2p���f�1w�C��	فE	Py�˟�����J�lB�-&��Y�N�)�k��q��spf�?�h�m]�ziO��|���2aH�fmb�6\Ǥ��;�Ol%�wt��������w�<`f�X�r?֚��D�hS�<2��O��g���6�.�+��j��������G̨���H��WG��L���w�j��2�G��=e�����s6{��o�����JL����c���@�9��=pV-Q��fKٴh��<���>�K��]_��7��g��rZ���YGł���h&m-A�f�X�o�����S�ƛ:�W��*��4G�EZ�A�~ʇ��}hI� ��rt��<�t,�˄�-&�D`�O���rH�HB~n�Hr���n��CՎ���r�vX����ߥ�K@:�t8S���65F�w}"���W���gV����/�Gn����ג�#�9�L>����u�[�!�t����G��ׇ�K��_�A�R"��u-`m���"�
d��?���<�����T�������}���׾��ʿ�Oޯk�t�+^���m�|=_����9�O# ��{:��'����}뻿�[���_|s���z��@3`Ώ#^�į4��B*��;9E����������\�`� ŕ�\��ei��%2�z�=��9 ed5��Cʲ�ƾ+0���C�����3�-���ߗ��U�SFm��lfB;�t��.�'�U|Fy����ˏ3C��Tm�|����dԽ�1�Piu�V���� �����Ѕ)�E�3?}�Q���cI��rb���l�q�1J��N��H�#��R̰L��=U��e�-���e��o�t]�����W�������g߽V�j�'��z"�%��P��L��?� 2SR���pv�A�XSb� (���l%;����ZJ�U�]s�U7n3��&�?f^B�N
�bS�X�:+�^��ep<�΂���׏g���sH� B\��4B_���|���?�����v/ץ��'+��l)�J�n$H���|Ń����h҅���"B�v~v�e���R��k޻!ˈ�J�U!���m�@��hBy^���KZ��`Y��h�K]��:`�[+��|��9��A��.��U�RA1@�l���	�Ƞ��Oe��YT�X^vX�XM�3NK8�B	�1���{:�������<W|iIs�/N������L\�����+�h4�57����J����)Ep��I�D�у��b~�&B�y�N	^6_����Y��� [*�� =�|1�7���L���PS��DǙ�z4��0H�C�S��AAs�O����YU<WdJfُ���Z)�ęLi��Wuy�����,�]� ק,m.�G��+:�E@Ȝ�ַ��1�J,ga�F�1Ȭ�\n{��W����f R
C���f������9vSl�����R�-��a482����%2	:�>�N�y]l�lhg@��F��-�Ȏ����-�`�QR�+���Kr
Y+JA�Z��.]%��Ý�j?aH�ɚ��9�9e>m�'c�2�֔�bd(>�kx7�k3�AY�� _�mE�0��{�3�X����j@y4�{;1�d,�zI+W-�o�}3��ӋԶ�{/>�?�������{㴮�vRlq�&]<���\�J�aPLA�Nc�.5Ϟ����y^|f���IH��D���<`�b秵�юm���ӯ��a�n�\^��-�⩪��}��Z���g�N�ƞ��1׬��~�?��m��ꕮm[�Z	b�a�����;�z��h?y7֯#���:�ЁL�IΌ丄�0gOq����(�Hbk�|����6�eC����g����S�xQh�������Tf��B��7�b���7��DOkI���~b��eW[�"q�-4��f�r��<�,\��\Y���͠<���U�]�S�i9�6O����gsVP']o��� <����K"D�,���a�zk~2tʣ^�^I<ԃ�?�(ձ6���Z����?�"�	g8��|��6�)�G2�*�F)���{wy��U"8%cm괊�x/�#V<�HB�p͗s5>���@e��b�Yr�4�=/�
��P�o��bm���Q��?�*�9	9o�x�]ˊF{f���=���>@���M�����<�?yϢ:P�^�6�]�ؖg���?�o�c`��!)h �N�Jb+���:mz�8=;�تiъ����:I�����`N�G�SAr�9������7{�A�%Ə5Հ8BY!����8ǰA�'-ٙ��cO�~�pڃS�:r�5���3��8Z�`��ebѓ�r/�t<�ÿ���yy��;���+Wh��A���f���]$�'^�����p�]\6���H��4���v'��ޒ�Ԗl�ރ���-'��>R򖿏$'꼝��5%�np�����[���Y�&d�����<0��Y��Ӷ��ܷZ)i�׋<��˿������_���s�B��ֻ�Yu��@P�����e�#�"J4�nBY�����Q�D׍zDR��0pΦ�S��d�xd�9�ձ�1��l=��_yo�#I?��2�F��.o�2�����=l�i|eo��_�I��9�;��YIGy���U['jp��IS��4^�/斯�>O]"�$����k$�����th����̕�u(%��/������<�b�̞���Q(d�nv	l�7���������/��?��׾���N�|��ūy��=_����|��' 0���q].��U�~�O��������~�y�?��ŕ|ɍ�G5 :Ȩ�P17 �\�QߊA
:l(��C)�}�lFT��m���]�r1Y����Z(L&�87
*g,�W�Ɋ3�9�X6 ,�y^��]F�f,yX���\�I��@��5�ȼ�9�Sd⢏��������p�T�'�m��C��`F�C��5�W_n��*(4���lܸ�@7�a�S����3�k�2���� ��h�EN���K�Xߪ��-�8K/;�=�ܽx!�����x�z����n}}Z��\N���SZGz�<��3��<%�5)6E~��@Ge�-��S�¡0�op�o~o��5��bR*��?G�)�6�<θ�dHf��-�7D������*IU>�:Ӹm,L(�- p����P��?���o~�o�$���\�ai�Rf��[;S�lٛ��#2�WL7=W/���<a?�kj��Lw�#c���n��E�yt�3S�=ඪ,K�.3��e6��1�����L7���!.P~+[D0��N6L
�;����=V�!���韶�Y�a(J�թ$NgBk�NEH�pn����A�{
+�i�W�.,rp^��c,��L��0e�O�?{X.Z�q8��%O^�J�X��t�b�`9�a��«��^���N>���"�9+��̼X@�Uf�1�� ���ӝ�����w	�?	cK��:C^�`r�01�M`���~a�-��hߍ�	��4 ����1�1v��=àoF���}p�$�5����tF #���&�w�I��p�F�eD�X���}*+�:珪0�4��9ޔ���^�k�̼T��x�	ϲ�v���l\+���?��q(�2�bJ�9v	x��e����s�[�Ť�1�`Z�E�*�I�h�ɭ�:�ƑWd/��v8�!�)�e~jM�N��U#��iY�dʵ�`��	*�F5u@�`�{���(�;�&6�6��z���w_�;�J~�k�8�����A�ݸ;��~�&Rn���ʲ>���5.L?t!�0ȁ�ӿ}�1C��B�V�J������7ӷ�-��q��c����wߎ;9���M��Y����į����;~_�9&-?\�~��k��,����ʸ����7��;�U_v~;��Uy�c����T��HY�R����%wLFƾ���M\լ �R���8�N����)+��W�&��=���܉i�Ϋ�˂�i't�i���sʝ��B3����w��8�����9��3h�&7(;W#N%n�S�Z!V�����[�&�V�ڣt���5^81��j��]��
����l-�K#�k6��L��I��>�����g�:_��(dNt�����X�չ�*P��4����vT�
�ߜ����rם˩:q�f_�
����c�7�B��@67B�6��f��=�C�&��b�9�3�Й�72󳻍���|�	��J���c+��b{�����q�8�Z-Γ�N)*�촔�n&#l�V���Gas� ��zM�׮���z�;9��hG�����p̰:MFf`��cl�`LPޘ��H'��P�]���v���Cu6��*-���� o�Q��f����QCzG ��iݕ/��U��0�Fu��<�i�@7"���9�������	,��?��1h�p/��7X��
�W�9�WG�>Ί�u:s��b-�Vw�5A�U���:��v����\[u[����o��Wߕ�w�g�{��g���w�;0�"�W�����trse�r�,I띾�+7��=
�%�������\=�>䩩����.�x𴬿����gl�z̯������	x���֖��~>.�����O����3駝6v%p�6i<۹k �V��Vz|v�֖j�k@#��\���2���I�ҳ�*!����jAWR=�˂������Y�@�fh�(�C�!c�u.�Ne�s�Q�!v:�Em�����f{S]�"��ꆈ���=��~D��M�H�#�b��n7;w�XP�k��X�\g���e�޳Ϛ�w<G����PBW�g8�\�V�_A�8�g2�$8�w{O�F�M^#�w^�J�y��,-���1u{��^z8��K:�`O�%�١}��ɬ�pZ���~���?�'��G����W��{ x�������F���ƮȌ�}��O>׳9��&�\��Z�aDዸPp�7�P�
;����q+t�"����mF�"졔��J�`q����wn�]�&S�F��M�D��G#�M��y0�<Ǔv#4+\Ipΰ��5�S�rhl'� d�j���F�9�3q�~G�K0�y�A�U��,������Lc��������J�[���4�AI%
��EO[����:��sǅ��I�2�+�˨�f M�ZDE
A஄_� ��)Z�l���ݻq>�������y=ױ����P+*֜]�p>|����['�-؏�)0�Y�~|�	5�����A�۴�[��)Ŋ�9�ߎ;�.y/�H��5��P����q��8,� �Q��Y�n�����?juR��Ӛ4<KtU3o	�u�/�d��8��bٸ�ʒ��βx�j�&|-a���$a.?k�Ų�ښm3T��C{!�o�<�"c����L$�h����K#�j�ٽ�1�Ee��>,�@y��ʆ/y�������+v��u��7�$��+vV��S�r�)xfof4<Qy�z�bFk�����r'B���֒eQ��[`�d��|��l_�1p#�h6t1��4�}���2�QUA��Y�/�i.Jk�2�x,#���>ڙl�x��<th�eI��8̠����(#�,�%�^�|�Ns&�,�q���x%���f�mK��9�'u���^�`.�e�w�Gv�(�>�fA89U_G�<o�F�����F#F��f6y+̞���m4�����q�`���u�탽Wkf^�Qa���kg�Ir���X���5�Y%5��` )h�0JA_jjĽc�b����16���l�x6ׄ���=�*������2�Zf����5��#v>@�>��;��E\"y�a[5(h��(�a��|ze6G=Н�<g�6{��<���ܗ�3O>$�ѫk��r
40�Ǻ��"Cw0�E|�U&�e����݆VEsl8��%�w���8�����sZ
���#���=p��.�i���^�}�+�����ǟ���1�z��<��O�����~�|��o���P?���VL�;���_��8�{*��ײͶj'��:ԙʊ!�3��W�{��ǸL�d5����ecv�_`5Һ7=d�<w�˔�pR��k�����RMg�B���"�W����h �`�eŃ����V��2wc�t�=�n���߿�5
|��t��<��έ��I��ױJ��w7��Ո�RVy�xl���{M�S\��g��wb���m`K��ZEB����v�����6"�C��5�a�Yk�KZ1nr~��:1�d�Bd��ҍ}��6O��:E-�1h`�Y����j!W�L؝.�m���S��7ײ��)FW AT���pR.��Գ��\V�˦�� ����j5��p���7�T�g{ӀO���b2��c���9���W�s�;�t
0�\���}��9��1�gU�V�y��Lb������A���.�?/a�I'� ���B���j�I3���|����J�즀�8{�7tV���ƚ9�A�e�BgimA�gaeFЪ��h��W�{��"(0>ҳ�o�Q�����p&V`���� ��F��J.����Y�ՋWa`�!���+�V}���9"�����?N:��V� �?lZ���N��ì�s�s�@��bx�4xd�������;�Nr��ӪL��݋�����X�j���S�<���<�~��[�+����o<u�<ʷ=��<�_`ɷ9ݏ����3>��sn���x�������(���Nó���Yo�|�ïK��ٮ&-Lެ��Y%��*�	���L�d?���2O����3�Lm[��ދ
�oTh-�R5^���k�x!��z.	�\ކCl�+�`��Y�N�ŘL���8O�Xj��l��代X�����xZO����#�u�Slg|�w��q�7�ta��2�fAS9@,�.\�e9^���|����f����o��US�9���\/�D�����������1�e���V?�Z[ֻ���Y��=q����z���G�O% `���v_�����,�ީW�Y7��fjh��A�`��ؓLX��<���IG�+;2dP`�G�,(���1t��L!$"Z=�? ��GN�y������K���>�`#�Q�9+"�u��̫4Ь���[�
\0*$@7�&ۢ�Ԋw19���z�&A����↴�5�31U�B�QEfA$r�:PtJ �"۱3���5�=]3�U����M�}�.,���R��b�}�/"�%�Z0�hхY�q1�7�,��i����K˺�X��u=�uY{Y����K'�'t�g�K���\�|�5>�-������a<yV�Ǻ��p(�uTL�W�h��zb*7����}���{D��{M��iW�/c]/e=W��7}iml�j�jUqV�(v�+���0i�j��"���هҌӌTÍY&p�a��J�"2���=@4K�撴��:���R����٥^~KLy�������%�?��9f[Ձ�� ������N��.Q�����5#)(T�h��>x�M��8��+��d{+�,q�V��f�Y9��O���T$�'�?&y�@i�%��c�!Y*2�����y �2]'�$D 
�{���G4<�:3��~2[�
o^J�<���+,u9�r��*# �Y���g�a*��+��ޮذ���[sA�qv 	�Yi�uN�N�ǭ)՟o%�{lUбW��LZ��� ;�*J���(OX��t���7-x���x˂0Q7d���j�=��"�n��������{�:7�T��,7h��Ts�XRq�"m��y�|b��\?˺�Ȯ2ҵ�R+��D�2���=�4�� ^��'�D��.����]-��ֈt\x�|���#��l���`�t�U8$��b�{f���g�+UEOۿ�P
�gj�>]���RS���s!{�k�I�X�)=�k�ub��l�p��l���ۘ5Z�t�s����	Q��լ���ց�k��rZe�'�s>��i8�O����V��k��S�y+|�/�7?��=���w���n����Ƿ!�/��X�U 7%��̖���uB�;3�Ze/V(2~M��&����мw�)�����^����5���>`k�Al�l���:���߫�M���!zݬ,����{�`�.z�Λx�����<��x"��{�1�x���WAw��w��Fg~^�>_��� dk��m�k�ǌ�l�0�l�aY���{aŚ���^��ղ�pD��y���sn6]:���
��
�@fO&�&��P��A	e�b���U�1\H��V�0mnU��5�6So���0nc,���#�h�
�^ĳ5.��|N��މ��ZN�R��l;`�|��gl��΃��0�X&�EE�-�5���L���;[��ZB�$b�0��n�
�(!��_�F�������ye���I���Y���ZOf/�&S/������h�������nbSz�ڡ}���j�M�:9�R�,����Y�������С�%ޱߌ���{d��}�V�m�/z-ke�kS�5��$t[��Мܙ���F����e�T�+�L�୬�@�HǾڞw̩⼳�3� �r_�[ȃ�����E��O�"�Rq���♭���}������ĹVK�BŞ��N�	$����~���sT;*^e�?p�]���<w�?{��4�G���/�x;x
}���pS���Bmo��ɷ��E�}
�e|��{���#>��f��)>�I�{��]3��<u���W����:�\���t9�O��������V�23�����RSe���e��ོ7�̀~c6�f�4a L�ƴq�5@g�����i�ֳ��PQ �j���ׂi3q����Zcm��&1� p�v�e�@ޚv1p�4�-�t@_m`~���!�N��t���A��?{�QF�����1�2���8�y���5���yϕ�~���Q0y$1u�S�[�L>x�f�պ\z�����3�޿��z�=_����|=q�D ������/�����Ͽ��~ᓻ�W.e���V����k4#�M�	��^D��trI���׾�n7`F�N���#�1�,�s�c�����	��)��st�0�!J��>v�4�zs���fPfo3UR�|iD`¹��h��zĮXo�Px��9]�5dV�*M��y|�B��c���JK]VȰ�Ge�Fo3(b? ����m 	���*���òBy`�6]�%43��зF�Ph�~Wv���a�sf��>E�F�rHsj���m���>�MN�_g���,�+G���&��w`'�e�ڐ� ���?��<������#+헼u��/����Ge/ P�}�ne3�� ����A@���<����<}��)��z4���4�'�=�i�z/�<�[��R�\F(e�[U9V� "��Z^����$Ƀ*��)6w䋽����1����"�	+�i��5CjШ]ܸ��"��tQ���a=�����5`D4�\�P��t�2Pj�lf�d�hr��_�����}��ɉ5����<ߗ�J��)��ʈ
��<��+���8#ۙu>3�z�fu��1'�*���"��{*lZ�w��d|��d���!�P�&��k4�T��H�(����:ge��[+﹭F�a����4��^dv�Pz3�Y�S�����bF|5�n�{��=�a��;KUf-p����~�i�Z�*G�x�\�y�uCAu ��%6ij,��I�j�7!�(Ot��Χ�9�!02�H����Ǆ3[�w���7��fIi���N̆uf@J��_:��#�Q��6C�h+K�ѰA:bk�i� O��M��Cx����D��l$IJ��\��c�@�^c/��P���V@]9�䱮���ؐ�/��y�d��x���o�����(O<��	f����������^�Zq���c�8c5U���[l^P)�6$p���s�Ab(��*�X�ʂ��{�Zu���g�q+�}��:� )���i-�H�8)h��� б�\qW]��	�P8�;K*%>yb�#Ey�*����4�Ֆ�\������4hg��?�c��#|����;<S����=y=e��q���������G+����b_8�/w��"���N3���]T��j=�u��c �\xOP��EP�\��iao_�b`S�]����2�
mt���^V�Z�y�C�S:�)7�93�h-��7�94Nƽ������??+�_T~�o���!��m�(����2��hY��"�mb�=N3�M�8�2ls] �ȗ�a���AH[�&�̀��p��>���C����V�O�d���zk	`2��������D噂��27_c��wǥ21K1�5qŔ]M�f����>l���#�r��N�h���!-�C�d����rn^��(	^l�t}�EXM���	[Xe�N�1�Zp�Cg2� Z/��sh�p�=U���ln��C�x� k��e��fpDc����9���
����d�%�д�O�c	q�KǾ܀��s��h����׉g���R�Z�a��F����Z��G��@�-��"(q�\x���:�`���<��&s`�)S� ���ƣEu.��^�p�)֚����[�gʰ $�=��é]�]�R�z���|Z�"	�n���3���k(^Ɛ �iA��]�괓a1l��������YŮ��#n�vmb�7��.�s������LVϧңW���~P!�U�!����_-����
�x��1�_���Rƪ����9�}�w��|��?��Ky�^�ܙ难~޳˗��m���׎�x�ݒ�
��~N;�~����/O3�
	L�2��(�6Zj��
t?�����8��p�����ٯ�������I��*_+��4 �����ߗǂ�VT���B~��z�j"2�����%��0�zZ��v��+h �H��Μa�/�!�@��%�-m�%����œ~�Ѩj���@b)�^J��܇bg��w��Xn'(nz��QB���GH��E'����=�{������=`l�0}Z	�H���w�q�]V��^��5�߂�0g�������������o���g^}��������ߟ�0�<_����|���iT (��x�W~����_^~�R߼�j�S���fF;�e��(��52P��ؿY��6��h��կ�o
(3���J=ntJ���Ɨ�����܂
��@���7��`~ ���X��g9���E�&��X�9��edZ�!,�*!������2��<6�?Z�GbA(MI�r��K���3�a0pa�|�,�f�jfkq�G�7��`�}DՀΎ������m�(��:��x����H�M�����@�����RԂGg��|gյٶ��&p�ە�e�%�r=�r�rڵ������bh�6�>@��J����VN�����5�/��)C�re'D������|v�O�B~�v���8����Z�yEIY�qi���\����}w�*'�Lw�N�a$��o�
�¨}68p%�9�y^�ǌ+]8gV��b��l�i:ix�F�"�;��	g̲�[���Q^���铱�����ƍ�SݟmF�1�����X�9�z�L�АeD	�{�0���蓩'/�;��&��)/�{/Ej[���P�W���/c����f����i�0�o#BO��ZY��"����K��+6gY��=�e6<�}�)���>65�M|f(R>�^���A����x(I�6�n���јf{tFtW~����'Ӈ����8E�_C}��d�]tBkY�>с�3'i5bPi��
��	C�����vô�?�zkЧgYs���3+Z�;PB2�D�Ø�48��g���\`�e�*����D��v�[6g�Q�ȹZ�C�$m�CPz�R|6<����;�0�g���\�ǃOJ2�;'z��`ЅD&JȲ�k����@%1�(�u��=c�>�,�u�5��C�'\�` m_3� =�?D8	�19���LŃI;�רt�u�s�_��;T��x�KG��fn?�C|=(t��[�Hs$]f���pv���#@O����1���i���F��h:Y���;o���p^fVaYwf;�p]��n1��+�4b-�n_��D3?q����}���~��|�����h\X�y�/�*םp��<L��Q8���Y��w�#�H�I%=��V��\8�J�>�X�1���t��Ą�uf�'�k��p>�Yȸ�EϢ�cQ3�QQ���V����}f�n��0���*K���^�0G�A뼳�R��<w���__��%}�Z�eae?��0�N�#��u%F3�(������:��w���Y�������cs�#��P��}�9's�Ol	z1Z��:V>>��:� c�x+*�@v�PѨ���y�;iq@�W�xU��,x̫	���	����\�g�J3��:�c����b/�<|ߌ�m͌N��%�����̌έ��ϩm�ga�x`_����(��W��Q�a]�*0��R������&���gt��sm2
�v�a����vM�=�s����Cm1�~=�L,���g�9�(;�ظ�����A=R�#���6�	,�g���,��N^��׵(����S�����jD���E�vg<�����P�c��ΙY&��ŏ�y�j��
�!�`�"�7�t�:��ҠjV��Y���d*���JX�>ӓ"��8���@ʵ3�,�Y|��(v�W��цV7`uTI�}��]B�"�!���#tҿ[�AH��5�]��xV˰@y&r��9�k��]�"�9g0v7z�*�v����%l�Խ9�ϻ��g}��e�͏q�/�nH��sW�A�B��򺝗LZ�-H&_�N��TAWm�U����E������z�ΪC<�t�c�9�O|���Όۍ\��qV 5*+��tT��yC�&܃6��9Y��?V{���OĖn3��F����h `a�S��������P�n)��:���'�/��٬�{�Tl+����a�3<�l6��7��/'�E�]�v�A����	�$�J�� �+�;(52x�W��ۤ� 봷�*[Sb�� ';/�k\e�|����o��_�O>�W��?�����y#�����|=_��[��F @������7���~m�.��fw����`XXL"��
��!aXA�?�a)G�EG�	~�ʐ�F���g�aw/M�ڦ�G3�}��`v{DHѹ� 	��ϩ�d���e�}+{U�^S���E�Qvks������5L�PK	g���
�+�M�FwI�F���͊s����
�T�v��%[ik�%@$#��w�Ip���ي��I<yˍk�z!���h�������и�],��N|�zډbQ�=�fTԓ*����F�}
�Y�l�5�f��ө%���}���[��e��[OK;mk�! ;BhKS�;Yel�H�d�@�t�a�Cr����(3,?�&U��e�!������n2���\OdQ'K�������Q���y5'&A�e�4h���m���?�֙2���?\ʵ��������?���9�Q��+K���EiL��-�oγ����T�y#iߕ�aܢ.̂*>V��F ��X2 s��F{�z���Y$r(��F��e�_�-r���.�9��6���pq3<��9Sf"#�m��eH��\XZ�d=!�g�:���/׾�@%:6ͦ�p�Z�z>S�i\[��݇g�c
ZVs~�zm0:R,II��k��tXV�Λ�#�[s>�b��<�M�Tl̐j�h�VWg�wxaȞ��|��lHK�K}�8�d�;�,@ѹ��ϲ���"g���E��_Q�nۮ�FT�2sf�G�ɟh0Kx��0>�>^�B8w`���yT�撟fv��8mo��9�ìvb-�� ��R��4+K�7+ 	΍�/0C�������C�tuç�Dfy;ʤ���a6����M��k��ō�Ӹخ��ڜX��2�����C�E��y�C7iUD�X�>�`%�����9���d�e\���
Z0B��?w�}[�0�pO晟Ys�'}fܦlF��`)��AÂ6s]ӒJ�g�nVu���{FGր���#J�Lg�Iu��D��>�a�c�k�sf�0�� ��/ƒiӅ#�l�E�p�y��ڎ�ժ+i9��$�Ttޤ�vF6���ث������� YuV=`�t��Z�Օ��dX�2��j����*KD�U�`v┶������foZُ�,��=H����KQ�/�	q��c�0;=q��'_K��	�����g���1���-d���t��_h}�ƭ�:�cǦ%��,�o��x�[>�||l��e&l�}\��q�L���o˵^�?u�K:���\��<�?�5s�TyZ����訆��[u7��m5s�\4J�c��I	�F=��/�.��<��ل��VTи�� �S�ڙ����8���>ʳa\��"���іٳ�A~3����,33sOP.3D�=6xV�������[.�q�����}^^�G�;\D��)�C����xJ�˵��^}���Uـ��S�Ӏ���>�k��u�k��͈�9�A�n�����w��0<>P��+�g��Ʋ5���͔��W4�r:�tLR���b}�MuF�j�����s�m�5T-\�=��BXX��"l�����z�V��Н�f1:o�]T3]��p���(�ؠ1K���L�.h��ub����7���*J�����1~a�d�宒6�!:T?�Qn��麱���03�t�
��5�R{cp��&?��W<�I�Z01+*��-��������d��zD��9?�7�&�{���6- �%�4�z��<0�2���bT�(���V﵂��HU0��6��<#\�5Pق)i�H	Z�DÆ�Q�	�3ԉ��S���c}ҁ:گt�f)xf@�V��͹zpq�jQ\;�ss_�mq۔W�]�*�6��\f�WzW��YpU�4�d	�k�Oax�0WT�S>�-'�]��354����u�2��>e-;�2^2��i�|�j�˛��Qm��ĚI~oo��c#�	���1w�ڇ��9@��a��8'�[������mcy�|��R_pe3�[m|7cx�oIc�:��bʾ6i�A^���w���]ǻZ{/�\�S�De�iM{b�������H���%��
�ND�X�p�ϖX����'�9CN5ZNZ�?� x�=0�h�SU�7�af�|�V-L.4��+�6�YT����XbY|�W�|��'^P,XZ����P�'e�H��	�:9���N�Qj�&�t�`IV���h�ܼ��-lZ��[4}b�zu`�����:�w9����Б�/�z��0���2�J
I���t�������Qm����Q}#���������o|�W~�W����d�w/����|=_o�~� ʞ������_�V߹�a��f�͕L�h�Ӓ���΁���:��L���3�R�,�w{�J���ja���uFE%@�޿���"�G�g����� �;Bё�$�.pl�
���j�[4�`yZ�(����0&E/n�H�2("�p��ǴV���Q���H<�0���ӹQll
�L{*�,[DA�.���VA`+ �X@����4�Ͽ�E�{���Ќ/0/ ��_�u�ψJ;ea�f�E����e�.���b0Hb�0ʷ�������m���W���z�/��~��\�U�^�����������i�8Y�J����O;�%��
3n�� ���@AI�����^� qq#Z�+�����p��p0T��U$o����ދÃUH�#�"M��ca���Sr��>���8�{kʁVc���8�O}��p�o�|R�����:N�%-�Jj�1���YS5�g�!J�br���y������6����js���* v-�K�7e�NU8�*oF�#�T`$p�o���7K�e��gYΒF��B�#��m󡬹���Y�hi�]����:�ѷW�ĵ}��}��~f`Oq��f4���Xc;T�SŸ�ܞ�5��W�Ԯ8�yndfkt�:�9�ք<�Os��)*9 �@I��u�lqR<f��*
w��yZhY�<���>�n�O�
��e���_:��B�3��H83e���#�`�ʱ�i���̧�o��[�
�=6��
�u��l��	�I�--���o�{�K;�t:X�9�=+�Ny�e��F����n�91�?-�ן�{�h�w�T�<���+p��+Z:�!�U9��?4�����c���D&�z���e�#e�$o"�T��_!~0��pm�.{�|�i?��x���H�hF0���0��/5P@[��l��C�5�x��ш���B�J�k���ER�G�f
zF�ł��0��^H��H��!���qj�G�jfŝ��O�L� �� �����Áϫ����3�_	�����Vi��Cf��C��Co�^�&/ѳ1q�>�s-���O���5i�$�2��I�^��q�-���{��@o����L�F�*N+�@�9��S�Fd!��x�4,j�8���BB/�.�\��^9#p��R��G	�lH���;9�l'Q�ob�|����{^�7��˧����J?]4Vm�c����V@AE�^�׍�%z��.$N��[YqV��F��m�ʟ����i���1",��2���
y�Ĺp�-��䙕���NEX+�<��0aE�u҇�&��PJU:l-ZdQ-�)�"�c�ˍ6��+Ώ�q��-�|�W��8mbK�b�ѠU;е;�O���w�QԱgA��G������X�ܝ���*�<<�,�ZF������o[V����M�߇e�j���nH-鬤}d���#�ς�:�70Oa�o�kq=���&f]@睜�欁!���}�w+R�뀁�l���ԅtkw5�(w!��ac�����<W1�s~s��x_��n*�'�j`0>b�m�{G�(d:V�
�1���b2�9���Q�Y��:�\�<��j�w/��=�|���J9U%��8�2i�� :ƺV�
v�����J��p%qO���t=u͊��w�Q�Ԋ���x��.��u�b|B���V=c]���ΰ���%y��{�׏�3`�6�� ���E�̵X+v*��ڏZ:t�����,З��k���
9gm��f+�P^��`K�).�Ń�y�+��\��Pٍ�펹ت!L�vT�M�W!o�Q�l�� �)Ar�W���ի�H��������^,�=ȃ��[��Yw���X�7,���x!����ʠ������I,V��*B���2�V��)�p	:���=B[O]�I���1��76㨽"Ǜ0&_/77�j��O���gȰ�%m5�m
� ^�
���������Ͼ+�ws�⛞k��Z�*ɼ�kz�����v^��1���n[ [z	��p�la���8؝U8���y���A@���_y!�WL! �e�'_օ��&Ͱ�ۅ�����@��~�v�A��'f߅����bt� Ἦz7���W��4g�6Z�L��݄�]6R-�N:!��q���7$ք�9�P�7 v���	�^H��DF����dU(�2
��9l8�W�������ɶ����坯��W��g ���qڢF�|=_�����t �r���s�o���?���>�a}3�Y��(4�yF��,P�Z�ޟ���ƍH#ʻV�0(P����@�l���ԣ�w���iȤAq�5V�:�x{�9$�N%Y�>�5��bα��˳z�n4U*�<���Kj5n*�`��3���;����R�
�0k�?�?�A�-�/n�� �d���tqE݂���3=��"�4�-�%03�MK��@'�\]{�D�,�j'�D#JU��@5yu�md�?*+�G��EX>.�!]u뽷PI[���f�?� <粂T��Z�wdՒۿu�������pǭ�V���4R��l�VN�fL��AT�9[�=*�ivVt�M%Nx޸^b]�w,;��I��b�@�)c		f?��إp^������&e�u�����lA����e�A��K9���qlt�j�2�kY�������E�W9�G�(�q<N��}+��v�w)cW�ݬj)�:�ų�UoʵDUҪ.�����z�{4�䜩�Y)�.R�3�`{��j��=�%��:�F?�������QvV�.�=qZϲ�C��<��Y8���x-��KK��k�gE�����M�	���`I�b�K�`����±\��C,+��J�0��p�Y'�{]S�1�V�gx�]��Z��@�j�\<+���L��q����8��2[�t�|�����#�8����-`�a�&���G%A9��h�wq`g������0鋽S㢣՜�3[����xc�bY�z���/[���m�r�j����M0�,G�_/��.��[�����AÑ�Cڰ��Rˋ�ƪ0f�'�:����4�툘OztT���������(�Q.e&2�}J#I�e�J�[ASA[U��6G�|�s	s8�h����lUaVA칶�γ��iA�Z��A^�����<��@�y,2v)׌�{�,^�U�!3d��z斠�!����M�Ö�}�Q~�`۰�<�A.�#�wƫ�`��Y��lY����s��Z�@2jf.z&N��s���4�j��l8:IRwdWˠu���N3�d��S�(�k�9��k�~�?�����򫿱�ݗ�]/��Ղ�
����6���;:�?$L.ąb�>���]�ub�8�A�A5��9��{�KP��g0;.̎J���`�A�WK=�q�h�r��uV�P�T�������P&�GS���&�WB��������J2U������ o�v�u����sjj��R޲>rA6��h�\1�H:S�0_�n��F�&7��܈5�-=L�즼���,�*���<�V*Y�;�b�pRK`�b�<��x�A��e�m�٭F�(/�,Ab�����{0�N�<���,5x.���|J��0�rd=Tmx��Q��E*�.+&U��-b���@)�V��U����y��Vp!���S��`ۙ�C����Η�{ �ғ���?�(p�
��Ra@��$�PyK1ќ�:"i��i0ڳ�<��i�6���*[��@��5Ͷ����g���?c���r����e�(�nggp8F��aъb������|ΆJVp˛=�E��ʪh)�`~��U���r6�Q%����֔E�t��3�n�Z�1��29�/���ƛl���U����2w�\��]OV=C+0B�)��1���3����;�3��`ǁ�=�����;�L�����@��VIa�jY����D��d��9���~���g�ťU�=D��h�_a����ۖ8��Ψeϋ�V������'h#]Q�����+SP��׭U���u�ӊ���ݘa�i�M\a��hA��熀��W�W~$���-'c�*�t�'n�"Ηۻ���I��b��=�R�	���q�;�lc���c�L����X�5�o�$�7��'#�,��V�$x?t/w����8�E��{�\�(��7�Ov(�,���������pܭ�4`�b=���m�ɦ�2.���\ΫVA��l��m�s#X���8;���ÄmkUg!,S��n�֯}�o]T�i|�3��01�{�:̋���,0�X`G���9S�Y�C�Wv��ql"uJ��h=��w��;mB���i��j����U�VbzQ�/<W��%�W�P,L=8U���ePF�8�5Έ�i��?_TO�B��H�+����D��Vg�_�@�`Arɰ��Ps��d��l��F���$����Jb	h<��$,�X��ފ����k��=8t~�*�Hj���W�����җ���W��|=_�����������}x���O|�����/�7���2�6fIkl�qe��ȃ ���i����#͠P�>U�l�@�]�h�X�2;���������O᪙Ţd��d��&���N��ŉ�О���t�%e�!"rF�O��n��������4;^�r)(?,�h�J]Y(�u�`	Pl��#@< [	�=��a�����a�0>���ee>�d�MO�~dPM�#��#`���J��Wd��^��B�XD�1�4�1.�GQ�.)ZSqEp�<�7��Mk��0�N YkS#ϼg_f��wY��#��Q2����Π��e���A	'�g4l5�N�d6'd�&��A���z��Q�@,+@jr(��2�V�f|�Y�4T����B7#�5�-�5Ww*j���ʺ/5���a��W��u50f����]L����S�'���+~��4i�O�X��qV�o'ip
���Z�=U�!��ގ'�鬺�� �cp�ޅ�T��Nc�~g眝�o��x��2�FM��ج�"��<H�T"���4z�Q����D&�h%�L�h��i� /v'�2�~`h��>���=r�#"$e���<;ÜT�t��U�ޠ��QѦ�bK(q4v9�K|g�M�����gjLPh���EC�j�,m���j$��5������e�W7\Р�>n�!�.�y�u�{ߝϺ�j�+���K�d�O6vؒ0cϜ�����9wH��̚Ϲ��f՞q8���9��dc�Cy��Iy��\��Wz��)=&����,���wt.��b��Y�/��F���q^�y�}l͇9,��*��XoF�mh��u^h��y:�+�&����Wރ'{6���:nF.1'����h��Qhhn�B�B�����>�3��=��cК�|�g!"@�q�1���$	��� ͒N��t�%��1Â��Ê�2���p=�Y���ğcr�@�K{�!�~b؆3a|����.�&��������E� ��:��ؤ���nNg<��rY +|]D��Nq�;��ε����傅k'�wf��� ����8)!�`D��ۅ%�Q�Xўk�Ϝ~���yM����2�Y󖩕iݎ��o�:럼@l���
5����X���4i�m�iXP�&V!B�-��2Љ�������L����E��IC�` Wa9z�Xj=�p�b)f�?� ������}B�jV��$s�wC7+��Q^dM@�:

]�i֪��(��>�X��ɜ���Ƞ��U�$e�V5G�V9:���V:�FOYZ��'u
؄������*��{E�%ʑ3s|�Q2�U{򕱛 ���H�
��_ˠ:Z�-��&a�Ϡ�%��W�6FȂ1$��/e:��/ 9b@&��^����k(��2��2A'����13�Bw�j���s\V̻T$b�D{�8�AT�́n"�Q��J�Q������j�O8G�܉��ΖL\H�P�5�f��
��RCV{Blu:�moQ`��}�ݡ�>�H�X����<���>-�$���M�"��?S����r���wp/���}���l�h|=��GXz@Aй��T������b�1�M4D�����L@)>�!���B�j�	�$�{�$�O�0ȳ�=�~��%�9%h'�Iⲇxp�gR!�Mg��5��	�NT3�ኌ�Ɏ>[/���R���Z�Q��m�v�<�!m:�-��c`�-�ٝN��q`&[_&}��0��`��Om>�!~� <(��v��ӆ���q����l���l[y�u!�`b��?�z����ew��zs�#��L��P[{�M���?3/m?��4;�x�D j��Ɂ��~ed�kN��.C�xZW?;h�-�����v���F���{\P��II�y
l�i\u�����Ž-.�
�]`�k��~�: ��=�5#�rs�%V5p�t)Nf"�Rݰ��R�:�8��Zz��Jy���p9����O,XKr`�[�`�E�r�lic]&�a�kԈ���]/\O���D�J�5)� #�� 0mD����}-��O�%󏣎C�4��[h��}�/�+��;`��?�^�y����u�야j�|=_����9�O# `����������o�������w�����K�K�m�S�P���#xq��L���Yi���°1�OL)�m�@�J¼�����|��T�Ͳ��i�rn���a������j3�ѱS,�mʁi3� *��c1!<�Y���# f&a(���jx�(���6��
K(�  �"����"�4��p�Jg#A���B���WU�  ͙�+;\� k��,�rg���5 ni����"�%Bv�g���:�3tʺb�{�6�I�1���=�_�h<۰�֬n�p� }�<��;���if��.�@��ݲl����e]�����~��������<��¬K3�d'%8F���O�Z�������Aw�`��t���y���)|3+t]N�xO:߶#��^_���t*�9T��\�E=�v��`0�>�]B���9�l�Aq����[=(Zs�tj���F�Q��N*H	`'e�AR�#rp��I�B׻�Q�=k],C��dY�*0,P�;20�J�6G;25���1,�B���+#��TF8�F�{W��g:Ϝ�L#4E-�Ose-d��ju%���+�͖�h �Hk���a.�%�x�%��-;�j �{�Z�l���-ַ�І��1hf��d�����4 Vq��a�]zmˮ�1������bU�H�Dɒ+v� �	� ��H�� I'�t�;���^��#0Y 8�)E�"�%>����{�^kf�1��c�[$�[g�s�^{��s�o�8l���D)#+zA*���f����ې��(^������1�Kd����W^�N�ޗ���q�c<�N�t�� �s�����T|<5r�����r<�;�:�h:��ɖD1~/�
w�Ym�2 d�X�"
Y�޳���h<��+�Yu��^s�ӈ��S|���G�%���0��?2�Z@���U�F��bVl��4$,VRu*^���ZU����S�=� ��W�������@/��q=�iy��#ʿ���1��bk匊��K���	iD�1c���\��t�Ǚ=�j!���(��K�(ه.�s���lb�EѺ��hl��M��y��ץfU��u;ZbB���|% �|�|�~����n�3ƌ��YmGq0s��
4�S���-yW�z�q�2�5i>�Mz����U�����#pm�@W���=YCƨ���ٛ$q	G�|�4�p|��}�����r3�]�}�̥yH�+�T���|U}0���>ij����Pm[�C7�I�aש�ј.2zJ��#'0���b�/:%����[����s��#�%�&o�}�̾Qa'�l���n�i�o�_��$�ADK#��Q�������z��<A���
�F8q�k�$�ҝ_����={��V���wS6w9P/lr����K���@%ʠZq�lL�W	�LP�LZK#�>�pO��N�"IZ�{S/N^M]���@"Co��Z-���ճo��f����r�����eU��7�/g���!��Wg����&��td�5��w����&�E����K΁}#$���by�N���ȹ�:E?	��C4���30da0a�9���k��d[	�I|^�
�8p�:���܏x�AA���0�ơ�����X;Ut���3(��$T��s��:�E ��a�E�]�q�w�Y�L��06׷N'�E�*N�=��Q��`(�c���������w,�X��BW;�����A=��2��7��v�;6d��C���Q�W�G�R��Hx�]e&�����������V�k�B@��9
����NX��z.�!��[1����� ������UG7�-��B�+�u�%c;C�0�"x�s7m�܆Ӳ]�&CV=ɖ��n��7؁�@+�"�;��5h�6yɥ�"����=�q��9-�˵�ز�ObG�k��0���Wr�gp�z����O�AN�UM���{ϵ��İ��k
*� 4PɈ��IW�y�`��Q ���
�F{�p�j�+k�C���ɧ���Ug�*��yC�v��$��4�rNq�g.�?e�{x�g�;?iz�5��V'�9�k� ��"�Z��6o����#�A�o��8��e7s�G�P�K�ٜ;�Ӭ+(�q�ȟ���fc�A[k&���{d�_�-	Y�:�r��s9gx�|�ԭ&� ��&��KnԀZC����$l���������^��'~2.��/^�����d���vZ��M3�}��������s^� �M&��ŋ�n��������������{ۇ��q&86*q j���p��+��@!,�9_���@dsR)A��@�1���Qy��3?W������}*��M{�c^FD�NA$�iH���G�G�5� ���~�[��� 0fu4��0`�ָA��������3k��^�G�]#���  ��$�L��aۖ�\5q���QN�	*.P�"���ڨLnҡH]���/���{K�����>eiYf�mڟ϶8�Y�nes�����2�0�ů����gw��?���&�>K�2�5����#�vG���7";w��-��F��Q�(j�Y��������ar{��S%MQ�Q�^̣�>ݍ�7�����b$U��<�#}���(Q��S:��i����'=M{���{������p�L��+�[Y���p1�Y2����u	���^��f��b�:fTLZu�YnMN���'MV�~�#4�^�������O�+�Q&���E�FϨ��UƖ�JG	�u�Nt�Zf��_-��Q�����%ej	��I�z�´,��"'|���:ҠgI6�/��Өq�|T�\f��P1�<��?}�0����_�L#֔�*<�^��rQ�h����.�]&KO��n�n(�p�/� ���-Y(v���yF�#>��F�gp[�efp^r�U�O~���Ȳn,=�h#c��������
��i��XrO2�J1ʸwS��.�?d�!��ѡ0������c�of��Xc���d%��o�$�jXK�{�K��˃ �d�m��97Zʸ��]X�����Xc���z�g˟5��ᬶQ��#��5tڦ�Uc�%�qֵ���>�UC�?{�Lq'M�1��%��Gie��q.1Oib�����������h�yӀ��4Ȁ�ZQ �2h��1X�����)+u)Ɩ��&�׌2����Ϡ!��Z�;�GTs�^.���S��9�����na<�`a��W�n��~�-���j�S1�\�@��c���*֕{��A�q�y�tLҨ؄�t�zȏ�_��ټ[�n�m>�)��n�����\a
^���h���G��p����F��az����dP&�6�Q߱W�S.�ï� �A'c�� .�R����2�`�����jE�����O�'�,�f��ゼ������*X�2P����*꽬����vS>�~Խj�?V�y୽�l�5�o���ك��z���!�f@����^:�¬Kg���Cy�<N�H5��F纟P���K�����`���l�E���6�"a°�V���~��\�j6s�������S�1�$�>�L~�D��í)s��>lE��k9��c�_R�`yV�Y��.�,?���&f�XS��J<\��l��p�я>-��FpI�g�i:�[KݓN�2����|Lc𻎰�,% cʍ��(c�y\���7�e��ŠV8TM2=���Lm�~����:�#o��-� [W5/9��֩?�Ɗ�F{�֬��lI�45��18_`��t�g��Y�i��N��Vv�4�jrq�Cw�6���Cm��YH�o�vV8���m�r��H
�lo��:ʉ���̳A� �޲"	�OۑW��q�0�A7��ZVe���ʺY�՜�jsaVi~�[��ʝ�Ck�!�b�ʳ@���^�.�ܭ�\���;`�� �B�x�\��jS:���C��X��-�8�3�	-�ϣcҝ��6$�J�\����F�ՋQ�m���n�Ck�]j�!��n�
�q<6<P,66>�]W���[1:� H�n�vr���?@�sGg����Au��h���J,�9�a����v2 �2 ��;���@�܌��q�7�#K�%���bŦs�����:�~ �}YI0��_x~�7oPY G�����q}ƶ9������ce�z�{�J�-�*ȑ�2`��'G�E%	*p#+��գ�΀R<d(��I� �,#BxO��l�����vA՚Y�s	;��Ul���Vl�T���-��g�uJq��u��,�UW%�M�6C�:�c�[������������O~r���>�  �ݿ�_�����ET ��w�Y�G�����G�Gw'�x�gW���PRl9�
 z'�Q�A=�hU0��^�&��:/;����v��.0��o����=9=���'y�����ַ��������K��������!ywځ��s�bM���G��m@�Ƭ��L�ٷ�$�����OY(� W��afz�c��z/�}����HK�6յ���|�B:2"W�3o�7);bL�`���kA��9$���A�798.��]Q(��w��co[^g*�ĵ#��k���ѥ셷� �'��,�J�3�f���+�=�>-X���DH�Ѹ ��N)~ �7) ���Q�aI��C ����`����t���3��m�tl׃��~�������M%�6*[8�iDu�D/e8���nnҡ'Z�s3�2���I׼�Gc�t�1�|��+B�����/��xl\�A��3�@Gc����L$Ew(���1�?�	~F�ݢ
��c�[Y��ʠc�����F&�⑑�2�����=���׈�a� oE�˲�Cs1(%^��)e$��H�*k<Ɓ��8�-�<f@��YR�!���������y��։紅B��5T�3~:Y@��eT�ZL�E�t�T�m�׮�̎ˠ<i�8���Rɧ��piaP�5c�t����7���}iR`#j��F���ܪ̉4���R>A!T�SG��B�dv�&�̔�ɘ�r�����C��y���m74�G��4tg��y�ne��&�f ��c�����%OΨ�cN��Vih,�Û��4�W�勏����y�o�ϘE�Qsb��Nޓ϶�p���W��\L�g�i+�z�������ڠ�u�j|��FZ7��;捬dU�䆡T1�O��|��oӳ��#���y-I8���[Y��2�]K{Wʐ\�U�T�p�}��<�����l'�A�0�z�z9�`�>�d:=�"�������q>=��+0�yoV����K?3x�K��{�픵���^�Jc3��	�!M'lo�����.�O`/�~�^�l~iX����{~p#㶯�)Z��^2�!����E��Egrf_CG��n�*W�'�'F-�V����!+���s@f$�C�5��)x{��] �|�;'�u�A-�,9��.'�U��r����sG(=��C c8��5U��t������Lg7*����<����h�52x�%�e�/�?��'��]��?�s�r��d�\���sf���ƀ0��%O��w�3�uL�����4^c��p�	���k>>+�,�k��+#{��-{+��Fĝ��;+|�<Nt�g&��Zb�.��q�w7���~F��{ pi�\��8�Qi���k�`X�r����.�F�J�·F�fڳj�`��zRK�)�� �L�㘲�@	:/r�SxV8/qoҴ����E&r���Jnj��U
�ά�o&7�@�:��
rZSP��(B��z�+$��k��0�U��	ԯ��-i��k ��3֘�;�K����Wd���гigʳU̖r��>>/��"/l-ʴYn�����JC��6�<%0��+��V�%�6���\}mH?�:�ǢR�8����yp�I
�$��)+�#Ω'_v������ �lݤש�B<)y��%��>F�8KŃ[)0�QkH\�Q&+E��h��Y��3�:�?Q���fx������y~��	��m_�9<pi#~ʀ�9ow��לnΒE���2[b��~QAj>˫��x��B����������'p��G�,�~@���r����^H��#&��`*p��뜳W{�6ۘ�,|^s����sz����,|�o%�O��1׎����v�Uop~�b��|ʹ�NRF��X�q�:�ցUn��������tm�#h_'v�LkqML!>�@��[02�a���8X�k�Λ�9׍�X �fVU*��_����(����<#�)i.3�s�S�j�<��gUm�[�fC,�i^�1�(F�����NC���_{���h�G��ƫ'>y���z���5�w띟�W�������}vwk����M_άH�?j\,x�xR�!?S��H���~[VIIC�_�KOX�A< �'��)�����7�~��?��²�����u�����/$ �+;3�����w�������?\׷�������f��|Y�k,�����pi��q)вL�|yY����t"�?ޚG}>܁�[����O�����{�Nw	 ��q����^g���ww��xi?������g��/�]�����)H,���d�FýZd��
���4 )�6��g��!��4ؾ.�-Aq\-` ���iyBK�n$���]|(Ik���,��ƍ�'\a��5F`ມ���89�k����_� �5m0$�ҷ4���x��0n���\�4�7��Z���+��e�4�Ō����p�q$�)KG�0�c���u�9�ˊ ��P:ܡiC�����qd�p2G��	�V z��d��F�״�h���㼣iX(�h�a�^�p��5"Zs��s^���gֵ��m��d44*"K6�W�}�����J�=�`��� d�!����T"8R����ն���kW���T~�إ�o���R���0��8ϴ���M>� �
���׋Gw�x��p�.��-����d�S<�JMJ��Ru���u�s�����@Y��(44�ٞ�u��>���Y�aY�.�lh~���`��c��8)���TJ�w�zB[�)��{��W�-KQ+2{irs����Y��=
�H�5#�a��\�>�l�s��֍�"۰V�=*[��C���~�Ш�ʴ�#���Ys��l�Α�e�<�Ρt2��@#Xf��[+�T��1h�r�UϾÑ��g��np:�x�3��8K݉=X-�(><�e���v��Z͌4b0C��\��\��n�~u��߹_� |��x4�:��C>G�9>/ 0����r�<�r?�q�x������{���
��׆��)����u��50��!:�l�<Dr����4��h$D�^��(���hn���i��ʵ�X����=T����P�B�H(]�C�F9�l�a-A��gsc&V&*����K9X�2��� ��� Ȃt^��
�m~�D�k̺!]gPH0E����`R������sulV�wy�QQ�?>�%#9�.2i�̔1�<x~� ���&֎us��쬒%��d�3��\9���UB�:�-Vr���N;�7F��x�6�I�ƚ0�8��i��;��-�Z�����ѱ+�&a���N��ϒI��!���wb��[�VqZ���t,���C;%:k�Z�Bgd`�Z�YW�꒹��X�-N�)�ay�6��ZQAy5ӝ�`F`R�si����z�P�f�g�P8wbS�~*Y���
*hMsάO�1A��F�x�8�m�
(=�|���_v�}�k�F��8�b/���{$Y@G��_Qn�e�-�tl���&�Mr��Y|*�f�s�{� 0O�Cr��!>ua`�f�N�x�q;����<C9q�7�3���KZ���O�� �M�����m�p�g��K��d�@��Z�i���u�1���~M:���7�>;��s?ೡ5&!�я3J�׉O�U�A#��>p}ʹ���V�<C����U�68��(�l��g	��@�yi�5�g0��:�9��y�|�q=�j�帉eӞ$,i���q�����ϣ--������ER ���-m�ނe���k�K1��i_�&h)��EF:O��?PG��A�2�e��5k�uʒ��t��6L��>u:�#��y���I�dP�9��!������E�Ȗ9�5���i#�L��+���Lճ����\[��o����S�*i�a�x�;�*nB} j����&��F��L��^&\luHV��n��I�n�j�̍��TZ�21��b̎ʹ
]`h<a�#�*�ϡ��q���mhmc<�p���s�k��#�Lʬ6�v��H�3,:y&1:y>�_%�H� �8���ռd25���Y���ɓ7��o�GO퍛G���p�s[B_AՏ�y��N����g�}r��>�}a?��G��.�^X�cN_��"(��^#1l��r�Zjq�	�'���ρsWm�\���/v�^ܽzp������x�g �Ŋ$�ݿ�_���{�B >��������/�����g�٧�m�x�"�Up����H(�lFSQ8��[S��`,�8eN�f�����=_���b_y�ľ�λ������n�]����^�h��}`8 /�<�% �.b�͇'���;�Y쥭��O?�?�����]��=Xl����y�rcDݼ�,)n�}gXr�J�_��ם6)>R���q�ٿ4�/F�u:�R8�Պx��G� !�T6�ܓ��?N��y@�d��7J��}����@p�j|V��u�L*u����
�QLcu]�(��S�+2�hh��7T�h4^Z��2�dń���*�֗ixK�ࠕʦk�Xb�3�@п��}f[AIfOo��eY'�;��P�i�0ϼW�#�a쁶�Q������ڐya-��,�v
��)��q3e(���|�呩�Dpo�W(,�����f��%�2�+ʪ�Qd ���D�TO����d��%��|SF���R�P����:�c��4A�A4Tf����8˗�gv���9�����`�A�/0�-i��*���^�O�;4/*��:*��d�X��TwR�!O��[zm�����dvSk
�Y:;��Yj�F$k�le��R���P�Yfw`��QƳx�b���W�����N��QeC	#_��4�p�6)���1Jxz�+�VT�����i��R{m)����m�4>X���ϗ��r�,�8¨]���]]�}���Ej�R�Ϗ��F�aI�4�ӨZ��f�¡�*�@�i�7:u�b�T��K�8g	H^7#w�U�|q�M� �8ߚ�mIG�t�,�+��a�x�sc��m�K�8�����!㖜sCHV�`�*��ܮ�bb�J��焸�Ch�ކ�(���w�w2)�|�V|���3�x(K�:��t�����I���E�*fkb�4T�X�f"KC��{6N󤞘S]�,�����a�� �z������i8V[�#̋�7~/�4��8�r�����~F[�t>/��^m�l4Zd�Y˾����6;r9~�c��~�s���^�L6D{0���20��O2^�����_�	<`�Å�|�t���6����4t�Q����<~/�[�cT��-��pց�um���׍��yT�lj_�؟4����� !�e��󜘞CL%:D��eDk�������g%����F"0��K>���4��u�Q��Fz%OVv78�|;���YZqOj9�{����0�o�~-����Cvל�#�/V��X��:�Q�hE� R�c���:�y�Q��m2H|��� M>��[ƪ��S͊������k�#����W���Z�,�B��䓁���ۑ�:�72����T�C���-����Nk�rf."�ГW����v�K��t^Iw�e�*#Z��[�%���idMt��f� ����G�sc<��dʆ�@:u��+\����m�U��������#�,��X?�N�B&��4�p��Ӧ���wљ�-��=JPk0�ɠ|�5r$mi�g��ִ�5=<��=�<7me~���T:#���@���Np�RI�q�~�ǜ�f���H:KPi�g��K�8y��uX���ր� �1HO���+�T�(2�%	K({6^�h��ӐϪ7��c�����=Z$�б�,������)طi���Û
�,��[���ASm�餉9&c���V>*|�gп�0K�z"��v��x��w��$�}@bĽ�f�uW�h����V6�P����!����0��k�H�vQ[���y6�T�Y��bB��f�)s:�̓_K�
��D�N�"��ԍz�<3�>d�`0���9����֌T:�[��Nj�?�6�RS���(����s��6��ZĽ�k��C��2��:�0��!fi�z���*��Bp'�\��^��G�c�sj2{�U�5p΋a2PN�e�-������ϣ���4�|����|��~�����v����-��8^m=K�{��P�k��=;���Ƕ>���U���K{�'��/?������~n_��'���U]~j��t�u+��4��%׭��[���v^�^�ݞ>z�ٓ7���rjnn�޷ �ݿ�_?���ip�{�O��������//߸�q�R�w
�V���E����~ŀ@g�P݌%�]�N�7��f�v�_����W��K��7��-�ګ������'e������B��s?F���Re�5O�O�K��5{y���~��ÿ�s�d�	ؿt����`�Qʳ��-_�㢔�`���&����}����� m0� mT>���䌉gB����d�53�i<�r�H˖����E%����uM�٠�4+cq��5K>C*�w����1Ͷչ��X8�+:��*��&cm��	B�ю
z����;MG�`�\��v����f�Ө��_�%FC_.Z��ve��m<�0��A��n~��з�����Q	%Ĵǘ�gs�,�xi�AgQ�����C40d��h9�,d�� �u��ǆ�Xe��g�z�wY�\A�z���p����nN')�/�x[��&�9�:�t�R�TJ�9-v5xgA����QI������t� ��*��h��Ȑ�{&��2�i $�c�-x�6T���9c��T�Xc�W���U��y���%^k1b99�(�I^ǹ��/�?阤�"o��A�P�b��f���S�4jg�w��6?5xH
��1��KGtc8�7U#�^9{���8��<�:��5��춑�[��9,=#�������&�L�|s�0�����,��n��y/�_��״1F:8~w0�.��Ʊ�5K �W�4eĈ��:-���0Q�z�D�g՗zy�t���3	#��F#*2w�\��n���$3��@̕�a�,�tN���4�F���~��x\��p�{���cO�9�Ϙ;�J��!��\N\�)`��R�Otݧn���qܺ�3|�|�+�:1xml���v�<΋y+��g,�Ώ�1�<���x�8L ��q�T���F���UYl���G�M0n����iG�\4�i��?�'�.d�r�(̖U�c���4M	̽��eI#� ��������=	��o�0u�y:�,x��J4�}�!�ߜ_�[�s�'��i��Y1�A{���O��k[(��k���K���ec(Hm�͞�"�1rK��CVwZQ톥[C�C��2{.�Wk���P���/{��ZdPG����)���k�}.�1�$�.n�a���H3��ᡣ4���NWy~����dq�ج�E�o������al�s�4K�*@��[�ߌUl�����O�xY/n��a�aɏF:cOخU�zf��Ic CV�Y���7Б�@�C'�.���=�=����0��p����˲
A�2�N�ZA'�@~ִeM�j@!׭pe0�ċJr����ΆV��VE�o�ˡܐa:vg;K�Cfʸr$7�G�]�����d��Ĕ\S:{����[���� ⋁L`�3�q�N�_+���G�,��}#�����Np~#���O{��夶�*�\1\9���.��lh�`<]��B��xNc<o�c%��3>A��HC$���V![L�sl1?��L4����r�#������|�Y� V�C��ָO*�o��D�[2Y)Ġ�֠����3�k�y�¦P���{�������k�	�(�+��t~s?�\Tl���������e���,:tɗ�<ʻ�3cu��K++�-eߚ�FA��ߔ{ɛu>�$eY�n��16ǲ,�T��l�|Ѥ�Ă��aV�;֎�v=;��l��{���K\�!hqAP��Ԣ���]�s���r~���*��.:m?���~�3�8Ȣ]�l�@!��%�I�/�*x�܏���Ǉ�f�jnv>߀΀�fP�ĜK�]ܱ�r��$:��{6�"!�7?KXݤ���[+5ļU�S�:���>�y_�m�����5T��1N���^���<1��c�J頃����Ö
Ǒ�S���ɾ��̯2^z��>���3��^�������E������M�<$�ŀ�A6'�'2�S(��*؇��s�W��͂�b���}�{&���������B��Fsf�/��x�?�����j�=n���W�;٣�<o�N��WoVE��-X8��v,"	�uw�����{�_�������3���o��͵��&���[;pi#�o�U�0(w[�O���i�`gMt5�N:�m���?������~�dïwk��������s^� #��2.��?�����>zt��g����.mmQ&���=������H�M�J�c�o+e��<�v2�s�H�������l���ۻ�����j�:{4=���S�@Z-0X��h\��|:��v8�X��]@=�qȳgoٯ��E�ާ�ؿ���>~����.}�Q/��b�,��m�/;�v��K� �Q Ei
�ZU&���r�}��%�
�W���މ>��1�/��[��/F�u��cI���%hK0F�����2#�A��	��l=�1Q�� ����oN�	���|�@������� �DÙ�Yr�� 3A��GPpwzځ�&���cf��K#z�0���Y��ޤ|��逹����{����F�����(��s�ޅ� �KC�]Eҿ���'���,�+F��]�06�18�1�W����K8Ϸ;S79C�����͌�md���8S���+ؤ�9,�ψ�t�F9wF��� �X��wd��A�0��A��|�R��)��t<3����Wd͌I�7�vKǽ�Ö����ǂ�42�s�Խ�h�Y�4F�96cE�1��� ��&���De	p�:G��g�D�����>����9��-�a[1��d�ѧ�#�tڒ�;2����� �W��a
ZYt�P���Q|���*��,�=ۂ�9�N�4�p���6��/���!�Yr ���M�@��W��B�̬8���N�y�z���{��J�<�/$�,�>tNh��`|��"F�	����׃�x�:>h\RUK���l�/�,s�P�&F������8V�gâl⺦A�#��)�*�Դ�Z���|�� �&�:���1ƚ���`Ah�/;>O��̢��/�q1���!�h�.�<��2�kˊB�e�#���)��@�/�r-��k+�%����X�j=�.�������RLB	��秲��z%���fֳz	S�� h�����I�s2N3�P	�a��%m�9�G(��jIО��x&�Hڅ�s���Ҹ�:��ғ��[��8WC�	\�;~gWCPh��@�Ί�4������x{h���J�rJ�BA�}1Uk���gt9��t����ޗt���4�A���`f,`�51��b����-�\ւn��T��U�Y8J�sg�2$��C�ok�����`�}Mߗ�q ��kE�jt��� ߸�鴈�>Y����[�m|o�����XG���/I�0=�a�,�r6�q](��iY�}_����K�O�,�V���V�[����|)�dsN���ypx�0u���M�f���t��ß>>1��Fe�&�/���~�ko�������V�cY�X�\3�� ֽ���J���z��},�~-2���J_�5�@v��s��T̲� V�ʌ٠���꺐��j�H��`s���1���uefyN���gky�4����b��h���8�"�X�
1��ц���j�I�{Ӓ
pa����?��
 19ΧÞ�wg�J,�9����-���Bڬp��(����P�5���Ў�x�=��HO�E>��n���:�1@E��蜪Y�C��-3�yU.;NN�Ȓ�H�H�!=(��Lf[�nTZ����ObXE��3���͝�c��̯tM�h��m�h�C��� H�)�Uޱ!LQ����JZ�l{�N�<3�����b���e�6[$�C
��EL1ҹ6��I�{���$t�1��g�;�r�͘������fe�hW��g�}CC]v+:O�à^��� R
����#2����N=Ы@� P�D}��g��u$�4���`�-m|�qo�2���?���&�{D�䤍v:���Ϙ�Ӫ��N>v��zp�v��O�c����������C{��Z��d%m����5&:��p¹�9Nf��i������y@���	b-q���?Ͻ��vJ�,�������R�]�]��a�e��ӟ4Z�zU���V��B)�Q�j��Ɓ��,�ƕXd�3)�9�Щ�e睸'�s�.\K\�gŵ��Ū%\3�db�K�G34=�JU�:*ª��(�1�������=��gH��~6�t��7�`�����x?��;��=Z({���D �!����T]bD�y�C�������p0/]/����㡽��7�7�����i�������^�#��4�*�y8��iC�4�չ,4�Q$�UL[[S�%�D��w�On?x�?�/�����_~a?�O?~< � ܿ�_������� 09��g���ɏ_}���s������63e����5��h�da8C�+d�+�}�<]ܐz�u{�B��ߟ��������Η�oD��;����h�f�^K������:�����,��0BIE��]X��<�D��]0?}��~�7~����'��?����.v{s��m {�ؘ&�ߙ�H�ി_N=�M�:R᪎��H!_��P��$����-�sc�!�hT���A��7Z1�"����
<�	6h�`�hXą��u��T�٢�UII��B����;,�:�Z2?jvI`�Pc��1���@k�@�Pb��(ѦF�,���s
z*�e�,�U,=a��3�0h����g!8 ���1���
����I	�H��
q�-�ɱ �l \n�@�L��	�$�y!CC1�+���"�4�i(f#"�[T"�7���gv�EC�!Pa�o_�N�9�k�؛<��\��°�`6Yxx�gI�BMc�A%J^��z�sڕT�go���a��QX�7���4���|�����
x4~:@h���b��H7Ь�u/��k��ޮ����dS�X�7Ayg�2<��P��A�vk*4<%�Y_Y��"3�ߧqmdFt�I(�s�M띆���
�����N�jx�=oԁ��/�`����y���J�g�A\G��VRLӀ��Yr����Ƃz��Ǳ0(ŝ�<��nd����{���r���EEV �,ű���Q��wN�<��p���Ȋ4�U'��?�g�CPR���0W�g���{��qMO�k�glsm��80`��ś����GZ�LBc���s�!HFV�F��Q
#Ca:��|�����w�x�0�����D9��S>s�eXcL�(i)3)X�fD	�ro������N>2?�� ����%��wZ�3Y6z��A�|�J��Lk�E%��<�%ƨr)��=6�
�8��Ӊ9������>@����Zn}�3[�u0���]d����
6*-\!Q�V�$ic��Ǚ���8jo�'���;8��J�d��4�N�qZ�Z��F�a�%_�G`���Gf�͐��o�]�a�FΛr4pM<ۋ�n� '>u=��0V�ie�hw8�Ȏ_Yx��lђO��>�-����7�-�Z�����Ľ$ֺ�fL�aU�c�~	x	�4p���E�9��#�B"��Wus�)��N�j���5c0��"r��1�8{�wr�qG�4�K8�;q�XMc���d��oɳ8�!Q�"�degՍ�_�J#3�&�R��/)��$��C��k)S����'T����c̝�Ť�����(�����X�lgu#�=__t��6x>3�[��f��3e�0�����@X*����R����a���h �\��>��ȅ�ޡ��;��^N�=<��0焊QS������,m�L���sB�pV}n�|��S:f�غw#����fVfظw��(�b_��y��\cm�A�74�#eU��t42����Op�	k��d����v�
�>2\)��ǀǈ+:�	`�:�7�h�tV2?�b	��Uܻ���T�w`��v9�eˠ� ���-�m���h���y�mf��B{�{���(X,��(�c~ƯS�d�	�BY�&�@_iN|�i��5�2cq�Q&Z&^����1:�x"�
h!��X����VB�ĺXˊ�C��ҹG�x������Y]R�T����~֕X!hy��~����U5(��CaP_���3�|����L^6�8۳����-�U =���ɨo*� &�������>p+�Og%���z^;��-Z�0��I���ˡ*�x�����jɋ|�Y���Gu�v�2��1J�����3��!uۤ/'*�bϷ��ܛ�-J�,'��?��T<��5��ß3j[y�h�:�u}�))�\�m��2?�F�C��_`m�M\k���
)8��Á�#�0mg8�=�o�l�gИ�t�y�񕸋�2�}e�&n��f�����J�Vp�_�ދ�[�J��<����22�fW{����ҙ��]Z)�_��W�5*�n�lMgc&o��f7���o/����7�ן�m_8��i�	�g7Um#0��j��Re6�%�A�@�j�c��X���}��g{�ͯ����W���?���a�ά����:mf����<�:|E��S�3�pkx%�H�+Is.�z�������٫~{�xy���wO�����ݷ��������?���U���u��ݿ��������P<mw�2���O�a��A��ed(
(Y��ef07��eoW�'� ֝w?�{4{�v�W�|۾��/ۓ��k����9��n��'u�`N��/i��\����j�`�o�(���i��������G?z�~����G76ә��{#�r�@��'�繕��j����Bi4�2�1�W��+�,1�z �= ev |E��w���>�O��(��`�r-�2�qC���*��%2�XF�Gdif��� *G�5�Y���������)�,�kX����(����RA ����ߩ�1C�X_��e>�0�T�.Jng٬y��ё
cD�f�+�T�0ǖѣ
 !�����_8l�o�w�ˏ�<W��{������I�m��WZ�0sǨɚ���vT��_�	���A�Ȓ����%�y J��tp-� qd�e�9\��i�@/B�.�1f���2��e�e4� �Eo-�c|m="���yBI먮g)���y�C�
\��[�ȝ���S�tpf3�U�W�> 8H[���J�I(=��h̩k"c��!�kFQ�&3�����`���!*MY����^�]�4o)�647�	���Q��ݠ��u����#�Po��%T�Cd>~ֲv�E��,d�6W����D�Ҳ�����g�B^V��d�T��)�h�"	�NbYb��8&��+�X����5?�������P���rnc5��߫2`�L��fVޔ3��^1�w<�,L:6�L����t�L�܏R�4���@G�V��U��A�5i`;|~hKa�'�f�*�\�x��x���p����)�3��"�'�9t��3�rλ���=�Wh�"bSPK"���6qH���!��X@|J$�U���e	n��|y���|����̬F;��K�p�����s��_���)��,��������N���bZaP5*�]�D���>�(H�ǀf>�fl����֤i�5�7T��A]|����p�!����xʼ�lS��g���q��NI;��ۅ6�mE���g��)�I�p=��=�,�M���܈5޴^u��oP�h7e�T���$���,3c9��.��5���Q�N�y�ӱ�G�\.�{^2�\�Oz	�+�=���on��Y9d����t؆J!�U�V�.�0bV�`���	�|EGX����C�rю���,������YXM-^�r��m���f��!�9���v���>
ݔu'=e f�%��������q�M�$�}�D��c58:���"�D�E����4˵�t�zd�x��#/g@�>�� 8bP7���"�AL�c�:�SR��y}�D��Š ���3-��<�� ���{UG[Du=.���UF�+rЪ����wfFl8����1$P2J[��p���S%��'[��-⎼bN'�1��ԭ ��j��b�#�pUb���GtT�L��65�~e]�+Vf�k5�R 6�hv|ׅ6ɔ��"�������2����@�غ���\�f:��r��;��TYI�Y�e5��Rg'�%�Fb �A]n�1�����8tӸ�X:�y�H���"�%q`�eP��*��	F�V�2��R���@'�1�k�[��HS�	=����k��q�����E�����W�.�6d<��\�K�D�%�S1��_���1~�M����9�^��u;b��zШWbr�I�\ð�iG�Z�b�����Q0����Ld�>w�U[Mڙ�p���s)��4$m����kƵ�z�~O%D�H:NB��<�v�,�\Vwi-��@o�yZ�.�8�Ȁ��~&��9��ۄQ��S��bg��w.�7�߳�]��������w�����_�/?}�}"�^٬��Ե�0�i��|H��x�إ�;�mH��uқY���F_�e��|�����_�?��_�_~��}x���h��&���'���
[<���k6�c�Nk$��״�ڗ���ˣ�G��������u�*�_D @{�s�/>x�~����v�:�dل�	h��k�.gb���FH#B�� �����~i�n{d������w�Ox[��Ol�k  ��IDAT���hM�� ��M�˪��2K��0h�Y����#�Q��>�`�w���}��[���'�����晙sq0��fߨsdv
�Z54'�pC���Gg�=� T��:+F�
��x����b���)j�X��8)����B)�@��u0���a㕒ޚ�C��9�� �9�z�(5��xD)g�����Sk��Zʛ@��sm�9�[��R���� c��yݺ<����1� ���%xNe�����Z&I��y-��/�[T|_Ϟ;�؀էe�EH�Ð����Ǣ�p���籽Fm��W��%���T��0��������8��������q,}�Ry�&�`W�����~P
m
�9*3������̃��94��&t@uM.�n����V���k]�Ye�E9���g��O�q.��8ב��{Uc�q/�z*4�����֬:Nj�r~^��c��8�G�㎌}O��5a$y=p����,��b �X@�U�<Ş����a�S;� ��@V3x�f�ܖ�#]���+3%FX����6���sA9W��(7Qޚ3�O�@����<ĳC� x����P�V0�ߜgt��a�|��䩵����b��t�q[2��"�}E�)� U6J�#3Mt#�C�R�Ʋ��YY��(F���s�%Z�J��mE�\Բ�3�w+j3׮�y屜����ƖUʧ�5o2<T-��f{�}���p�����7�s�y���!.L�WKf5`�t"k��sI^�w��i��m�<O4�F�]1ph�{4����8�bOY߃�4 :���Z:����^s���r�[�
R� ������.o�0Rz��$�Ij[�/{��A­�7�C�:� �S}��O�}����ͫ����Y��B�X9r����疆j��O�sURB&y�h�Ǳ]�=���]�(UƐ7Oѻ�Gs��+�H���]x��Nt�J�����Q"o��n���%��
�!]�-9��r3�l�������4u�2��扌p��s�|*�"vZ�A��H>��1ZV�к����,P7�r��*�`���-��0�B3O�|�X��9�n��?�Ƕ�~��s@��-h��2�T+�^K�\�◔M�k�g��E�=�#�}-X�s��:y,[�tc�R�	���72�g�~�{�i3�&uy�V�>6b�E�0��e�|�NQQ,�&o�>䬞�^֒D��͒�P��Ӣ���Qe�ֳ��ϗ���Vd���\�Qx�Z��I2�|3щ!k��|G�Б�b~�`����课ڃd�&z��2��^��4���8�Vn���ţ�k���U:��P��gȱ�˒*k0���hJk�"�aC:I��\+���^Q�n�� e�N~��wYe%ֆw�d�rpa��-�^�|G ߑ^e��W���d� �q�G�m�������C�_9okL��)��ݔ)�ۺ��~E�
>��y�X,bU����!Y%rKX��:c��<Dj�G|�jo\7�_��;O��ِ����[�1y%��J�A&����g��޽e�9�_+�1�}P�A��붖*oٽJN3���p�>�y���dVH�^�:,I+:3L�@ ���k}��xƎ�'x��Eq�y�+���O^�x����h�IL�%�@��v���8���{p�MtOY��l��+>�q�wb_��l�S�K��c��G��f>�/�q�lp<��^��2�E���&�M
1h��6��\�n
��<O�<��ғ�|��3�o}���7n?��<���;�N�Ѧh�U'oj���'ρ�w�+�B�M��6�^�j �����������oٟ~�C��߷��>&NY7�2���J%��n/��ǙZ/��X�h����5�f�ϸ{Жq�|�W����j��x��ݿ�_��E ��7�����?��'����_~���ۣ�󻭅�Y��ϗ�� ���փQ7'(ⳟ�,����#��3�����w;mq] !c�ކ"�%��f|ެb�p췄젢gf�5^��-Ɍ�=��T�a������oٿ�������Ӱ���.h3���4X2A��y��tH���i��T� ��0��d6?�n���X
�jDj0<+*��E,��v��@@f�%Ȩ
u�g��fI�V�{�S��T{D+3Õ�x��˝N�@���c�R�
k����72Z6�����k�^l�L.���@�p6���J���tp�RЩ�l��Bŧ���(�x:=�<��f����#�� �1SzjSoJ���	���J�Nc��P1
�5d��
d��XΛWW�s1�|*e�Op�����KK��+BZ�']��Ӱ�#SP�ݹ�P���L��|�F9�R�h�X��^�`T�!v?"ˡ��eU����j�R(q�[�gC���wEi��y?�ņ}���3A�m�#�>{�C�<�<a��=؎����{5C��=?(�vU����>���j���E�G��tx�c����jF`��,d�P�K�G�9w0����Jq{M9	ř������̓�b�ss���?-KL��Jt�)��n��4��y
P&��?�t����x���tv=�����-�[��7(���,�G�����c�����2Q��j2�ӠD#p��EK]r����	f�f+��)�dfջր
{V�(r�L�A�D�kuzTyxܣ��|Ub��(����?)CS�f]��Lr�bh��G��s4д�>i��I��5����^���c�llM`pƀt�A��1J?E���i���W��&��kX��Lb;*��!��Hfף���_Ϋa�t�(M���9
+��@*x�`؟9��+p]�S��Gp�M5UK �ԾeDV��鼢H�^��t�r�ͫ�\��,'���1/+}'�[K|&�퇘G��ٸ���:1A�dЊ�;�1�}��Io�c+퀻��֤+_E{V��3����-i2����j��5��� i��!z=`�EXI�V�;��BNt�C~]U��Zp?�H�V�{Si)�#ɳn�z�{*ϡ�m��������_�+��m;=T�H�Ƴ�D���[?��T$H^x����g�I�H�p:��Lc�t�6On�=!�s�Y����˱�08�3݀���'6�m��ԏ�$�k��Y�ν���t8-N���:��Zp�s���
��F�(#tG߯��\&�d2K��B�)����Y�w��l\���y���ƽ빝���8�ǰ� l���)^ò�M��W8��tu�rB�&�g�ǘ�#&FJ�6�S���(����G ���M��A��2n�����Gz�������m��G�b^_2@�S���=�sc|L�"�j����
(�6�\��+����)+:%��-��~���}�4y,{�A7���v	�ڑg�c��_8qc�%��
�z�`�l� ����yT��N�#�@$U3�C宸�:�E>e>zO0'��"��R�1�^%�qϪ��Qh&��1����*b��?ku��+Z����9>C`efS�,d��@U�T�d�{B ���;o�����gK��@L�*�m�97�l���9I+�Ԓ:����K�ʞXq�H\p��J���ak���@���ڻ�ɹ��9��;YY��ѰW����`�+�,�ը�Y��S�dp��}�gͲ�fT^�EPʧ�!��x�Ea&^_��_�QM +�[>�M�m���I�Jڳ�����EI�i����\��s$�/�I��e=[>��1bRZ&�a���Z>��~�ď~ny�<����nOv��-������޵v{F���nW�C_���\�`��WRk�k�tM4OLuX �6���{J�~��}~�z�K���o��~�;���}�c�;}��,,�8$�+ct�[�e0ޜ׬��=^��o�����?��Ko�Ý�|�z����߿�_������ �h���g����������?��������l�0�G��E�=;"6���c�pd�>�o���o<���W~ɖ��.(��H����憟�S0"��u��+*�~��1ft����/��L����t��n_��G�/�⏬=�^F&�]A]Zt���wid��,�Ī��@�/�ϒ��B?�͍�P+@�qta�kBC�#�PS	R�,�7� �r/%�4�!e)Q� Q	c*2q9K�2S>͂n}١��+�\v�n���2#1��Hg���6|��8Y���@�5T�y�� �,U���oRF���[:أl��/0�o0���y6�t��\VdEi�A�{0`�5��J�58Й1��(tF������S)��@3+kA��,�ϩ���,1��lÍU9��O����A�fi�B��/���z*U��X|@:�����̈́�A?�K>�kF������4dp��̜������ �mV��pB�Q��A�0��Ke�`���P�ι*K���� >Rj�w�M1��k'~1��i���H^�����p"e)�T�R鏳5�z�ĞyFR���|��;���xOY��[��L�q5��#9�y�Შ"ɼ��)xYk��Y�Z	�>=C�<�5�_.����ٯ��V6A���Z�]f֌�L2���HQõbz��{�e޹4�g�x���2����:r`?�{8��F��Y���[Z��ȵ��6~/�h�̳���\j���z�C�d�F�tj�\���6�yVƱ0Py�����J���:j�z���)3�ZN��i��S� ����?��2��~�To�J�dytJsm�mc����s�
)ֈ��S��&F�����~���v]�[��0Ȕ@N)��C6
N/2�W���-�6��ѯ���ȉ�^ì�{c�,��+e� �L>!:.�^�Ѣ�t��8�lk�X�,���k4�"�#���z�b�4���0m�09��	�qlU���R:��r�/�o�;��q-��o?��_���<��Z�&������^2���+N�Rm
����#�֙x��Q55�a�_]K�%�����o�唡'v��1�5�Rه�:��G��\����o�Ҝ;��ck�TN�9�2s�^"(6�rc5>�Y�rhA�\������^�or%m��<�G�M��ڤ�3��A]�xv'<'#/�i�7�I�*4i��,� ��N�%��q�M�}&�j�*����؀=wf��	-+�KHX�vRU�H�V�y�
��0�6��<�X�ca�P%CS~^�F=��5&6�U�|n]��ǀ)zуҹ�� 3��+��k�����gu�i�X�,5~\sV��-�:�k\cUl�a�'*���9�8�V���g���7V�3�Φ����̉�R�hP���R�R�6���8g�M��d ��6.��K-(�:1Xo���t]Q�������AM[��9�u�U��F��<��!�:1e�*Mf���hD�i��&��{֦sg6+�GT�گmY�hp�@�݋%�x��X�P�a.f ����>�.��7|h{c����<�f\c\B���fýd��b�~��#�jX��8��}��bd�<�'�
���r޻��{�,1Ej���4�*:I��6��-'+�T;��,��^�oԩ�#C@\q��KH�1}�ݯ�h</������jϽГ���4\�v�u����r�I�̌~�s*��\� }j��v�G}�UZ-<��?[X�<��Z��:���V���R���ɓ˹&Mf@V�Mح�/�=�]��#��`�ey>�ƞ�l��i˜I�o����6���};��[��`�~~D7z��/Q�t$�*c� -�8T������m9�YJ	�'��/��ιc���b盿nO����/~l������^&?�U �w�\#��b�/�\��}������s{|�������[O��x�O>|8 .v��ݿ�_?��W 0#�&s;��/n.������������z�l]ۺ�3��H��� �Gw���-��Q�S�H�ǣ��;W����e�x��-�9�3�e�!~E+��[k	���H0��J�G����V�I��J1VFIB�EI�),�g$ق,���/?ۍM���w���^���8�E������\�$Rɢ��8�3�B;c*T�m��̒��(�s6(�\��+',�W���E����O�42
}��n������U�6Y*0n*-�qi�jOF�R�WP Ɓ ?���i��e�=�5�WTH���#�! ~H�R�K���Ԗ�z!���p����e*��%U�,}V�?���	�q)�����d�ѹ��� �N^�oÜUb�b���̪�˞m�E���:��C�A��Kxf��6� ��4&p-�Tn͌��[)ϕ�vt�q=�J@�|i�Z�m@��Z3����,�af���HP��ݱ^� �ᢟrx� 0������z�#�$��0���\+��s�R��Ӡ!����	�u���X̙����h�3������'�kј+-����wpr��F�E���/'K#${$��!�za,Yt�X��,[����R��F��>N�-�ȍ�k�Y�2�v4�)��[S����[*X��\o9�e� �z:H�gekT��uy��y$� ��b�t��0y91K�l�#�q�����$֡�;�����{%���(�aĂ�j$�JFHLN%��:���
�R_�c�$v˳O�5�=���I5��׏�Z���hQ��$_�(�x��R�4*Ҡ��l9��:i)�� ���"���-a��㌳:?����-���1`#��Gx�Ӝx��uq��e��c���K&8�V�2��4�½���\�{ETW�S�f��1���%d)/�EU��L��.����b�\7fm����[���C{��\�4�r�\I���a�8���-[��T��O~iĹ<?��q~��AFu��	T
g}~�x��2��٢�� �����k�o�z�� ���aCi�Ut��\-�C.�"�z�_��q��W)|m�g�n�ŶZB�xZ�g�hִwy�%�1�:�!�+�D���v�yz��`�V��wD����,ĸ�*�k��k��>��V[�s��F��N���yɻ�����;�5�L�&�}�Xs+�-r�Q����\��I�m��6�n�*@����f��-��tljk�#�/Ȅ�s���!�Ju	���s��|�z��q��:�9ߒ׈���s�������Z�!�1��ue`��Y�Ψ�ם�����m6MT�ǀt�������g�r���8└���F�@`ўؽ�ފ��<�~�s�A�$Թ��=�E
��]z���*3�W���$� ֮�O[�W���Ҍh��I�h�N��r̍܎2.m�'���!K�W���T���%�l��Nrpz�����\�vN�{o�EL4��1��ڈ%H{�"��n����Dl�A|�@}:/<�j�E�Ԙ����av�y+v�����!�]���T[Uqaf�W{M}E�h�J�b�� �Z��q����#��{�t
�?�`8�3��T�mk�!�J�/^�jd*�P���Y=r����=8	�V<�ek��.���,]b�R	���3���1��0�?}�dMű����N�-�F`��ߢ�5 I~naO�F�.��,�^�VZҟ�_O~x�6�vk�=�`�:'M��F�g���t����(�:�OJ&�al������/f��.Z��u'��''O8�,�$=�G_�����-��-���$��~�`g����o�W���f�kv,��L[Sߐ<��.�u<b�j���2�&C���s\����j�>�fl=5/]ܿ1���ٓ�o���~�������>>���s+#P�#`���[�P��Ԉ!<�t➻v�o��_��,?����G�V���_�������^�� ��g/ڧ���;o��ݝ�}���ϯ��n�#*�RBbP�M�w���W��g�v�������7��e����e�$�G~F�BM'�[Fp5$6�QQ�������|��W�t_�}��cW
v�rݾ��m{���Ͽ�����[/a�.�ѩ25E��2c9�E�7,S`��
��4($�x�_:�[yG�X�1��]ʟ?c�L3ev|hFAs�T�#�����Y	8��/*8����_;�ܠ02��cI\���_[�ϒ&q)��N��Z5��*�>Ji����*_?�CACp�M@`���z���\�/�{�'wK�F	�A6"�Y���H�;��ܐ�������z�����Ǡ�� iKoŘ��&�mCY��Df��x��2 �F��� =J��3���m[�C������^�1d�V
:�-��ZR��l�4�\�����?\(��ΝU���~��`�J����ސ	ݩ��k˺R��JR~��������RN�)��M�,`��di��{�A~�ڣ=Ow*r�oW�--i���6��9��*���?�Jn�?W����h8�V�Eӭ�D�q*�TZ�J�Ae:hp��k�Uz�[�U�h���d�83�7ױo��� t�4�����6�a:�k�{Ғ�7$7�C@@T��g0⛣Tfh�0���#�zIC@��l�p�ו�ֵ�c�2b�a�|'�Q��,��U����%P�`4`_�c5�Wq���՜�> (��Q�C�����l�T��MנzN�C�gT[�'*���	0��`��_ۧ(oz���1濕���fe�Gf_���� "�=
�N���i���dX!��nZO8c�o/:a��`(e��Q��:q�&��<_��N�%�
9W��IӬ�S3��	����{��.Y�|~K����Ԫ˒��{�28���ע��c#3q�K�j�L��u;�l� ��8��ȧ���G�MC�8����vM���pe�ضA}��`y�2��Gpಡ /޹��=��V0a�3d4[�U\���/���oWݭ�f�����Z�B�|��W�f9l[`-���s�y�+)#X¸`Sa<���M�W3�+��D֨;r�0��"w��k�F�����[Żjfe�Ue����0�"��M�HΊ�Jv24�]#����/K(z���3H��_��Z�E�4tx�(:�@����y��a�a��T!l�O>�pd�~pY��Ef:���c-_g�q�\=öEp�ko5�#i�Ҫ��m�b�%8����^��9W��Y��o
��y��������KЍ�:�p��( 60�A�P���8�d�:�ab���>r�2P�ñ/`�+4����yyA�nl�˚Q��jE������}�=+k��-�l>1*�%�S_?�$��]-#:Zę>�_�mCGl���;`�Zb2���ʙ#dU=U����Q��f1��1嬾Ƭ��Ȩ���\�ߴ����e�����:Q��_��Ĳ�ˌ�:�y֍T��1�5 �i�K����o��
Z��o��J >Wx��|&j��9u��EE|�et����Ԃ� �$}�l���v����1U���嫔������
�Yu�R�3�cΕ��� ޓ�RVh	�>Ӑ�E\v]�1+�6=��kԱj5<��vu:k<;�	���ºת~q*6ȟ]������g�~o����~�6�����k�:�jpu�b�9�Hh�ޢ�=G���({H^UD"y�%MM���M��h�E�/�}i�����_���v�6�����t�
����5��:<�؄:��Q��/�P�[T�������2�4�`/����_������O~�������Ĥ�H�3�!�Y�'����O=�������x�3� �ݿ�_�?^�� ��~�\Z{���_=���g^=v��.K��O����pH��q��yW���[_�yd���~��{����,uM�c�ƃ`e�\*,�dÑЅ�;D���I����ԄM�.�%<}�a){"?��{����o����?���a�  ����g���Y}-�^y
�2_�E��{ԬE+Ύ�赣A��DװF��K��F�v~��9�;np'A���
��������&�J��Q ���-f>�gUa`��oEZӸc*!#3�\}&��̆	�d+�	������w�-���F͹�����f��l���&)^$P)K�$X���/B����=�'zI �I90�N[�b˖e*�LɲDE�H6[;�>g�5�2�������-*H��� ��k�5gըQc|�Z� J��.�GK��7�
��x�]��ޱRP�1gz�|�����G;m�%�P���eM��UZ4�8��jFƳ�c?�֘ �Je��l]2L3�2҇gCC	7*Xf�l��,`�VY
��߶�s@�|RX��sЮr�i���B��d��}���H  ٌg���cVe�a�'��:��:Φ��]c��C�}d�N�I��!�Ffa'��3�#�lM�R=�R-^
[v��W��X�1׃O�sg�^��z�{����<����9��P�A��
^J]��$o�j��Ng�?�P[קC"��h�����	1Z���a�����|�q�Ai�1� �xo�9��"��B�s�V�p�B)�N�B���J@��~�:�{�H L>Yu�g4�]����$/8�]��ᘼS�.8�uT�m��F J��&M|��|\kYQ����|o�1C�&�ʠ��{Y����A��Lg3� =���q<?� ���Z���W���D[�x����ҡ纨���'���k����#�i�h+�����2��K`j�0p�����N�9�D�a�vO�=�
�VT��I�'*7�Xj8>'+����d�>ά���O��G�Ur�伂*�t6&�*�9��������a���/�	�x]4`��8�5`ПXR� ���1i�s�w�W�-��۟����|_̕qŅi�ʉ�z�*t�"�C��2E��N��|`�;J)�b{ps����<�cJ�Hԕ�)�v�@����W�.�=�t��QV&�0�����}��	�8�M���j��{0��{�s�t���ג��?�+�$,#�4�6<���K�Gr��%�?���P҂�uY!O�fl=���cnH�.�f���n��FEK~�U3WG���y��á�V�m�V?dd�H�>�@b� `��x��[пF�h������ݜt� e=ca�%�S�h�lj�W�^]y|A����N�� �%��d�A��X�t��W��CC?Śg���I�'��z����2������Ao�(�.�Ҥ+���#q��<����'�s�x|�J���v@���XrH#�U[$��F�ڴ��J�{��L��w�SF����I��%�#�H�"I�W#)��d����E��8F|���V�~���/`��9#�;e��PA��s�fW���<�������4�do���@F����`���D�!��H9CYK@�r��N^��������<@;��U�|Ϥ��$�3?��6O6 �z���/D�Q��蔐��8IK�1��"�ǰ�ځQ`�Jb:^�d=�7���v#��]���D $�kg ��ƺ�h�B��V��/+���@��u@b���}�c��GR��c_9��..YE�%oq�G�\�[�gb	������ᗒ�ׇ'�<����d�Р!��ޫk�c\ 8�)�� 9���ʙ��so�M�q�4�w�&�-��{�����Z/�,v�.��z�>���G'�޽����]��&��dR�S@�(#���}���"�4�ts��?�L��ё#���������g���]���ʟ}��#����iXsK^�L�Ze=�Aۃ=|��~�Ⱦ'Wv���5;Yԛ�溹n����O���፷�x�W�ٯ?�޻�����#�C8��.��F�7w�/� �
��lo�{����/������8��@f�K�x�
h��B� �y�"?�`��7�o�ݽ��I@g�`g`���}Q ���x�Y�K�x�+�j/�~�~����?��/��p����hi@yÙ� �̌��J��R�tpe&��`&s����3�9��j��&1�ɽ�;L;(�@m�*<���!����U��<w
@@��N�������"�sh������%:�0ATw�!K�ԟ>��` �[�0�F�A��:��Jdo�6�-:��UVͪ�IұVPs�b�N FV&sh�pa۴�~<mY�	��qCN�r�Nڝ@~ΟWm��c����������!+�xr�#��L��{t�.
��}	�b����V� �< "!`u>%a5��1�%�ۄљY��ђ��s�!A[���Zo0<N�۷��'�EI �_N	���8�<�w�qd���^L��)� ��X��
%_�A�����w�@��CA�?���5�qƬ��Lg�0�F�6�kT���
�rjY?:�H	Ƨ�5��|ȣ�U�1��~w��p����I�����}݆���@�U?wv��i�o�� 3+�����_�"��#B����#�
kgIk�?k�����.	�c[�/�e��hWn ��F ���{)G�V�K��p�!*U���s���g "�t'�L�/�~��g��î?�ߢb�Av�0��Eh��I̤�C����'��@��I�k��MF�>ƃ#f�ڀ�� g~5����mN8C�Z��R}�I]��_C�B�Ȣ
��gޚ1�?��bܿ�{N�L���0�Et�����y���A8�1f���8�o�M����/����(3���P8cMJb�����agg�s��D0ӃCOŘ��G�XVwC���SN�����&�q=����V&�S��yL%eH!�iī���~A�1�-�MH�Q�#��5(A���bf�U��M�EE�hL��Ӛ�WM��{��<�����e���H���0R7c'j��{&�څ���h�l�S~�X�������b�|�	б�L���_��x%A�^ݚ���Oȯ�� ������&Q{Qu����l���L�J�1�%d��*��		}Mko�$'.�	8��~81.��"�&�aà��C/���6�N�'<��?���X���[���ÙA[Y_v.��'P[I<V��}��9<�7��H�����ʇX�-���ޑ��e56u�pk�b���;8�0��q�Ax�K�P_�R28ͷq��SL�0������ؐЛ=�v/π=����vuuG�qT>��W[��<��c�y��CҀc�͏�j�W��dl�:��i�����@�	�c+�׷HL�:|h%žA�4��%%Zp���53B��TĲ���s��L
%tܐ�Rl+T�x�|g���ԏ��	��W��"�{|��P $��6��Z��R�~�r���1������X�1���tJ���S�(p��$
B_��M�+A�GބsM�����~Az�P]�罥�$�O�ФR�u`���)��x�	T<���g�|)2�{3������E�M~/况�t1���1��w3py�;|�6v�v��E���F�����.���Q�8:2��>�H�Xbi����O���vzT�H����p�[�a|H�)L>+|�8�ɍ�������a�������9e���;������W���z��/�N88���o&��ɿ9�gE�O���2��������j����Y[M����ʹ�K�C[��XN������-/���-n�	 K�m�w���[c�twR0E����C��,�oŢstG%O9�p_}�8:N,��F���}O.gC/����	���C��;�ڃ���X��K�<Z\�暆����z׼�&o_����7�ϳ���?+�;;ys�\7����\�k@s/ٲ+���������;��2�x�]K`pw2�2�������~����[�qW������W칻��J��� y+,W�bA��ψv2P��L�V`&�[d�0��&�;"�@l�Ȗn\u �V�5��R�%�d�7e��I ��Һ+��ݷ{�U����5{��x�r�*�^k�
i�J���0=�7Al	d��
.4�
[л]��5+��J��E�Р����+Uu��U"�U�c_��ږɳ��ZVxf�-�RZ��
8�J@P��!�0���	� R=˾Ol�3�p	^ق�Zp..��} ���1:�PC��e��Z&Ռl3Ygm=%�59K��k�%��)�^����aЦ�٥$�t9P|���sɁeVqm��j��cBK��Hn9���x���L
2�%+eB.�V�*��oZ���5�R� ��Ĩ�ͱ9]����2���d`s	N3�3	��M��F��� �����cah:xM�G�V�
߁d�D�>>=�<�!n�#��7u�k��A�1h�W�`�� on�y?~/�)���3ka!��VO�HM�F1Z �aԢ��	I|A���{8k���1�*m�[&|�=���L�ǽ��8�^�(���0\r2X����������������&~�}'�����+-����  ����z�¡_3�16_V� �?�PQ�g� t|ƾ�a��؇^	$kY��:�!2)��:����n���;��|��Y�.�?X�3f����8=�����F�#g�����Ι�/w$��l��8brzS]':�ϑnFg�y%\��d[ն�e��!��k�d�+�SH(��X�D����*�q܀'�,�Ʌ�b��%��I�pڳ�Z�.^ ����kR�*p���Z�Z���.��P��^�CS�[ڭXר����7Sy�|�σ3;�>���T&<�3��5?6�?� Kt,� 3��u�1�����ٿ�4&8փ'ٍ,���3&��zr�bv��!�נ��xl�G4T ��6�Z����.S˚6��{ �ȳ(�|����q�7x��y	=F>=��M�LȜ�"v�֤�)�(��dK=XqjẓNxn1�`p�v�Q��b'��tL�!��Ka#�6H|��%��7֓JAKy�q�sqӣ�T�ϣ]�vd����|��Ʈ]B��� .�`�M<�x��ř(�/=J��\R�:O�yrc�L],��`o�e4�F��饺��f']i�ށ'�?��vɷ��,��n��_�Eb��^4X
r<��˺ξ�V�Q.��?�Dj�����<�����vt8\!?���3fK= r��������,L>Z��l�"8bef���(�~&�2O�4Ɓ����e��@�Df�����7�̈{Nm\`-�� Av ��ޛ�_�/2��G���J�Z�$[��zɻ�3�Nq490������3Ua)L|p]�{ı���c�����<�'� "^v}�x��E�A�S
ֲ&�s�*d�QY�z�94�[(a�bӚ��� ��g�@{����im����"|�2�`�?��0.��v���
ͫ��w�S�5c�v:R���ԕ���sd���|�#
�=�k7�b���3�l:I�� �>�%e+�¯A��ݛ�?1�_v��Au<b��'@��_�[����� �����5[�ލd�G���F�W�6�k>E�����D�!�z�:,Y+�ac�2q=�_�p�P�PcoI��;�����H@�y����nV��L{�����J>��s�e�X���A��"|�$!	(ך�̜?P<�uh8�bH�?}��K%p��*m�^[�Ha��1�F0Z��U����m4b��z�XI�d&�<rOF��)���S}}_b_9v���z��Lc�̉��!+q�^� �͋���d��N������3�c.{�~�ե�jgv~v���}�՗m�1��z1�}��ٱ]�@�x[$�mt�^ ؏��cy�m�è�����q����Λ�;Ԕ�>��i#	�˦������x������Y������s��?.���?n��G_�?|�m�+-��3.������B~Gs����{�����W?��������r��}�ܽw�^'�f7��us�\��~w �"l�ƣ���֟�ۗ_?���C�z�؎˲K�"���$in�,Gwt�����8ڳvn��������l}xgŴ��l�@�8sxx�vvC1�⎴���b�ퟟ��J:��ߢª�7��;}����ہ����A�>G8M� �Hi4��]m����S�?~�M���ٱ;{:Mz�R�*�]�� !����,�>��@:��e)�R�-��[::�np\�QHGR˪���@ژ��_���Yt���si���t80�Vaxef.x�+��� �FRs�p���t�u�B���W:H��5�3�b�j��T+|�;�6c.H��� m�	�F���XiC4 ���C=x�\] ��/j ��
�N�Y�ܣ�(&$��Е@��V_��'��Y#ZB�ƹ��Z��f7:`��:���KGC�������`�U�zn�1(���- �����@����:%���m�aߑ?�F;�FU҆��h��n:$��)�C(���\��ʉú�����!*Q�>�+k8�+yS���!V�%�A��{�0�Hp�Z��w8i�_���@ȧ#�~T�p]������]�d���Ou�W��:��7�ǸFw�l[�Ak"�38�r���?f�}���l�/�xy�K���s��e�o���v�ř�Fq�$	��Ft���P�D��V8V܉�x���
8ƅ�:O��\I;U=�8-M;d$��!��֠�;~�p�q ����q���������7TU��U_#?�s�����,���WwRb��C�b�E�dY��QYПQQe���s�j�>w�����Pbゼ�	9aF@^M�3~Z�
<�D�EqO�n)���XJV�!������{��2>'Od�M��9�Y�x�%��{���;�zl =`��C�#aW*|�D�z����ߵxР8���rf���	�L<�c&	X˄;.�`��C������L�-�[�i��ej�,+���c���u�5��;P�=�
�e�;�H�Tf2w\'�ِ��6�Lgb6S~@ `sSY��������^����\��n�sW���T;�K~�]$�&�~r��,:x"o1&�œg��ȱ?ʪX0L<��e��n����
;ҝ�^_S`��jH�8|��U#Y�I۱��]2�{��j�Q��q��ٹ��)�G\�'�@W$���d·`��^dI�?U��	݃fC �߿r�C�m����N<���n/D�eҐpR�S��9�!���g=0;gCpGO{+��	��Jw<���kK����-��rB���nK)���2�-�����4=�H���`w�隝f���^�E�k�=�� �R#��Q��F~�<�X�$P�ɇ#}m�䐯Xcʽ�!�	c�O�0��n���#h��yD��Z�I�����zwqv�$|�)F[X �UХ9P��"��ج�	9���Jmǲyo����L��L0%���ecb���8>Ao��D�G����/-��D�y��Q J�����������@�63_�-d|��s�A�9��8�>���Aۣ��+Ȁo�O�P]�k�&��I�4�o��Ɔ�E���j]"q`]xtI���&��Y8 {�,&���)��}�O�1�$Y<?��%i)�2i� IxLY8���ې�`��Nq< ;)�{��N���9'ϳ�����y���Ϲ��e⯺��˃��I�},�ٵX&(���Q|��RA���,��������~�S�'u�&{�
��v��\mީ[x����8����]����,v��;���������ě){f�IZ�ܧ�3H��oh¦�� <��X(T�����������;�ī?`wǗV;^mv��7�܋kʖH�7�o���_�򼌲RO~i�r`�c5��	����޷˱�r����Ov۟�c@W6b:r�-�{҂"��{������A�#���'��׾l�գ=�{���̎ɏ������N���!����I^�����^���/<��S��=��;�-o��ݗ���7��us�\�z� ��;��r�n}�^Y�{v��;ڶ�[������a �
�����k���j������ĳvvن\^����0+q>w�m��m����M|Wng��� �h�:�g�����ԟ]z�^߻�/^� m�v��Z���9��h0�`��po�t���'>�	{�k�ڿ;��+w���`��eXk$�|G|?����;�mL@��a��0�`�0㲉�h	2>w<p�>L�CX�b�C��aN��� I�^�h�b�\g�>o �H~h�ѺD�e�s2��5��<����+}���5 �%��N�+{���ܸ�6M�:Ǡy���p:�1�&�Op���_��.�тF0N� �cG��g�wR��:G�cdTzZI��M5#���ӯ5��0���LtA{9��Y�cm���~��s�I�W�e�k��>-�f�Q����4&�(�S��(�O���k>�� �
�p"i�X�5�hA)r-[I�vb�@|��B�VL��������i����D䒁tЈ�%Ҹ��w]=����Y���xKV��'V�`8�x�$�]�z�J�6����	��7�l8q����.�ς����ם,^Q�y)�x��{�	����S�f��䤜��@p>[̆X����E.��!�Q�ÂoC{���X��Uf&t�>�Wk���5�tDvT�/�+�[�+��y����rBw�8΢e![����=*���������۽�d	�����p��X��>P;0��̗����5�aw�p�/�h�i�"W��R�"p�>aK�H������a�,sR�;!�fXm��YEeM��8=��kGz���GT�8e���L�Hf�*V΋�6�Yb5�����evP��lp� Z8&����,��~� [�!���;��$����ć�����'���bfg:�8Gb���^�#%X-�tG���j�Q���� ��� ��Z3i��-��C�3n�1Qcsq�ٹF��
-�L�\ރ�'!��Ԙ�>��Kz?�e3��{���)ן�'-3��͟�]ŰR�k=U]c���� �I��u)�@_~mz�Y�Q>/u�Q_��c�Ĥ>I*K'�;Tt4���Ú�����%�1�Ÿ�O�x�2+vA�5�x�WI�!g��X( g�b���h�ڢ�+�O��0T�[f�
+i�S׌X�\�m%	�%�w�½�J{�roZZ˖��;|�b`$�.�M[�SG:����Q�!��&�T$x:��i�3�%�6DL����R�V$��@:ưj�Tg,q��,�`؀�MpP��8���k�N���i8�����?��&��i����*�#���6� �y5c�M�~�I��1���;O1�Xv'�	�#�����ydZ(|�Q��Q���oFN9l2�{XZmk%j��
q7��>-�����=^5�ְct9Ǟ܂⡘��H���NQ��4�M��;;�ɤSs�����6�f�Y輂�"Xu��2�E����H*��`�H���ڱ�0��8����˕c������cૣ��~*ه ��V�+���LvA��,T�pAg�a�[s0��f��S��ڴ���M���D�vY��2�ApC��� � �^�Z��v>�.ű���s�;M�-y6��lϯ��S)���A�c�hs�wU\�F�?#A(:!�tQ_��}_e�ƂV��U�Ԧ8�2}&��.��/�l��d�#yt��z�S�qF����DҼ5�]�G��jK���|��|\�d,�5�[�]䬬�'�T�"�S�u9�+��(/;뱜� �Ǵ5�uh����lϔ�QE�eEo��}m6�)tՁ�-�؞��X����/���?�g�ȓ�	r�]�g���ѹ�Iu�u�d��<�xK��ۆ����>�>��%�j�l;��?�Q�կ�g@�e����jٻ��"t��:�V�}����r�o=8��޸���7����ۿ��\7��us}��}O 8;{m}��o��^׻g��w�z�Z��H��zV�������k��s���ݏ�;���_���]X�|�A��� <��؎�;������,��F��rk��|慝�?f���og����':��ʲ]=��ˇ����xճƎv8X���>��������>׮�A�Ko�c�����< <��h#�l����x�{����{�+��_�׿�e�NoW��s��52��{��I�+�U�	�i<}�:Y¹~p��A+��6z�Ǥ�Ӑ5�� C�G(�+[G�����/A��T#��`;W���>���*�,̳k�*�$բ�)x5�	��/���H=��4=1�����I�F���5������M kJ 5�d��wJ*~�t���ײ��2L��q�3���&����}M�k� ��;Y��&�ɱi�;�[�G��_�`�����;儿��׌��7Ļ��p�g��R�k��]���4���ЀF���]��K��>��g<߰�@{i�.m�=���>���8 J0�-�F��`Gv�� ���c5���-rr����"$��~,�O�b����=�d�78YZP-�G[����8� �@[=�3�f�V����}�t�*���E���g���X����D �Q-�!�E��ָ|���<�/yhcXJ�w��V��Y0F|������ܖ/�*��`��|�����$m��G�i���?��/��cW
�^}7E������v�_�����"Q*���+��^U>�c6��-e���%�Z��R��2�j�н���Y����ލ��9�#2z����{6U�5q~�<��,����N��R�q�Ȏ#b��½?�x<Ge ��2wg��A�s�LsLGb������w��T@ƲZ3&�A�Ӂ�,�=�k�-p�,jy4й�d�����z�u��x�ђ��S�8ˏF~Rr~�3uD�xz��_�=�-��Y��~��k�o^)������'&z�������#U,��P�D��aXf݃wg��7��tOQ&�,�h��ԏ=����%�	�H�Uړ.˼�-`6�A�$C�D��	��v*π?M�k�3~)��Mҵ_��.��F��+��k��&�4�V#OJ�X�RE�����I�����b!�+f��`��{�=ǦG�;+Ԋq_ňy����Wk&I�y�w�vQ>$�Ȓ��LG��l��sƋ��v���H����l��N�y͔�Okm��N�ך�kRP��)GKV~.��P�j�<x�G�5,�|�� ��B[�8������VcY2�D�;�9^����	Mh�{����pʣs�D��I?H��d̣l��a�gb�q�����ȃE���Y�3}�쳠�/{cn_�e�w0����<q��d��g��
|X�$�Q�ip�D���i <�+{�m$]���޴�#IC���E<П�e���s�Ȟa��o��q�_Xm=��<��u��1|eN�B2�~C�0d����2�'t'^�-�7�T�=s��/3FA�,���$$���f�?�R���ﰹ���_�]B��N������h�qK&?PU��r�+d�QǵQS{UuT��"z�Ś*�E�W͂��t�Ϭ-U'���lE":ؐz�ۓ�]M�l���c��4�I&K��XQ1Q&���@����9�)	�z�G$X-�{R[C�$�LZ�(�I5cA�dc)@j�cƾ��z�ٲP���I62�'�7bb1��*q����Y-:bO����I����?��2���t�z����k�O>���|����.{q�я*�e�{x�AK�˃qLc�/g����߽p��N�s�s�ݺs���λ�1��K�z�ЎWl=hm{��ȶ㣱��vo�'j^L�c:L�c�������\{\��ޑp��cw��7�y��ŷ��./�8T���;�l�����^�>��x�ˣ�j]�...n߹��z������us�\���o!ўy���o<y���'������m�í��r��]إ��f� He�`��t!y������������YU�,�h��YeF.��4~���'3��<�H�z{���-�=����Ͻ�^��K��3h���������{�[�*���?.�}����?+��R���U{��Z\hCx���d�Q�j �%�}�z����O�>���ڛ��۽ʱ����j�� ?�S�"�K��)��#�!���N�_��79fQ��j%�s�|	���ۻ�fɪ����� �q��9pZ���Sc)LBA���.�X�����H�k-l���s�œ����?�.8绐h�A���ɀ�hX�%c�cu��8�4M�� ���7�R8��J��@�0Da\�R=�B�i2��2@�,N^%*��x��]��m��[O/���9��t�����敥6ڲ�tw�s,54 ��h��4�Y��Mx�at���Z� ���sd� �ƫM ��iG.j�d0j��P��h+�t�o�uF{k�I8OZ:��]H]T�����B�bO���b��I��0�`����@Dk?�>Yb�N�*�+��]ޜ�74Ztj������;t��X!��T����$?Rs�p�������ǡ7�h�1j�xgu��i��}z��rY�fl�����V�Q�@���k�����S�P��nDEg��F�O��e:OV��� '�0Q��U2��D8r���6H��V�fwg����s����s��U���Z�Y ��x�3]�u�������}^q��Ѫ{���7O�YqT��px%�-ϧ��B�'ԝ�"��.҄�6��~�b9���?KR���Y�8��b�!��UB:���|1�ķ�o�9�%�P��M�i��X���}a���A�ªI��L�r�e��Rň��=���-`A�!S���tH�2Oށn�[�b��q��D\-Ƥ	-p%h�q����k�!�5Wv�Z������o�J;:x[~O�e�VY�/삨�5�|�u�J�9���{"[cc�w����NO<\҆P��V���1?��s�O���ջ�5�J�����l�0�D���X�������/f�EufK�7����COV����].���gC2'�@fܯ�+O�Ү'�YȞ��)�,���8ms�F)�6W���jw�%�׊4�N�N:^�۞��@�� )�Rs|dG�Rr��b�k�<�#��2��_���5���'�3��B7�! \&>����`�y��l�O,��'A�Ȉ$O3Y_tb[�&��/�����؁�6#uU��kg"�Ay�(/��,�Ten![�T[/RG/�@����|k=UltDژ���C��F����q\�:���A��ԕGjPĘ��p��0g0���v����X6��7Ǡ?,e��K���9��]�l�oz
䆭)"�Կ�2q	��9Q����ކ�B���Kb>̣�z(��6���F�Ds�9���l��>'�+����C���O���b����6"���5|�㋿[v�;Q��z&��n�K�Wډf�I�"�Ӡ�C�C7W*�|���q��	
~^:�X��^��9��G���߃a���C	��f���Avl������{�t��Ģs��0��D]�H��HYt�m�j��FU#ѧ��K;��=:�|��!u�7��� 9���½��*%���gu�/�j���ϱ�~��t�P>#1���G2��$��7��mH&���X�x��~����Fu>���0�+����<Vs�[�k�<�bT�tl �b�$��d$��n�Ɏ��~�r��pȨ�����}��٭����P�ץMiH���9�5��_�u,㈓]~�r����={��ٳ�������{��.�Sf�C/���Ⴧ�ƛo���S{�Ͼi�y�=��N�^>�o�4I@�ԍ�h�9-h�m�����9cГ �v����O?o�x��}ޗ���Ө��.�떺�����S�}��^���zk��>v��W>�n]ׇf���us�\7�������ۧ^�����ş}�_�����уc�8�V�\q�z~u��>�~>ʭ������}׎��l-�4��I��Ma�^���Y,�1y8ۿ[�������}�����O�ԗ��Ǟ��z�c���9��?��r�\����?Q>��+���_�N��W�Z���M9��U./_oe�jo{s5��x�٫�a��5����Q5���:P�쇟��}��߶��b������](rg������B*�Y�lm�V���j��	E(F����8`i]с�f�-�]"ڊ�%8A:ϕ����-�"����< �<)��u�~Φ��u�7+4a���� �Y$54���[�2�#4`��y���3�z��M8��b�⼖��(ۦ���4H�s�����"�X�#�5�nc�a�� �N/�DWp���h&-�XH�k9wӤ�tR8�ۘ��jT�.j1�n��#`��y˟��5Z��խ!�XE�؛Ė����A�L2��9�OO���&���Ʋoi E�����|�
�1�0�U��'�ø�7h[z�-�RSp�8�����@���9�N���IzB��Yb���9�����G���o@�t�lɣh��5�'�5��s�Lvw�)�|�7�`��w�����E[�-�OA��bw��K�ӱ��[Tmq$�<��w�1��-v�En�q�$'�UY��䖞܀�;�%���!���q_��#�"2�[�Օ�ü�R��g*�f�m�~=�`j�-8����Ǿ4�'��b�P��_JUoEK���P�A�h�N��g.��c�pf�F�E9��ؑ8֍�Y�;���Mn�<RҦ�	�x��t荐�uVC� ��r)*-�6[|c�F��պ_�p��:�a�N���!��� .�� �E K���� �,�ӢY�E8���pV�� <�4/�F�w���F=��nIy�h�NP�x�fe��}§U�pX垔6�pfY�a��SG4;&I0�t��ѝW:�}|pl�c�E�����=V���;9�ۘ@���F�˥e�x�Y]��ɫ��@7V��C���ʧ]����=�f�"�*�G@���@��{5��tG�Ѯ�*T�����3t-�9����+��!�f��Dc�7�3u/��Xw�~�<�E�h�~ɗ��ٕrb��<,��G����	�$emCR�L{��?����7��{���b#`�X5�3v�����J��b����H Y&eݓ�0�X���mF2�vj�@$�����d�#`[��[kْ!'@�ư-�^�w�9DE*dc����kؾ!�������+	�Ff�xY�J*e�[������6��s@�d��\&������	�%�ԥ�ݢ|�O���܆]M�|̥���d� (� 涎��N��_i����Ϊ�-|��Q�KׂfS@i��N�N`5ʀ�9C Vb�cm�� )u��_�\������j
�{� �Q��Z�>�������+T�� ���e�b-�-Bx�I@v�@�Nx;$�H�vD�s&=dW��[¬c���	t���(��2p�ղbGO:�]�����1nȯ\�m���͠�1��N<��$8f�K����;���(]8�F�����!�Y��Ǖ�8�Gkur���h�5�"���oV��/Uk�+�ߒ��~��ir�ol�<�R65�֧Q�g纴����f&�ϫ�<H��Y�{c�'�&�����\���W�Yt?��	�p9o\j���3ǜt�<N�uB&�$����a�O2�Q�䞮����S��t�>XD>Os)���\���,�p4�ߛ� ��o'4:ѧ�W��C��h�̋{��n4�k��{���`?��W��¶����N����{�7�.�4�&	8+T���e���a}�^~��3��!��}k�|�d�LH��=���Žs{���^����o�7�����+���~{{��;�w����ut_"az@/Dm!���_�D���.�>��G�����=����_\��dM��v֮��������~��?��'���y��'�����I ��n���/���$ <����}��_���ç��/��Oճ���.�����E92���p����-����8�����<�T[��#��zd�g�j�|���ҳ�.����.���x�^����k�Ǟl��.�Vֵ�R27�]�������8�
wm�<��=��3�������W~��ſ�_���G��=`P=���	x���< ��$?s�0��E9�^������=;����Q ]��c�4>1
 ��oP����m:�
��X;���� /Z�-o���p$���q���'i1J�Ip���p��2�h�TVd���4& zx�9 ���3������t1�2C�B<N{��p��A��4��J�a���y�~�i\������4X-�h�yA �`�!S6�D@rTɡ�2�s����٨S0���3� ��V�&�a	#��ּ�R�Y����ں1����f��F�>�#m݄Ύ�'�"�`+q���,��k:W vu&��f���W��,��������s�ܿ¶��{�&O�V'xޔ{��;�|
��K:����,����5C���U�%3�;UL���2�k4�c�������QUY�xI�{��47�r�6�k9�KΆ����y��'�QŰ�J�c���8��4��,��jV��U���5�����mt&x҄����&�K:M�L�
j8�P�ޓ�S�S���p����a�D=+�ٱ�a�}�q4���+K�G�T��dPy�4�O��v��@F�E�9���.�W|�;���ӟ�׭����=*���|���V��X��;:,c�I��@n�\h�W'�^��t Gb�1�sj5�����J]�SL� �������-����,�j��}��i��Y&E��yr�,��N*uR��0O�St�(����Ð�EZ�ʽp޵p:$N���,c��?�yy{�2��$��i�bqx�0��&3�
����1� �Fa�_��-[u���+2�oI'����ԫ�@^1A3�CW 55`�<��!k�6>�j�9��U�s�f�����(g���'t�]N�]��*�ϻ??	C~Ώ�9��N�����Ʃ4I��y��7��صLvC��v$0`�u}���!��-WUDjr���Q���ٚ>�=�5ȼ���X#�\����	���OiI���;�M��odE:�Ɲ�ى���aS�<�뢪.�9-��O:��+_yCG :���Oc,�=t���-Iv��{J�Є�k�"2��2� ���G�����r!x��ʴ�&I���Ԗ�=�>�ROV���;0,��:�I,�gVǘ��nf������aWx�d�z���:4O�>��H0��� 	��cZ��N*89wY��Uv�( I���Iʷ*?��3=����w�܊��xA&%��y�ѓV-��i�~���	�B�L$}Xt:h҆,D ��FG7�]�e1��	��{�'� j�1t���de���el�FB�AǞ^�0�b3�/b���)]0Eʊ�sL��@�3��%��������Z��gR*�Y�i/#?Ǖ���������`0���us݇�X�۠��dި.9�ø�aG���Ο��ˮ�ۡwve��D��E��v�;p.|	��a�{�N�m���'%�GM=H����=�$�Q�x�P)�+��B2Fb2�
�fq���<M�źC�U�_�o�`���w��y큇N/�9���I~N���{��S����݃��t:+be��9��î��YʽP�u��J�%���)Z�6��������9n���{�yk	��i{���]�|h�e/޹k�Q�G��7�H�#捾;��>�8ZҼ�W���b���~��g�>�cv���H�^ N/�eX�~"ۡ?::Z�vq�)�������}Ҿ���~�7��ߵ���}l�l9��1OC�B����x��3^���������=m�o�[��G��ߑm0dA�с��DX��]�^��_�[o=v���|�l�9��:�Rދ�o���溹���& t�_�;��ycy�֗�K?s��|��}�r��+ۣ�Ȣ�� ��� �ad�v)�e�zu��}�U;^=�b���[ͦ��h�3gӸ�2�P�=��������9o��اۧ>���֝;m7��W��w��n��9���'Ӆ�U�k�[�]�h{��Wʯ��_܍�ޞ�]~�|��������4����.w�x��ٶ�է����[����) �`�-8g=[���W��ͦxO�q��9Z�����xH��̖�|��X9@|��MO��*�Y�A�ĺ6W!�B@�B:�4�8LgW���C�.G��ĸI�'�B�� ��nB�O�VI��d�T��b�~pK#:x}k8�Г^�8>'�MG�?W!<(�V�L9��!H-jTUC�&!��4��:���4̒>��}]{�Ƿxo�u��SK#�n�!������.�[���S�1Y5�X�X�|���"���u�@o5>�����[K��(ޅ�E���30k�����Jc8#ib��V�L/���w��|�|��1�%���kI�(ά���0j��N�c�E�߃9&<W��#S�d�F�>���;��,s��3���rk�5�q�UW�@���b�u�bѢ}��7�L|�ڑ�r�k��&�i��<��Ҙ-��4�Fs�İ�sr�Y�����ޝ!�	��y��
d�B�U�u�m����32F�����wC��'�A>�&ܢ�_�/pM�x�N�Q�6:���z���I���Q"��F@�n�/�ѫ����������`����,�7����C�e�$I�x�t} >�L��n���X 8wO�K��18ȳ+�h��C�*��3;���XȏJ���=���a��Y#-����\T�eh��9�X����A�	���fT���ژB'e���!U��b�7��|����$�T�l��1@��� �I����������du�����ۧ2W6��3�7+(�=sP(�Nqx�!�9�;���W��s	�M��X�g`ܤ���0�LX`�l��|���m�*U�B�\ȓ+�������׭�_�l:Fy��t;S��kY�~$ڵ��3�l���SCNB���uNm;���y*U40��K��e� �!��g�^&K��m�7�ؑ�����O��r-������f�^os��V�*�ۧf�^$Y�
|o�Ķ�I��s�,`��P��M��7�ؿ#��b�_���W��P�H��+;��!��=>���8���>��5,U������<�V�uu�k�� D ����D��h�^+�c,&���.�XO���Ur�cH�g@(h鉨�I֍�t�|+TC<L.�s\_�@d7�@�K,쀸O�.;����� g��E����&y�{9eu��2����v�q~����<H���rXW�ȴk3�f�}���]�̲�<�?�Oh���7H�֣Fl�[������q$[�sML@.5��|a���8Z�ՙ��7`�@���n�`�6;W[b��l�@��f׽&�w��AG,���I1����tn�&�(e>�YJ�{)��2��W2�Se<�8m�Mq2��=7'`���y�wT�s���Ic9�(�.�|6�mT�y�A�Xh�f���̓�tyM � ��N2���ˍ�&1�XI;_*ؖ���3h�:�{�hC��nM|p"�����x�q?��[&�a�\�5Y���@]7��h�_������R,���?׈�k)��f|>"h�ƿ7���)�s�ʟ���y�W#^����{$��Vȑe$���z�#��16�m��Z�V���@������.BBp�&��H��H����|EL�����>�z�U[]��m��v6��}ԇv�h~&7�'�����g;N�m���}�Gʞy�Cv8��h],t��������<���t�z���^�'�|Ҿ�����W�t�vuy��s��S�=>��^��|��zm�q͟��K����k{�߻xk��{|7dB����o>��{�xsY��loܾ}���/G��n�����������'���������n�5�n����\6q�*����]���{ݕ���>n�u���X1F��5G W՟�2����ڕƓ���+�#{��
���a���= ��������5�`;p�k�m���'>�����9��_�_���X��.��p(�<�9�D\��|��I[����/��I�G�{�z���n���[d� �Yu�.`˶���8J#
�.r'����ǻ24���`d����[�t`B�d�:���%U������7y��4�����	�[�ځ�Fg�Di �yQOn�k�pdpH8���p�;W�\�v���6���(�l���� -`I�
t��ɱzl=s�ZЖ�m�@gg%�Ӑ�<���|v (fs w2��.�5ǻ�ܴ�s-��!��B�O�W�X��f-��2[��/,�5��g�L�3G����� ��K#A��'z�S�M��Bki�����x�0��Y ��A�ltG0�7rGpС`i����eRV����GAn���Q��Q�'���!c���πza=�8&z��cM�LY�L�k���@��a����ck��؇�[�2��C�`07&{��2��G��� k�M���E��d-"q�R��s"��v�T_ƞ�g	���� �:�CM�{���:.w���.̇�N�V�����@$t�/��7V�W&NX���Gw�IvYka�\$�9���	���?ǘv�H�+��ނ����ˤC�P�(�|��(G6q�alp@���fΕ� yo��@38�P3��Z��ǂz�ɯo�\#�'���d%�1@��T�()�Ss ԸW�B��G��4�ϵ�#���,<U%T+�|d���,,�1��~�s.��i!O��tGe5Ola�Un���.c��]��)��ȯE�mt0e��8�K:ݩ�� ӣ?��x	�0��2('5�+xJ+�#�N�3����3�L_(cd���-�U�n��4��HxN:I���B����*{�3�N_����}��m6�T������c(zdJ��s���
�
>T�;�ep�L0V����\`1���@�<.ә���X&y{ ��"I���`�6�xĿ�P�h[V84]�eU �5In�s~�%�l���N��lvΤ`;iQ+U��O`��d=�t�=����9ֱՃ~H�"�T9[`��
{��욪�Æ��b�$:��GR��C|�1�LCg/:�Ǘ�2�#L"���ܶ �-���9�X���^�)�1�[^��"�-�	~�}�8#�Iӿ�� ?X�>9L�.s�b��pOQ������3���I�a�2�L��Uڅ���2�u6�9��H�����F��f�9l��B�X�vИo��]��&1<1t,���Lz�5��:�W�(�{k�c�"��P
�<�Sˣ"<�f�};��h|��k&��R6{kn�ʹӑ��C)�x��fR�f��F�m)���?�s��ф�wQ̽<��׏�d"G%��3=P���a;���1�;D�R�;k�����<o�wE���&HL��vQ�[+pךƺo���؅��*qn\���� H��}���xn����I��Y���:���7
���	\p�3���]��K޿���2����*���<O��Ie�,�����p@cmߠ{���!��1��}A10���P���>�!���A8��#����2^s�m!�I[|��깄O~ܖ��L�O�������HW$R���:�����:͝ ��Ĝk_u9��c��`?�ެ�L��'`{��x���O�����9��e�Bs��w�(�쾟�ݘ/��x����{��S�3;>z4ϱ^��2�_�(�+���a���)�ܖÓ����v������|^�r�\_�i})ZZh����z���b����S�<c��k�l�}\Wo����Q��G��-�[O<P|U�l����i|��}w{Ǯ����_%�L&ߠ0�F�_Y�.���&��溹n���/����~=�ˮ?9�~�_���7�xm{����/����T�-%*ú���.?��s�� ��|)�
4ψlT�p6WTՅr� ���Vo��~�'����?Z�����C�moI����)OA�5�N>2�zK�qV��;P_�ۏ�?���[�o����k�m{@sf�FG��1դEQ �cF�a���~������=<>�ˡ��|���;0� x�!��/i؅�V'W�K�|��0�#*�L�H���0::h�¡���d"y���
���3X��D��b@��[�� ���̯�r���3`?�!@⊤����g�:�<h�/�lf�r��q���X�֩��`�?�S�Qa�}(	 �"c@f.� ��&|�<��ų��Jӯ��ӖH5E�?�@�G&����7�VT�Z��N[�Y��Y�V���ʡ��{థc��շǨĥ� ���Sp��?A���d�����N+�$�$8��N������ؽ�02Jd��q��;e��E�75��-Hc�c�@O�ro5�i��xϼ_��0���Bg=���ǡ&O�����\AR�-�1�N����&oX�pLd�\�-ݤs`y� �"}����Qᾠ�yc��3B\g���P��@iN+�u��]�l��np|�X����P���~����LtР���N9��G��U�p2�'*��xF�D��f7	<�9�{%�<�+�Ζ��+�	�>Y4&+��oI�"��e�`��`�Pˎ���f\悮N��c�5�s��Y@G��|W�Z�	�H8����P\��$�%��Ϻ'��,:AeE(��N���ea����j-u<d  �Ha@x�gLB���h�3j��*������I�V�[��m��A�������$+{L�ϖ,6��_z��?d���+�8����������S��v܎슔�WyG��!�Uy�n[�(�0Mp(���Q�it��d�9b,�g|LQ�j�=L�i�ƪ�������q8���^���ߛ�9Ƃn1�C�&e�H�jH�E�Fޛ8��#�j���Ԥ��Hΐ_҉�IN'ϲ���/����ɡ���+x��l�^�Ah $t��zw�� ��d��_��2!���*��&�hSp���v�N%S�3�/��݈ޘ�܀����~��Yl��tpG�!���+��[1f$1�Pc%��Ƙb��[<g���9zDN6_u��	x���)hr��v�H��	&-~M[�mBގ��9!0S#�*�1�[�\&�$>i3O���1��&:��-�&�'�M|2�fT��xNyj@�P���H"�A�L��l��x��+�>h�u��Y��$�<��#�H�±*����3?����	�M ��bT���I���Q�7����!��E�1�լ�Ĳ�[�Ĩ��`�˹�X��	N�d��j��l�\�W���r	[�1�V3H�D�TN�5X.�U��o��46%�ve�,�d|�Q)��;���g�.���h��1�d�Bހ2��kAZ$ǚA�����7�jI�Lv��$.0GAaOv
 ��h���-��Ա�3y�֔�E��V�[�+}y�y��$�Ƙ���Bw�G��%MC��1l�'5����y��gP���g���I�Ŧn4�c)�[�W�L4Ml�x�G�a��~$;@�!yAv��X.i��3i�뱿��f��	{*;����#N�CP,�羣+����5Ħ�?\ɩ�Xr=p���l�P�?���X-79u�R%�����#�l��%`�= >�<�R����l4���z{�LtL�d�#����tB���E@|����-�8�&s0�ƀ
�5�L���x�\�=Rw����kw��?�}/Zyt��͇��y5J<A ;\ ᡦ���(d�q�^��^��������ŝ�o��:x��	��u再5�|�Ȗ걪g�{���O�5��_��ݷ�vu�;�o×�X��dЂ��y`3$dW����?����[�s:���2�b���n��7��;�����g'ps�\7���=��=`R孷޺�����W��?��O�{gO>��e�������8�PCX�6���g�{��cV/����y-Ct�E�I��� ��s?�i(ۋv��3���o�;�=�z�]��jeH��B��v�pe�1)?�m��0,�G��Ů����o���e9�Y�1�i��Y�j}��H��f/>��}�w��TG�A��]	���O�)���%��M���������fZV��Ѳx�B��QV��d1 &��Юl�L�]yvR8ƥ�������L��ah��y �U�����6�+�U�o:��'�pPdu{x��ۊ�r	��cX�Uj��&�qȚ3������������LUJ�Q�3���l��p�w��~lZƯ Ҵ��l��0pآ6�8A�p�&�3���k�I�Ǜ�6&?��0@͗-�b�W�51.�s,*�pxp>XKC����)[�E���N)߅D�Xc����P�p�b�8�N�m��7�,�ƔF��rIY?m��9�g�3b:�V{�"�٤��R^`��!�v���#�M'B�g�?��� ��p��|O�Aj3���KE;�P.q<�s�%���G���x�<��P?c��A���s^�,�H31�ÈE�� 8��M���ܢ��� r�P�� 7��*�J�V8xLG;I*	>nW�k-�ؙ=��R�=O���)%I\��55���f��P�E%wq�4�J}��ej���4�`���,� 3�Q&��嵐,2p�U�K��~�J�BO�� H)�UД����zt�s�S��xQ����Y�!m�Mǋ�����rwzE� LCh�z�-���i#��hedX�Qp6�宅�S���L�p��G�h�	ߞ��`���T~kT�e�gb*J�x'5�Y�s�$xb$�g��=������i/WG�����A18F�;xW:A�� �$���r�ј�<��1<׷�#�Φ11�!�y� XNu�kd���M��&-s6�E�2���I��9yLǨ	v��^�|�O{�Rv$M��ئ�����k���B_d"{���.f���q������r]O��ְ~3�ҵH�%۰��QhU�c��L�
Y���m�s��Y��<�����N��Oyr�b�b��=��E:���_���6:�>�����q0
��
t.呥�*�"�\F+y،��@�c��vC��`"k��S!��;ɻ��q�-����7�i���i��j�U۴1!+ƾ�������$	��,2��b�-<�%����7��7��.��U��B�x�Kb���}���b�	J�=Ӹ��T�&?1OK�c��z�Ӳd�w�k�Ĵn/�!�c��gL��u��ؖ��5p�^cg��G�jq �':�U�ƍ�����:�$��D�"�9�v��V-�{%��QV�����L�^)��������(��Jž6�(��d�'���n��>򱵹��'��{/����M�r�ԡ3��茦��8{'M����`��;�/f�XDއ�-y\撶�lsk%������9�S�S�����+i�9�Bצ����@�u��p�Aa7�	2��Oh�m�s+����Hɠ9�� �!���߸�����l.C�ȱ(���{'�r^��v^lA�,�뙴lĚ)����Bn�w��5,"���Z�MHPI��t�1.�T��>U�x)|mr����*��|n��ڙ��U��|'�C^������OKLۀ%�c��:^�v8K�܏�Y"�2A�I�BC�w8��>�_�����c���l{�h@��k*���i����A��'�����S���܏���n��vat���@f�ߺD�',��6��{z����|�o�/��c۱���K3�7Ȯⶑ��݇�����w���v\��Q�N���:U6"���]Y=������������۷߶���ٽ�vs�\7���=��5���Y^�����_���۟�ny���z�})[��+̄:�W�?�w�~�2��G>f��Ȧ�!��J}D����!ob���,q�Q"������?�����je=�� o��n�F10vZ-j���	����O��ϊ_�Њg�.�R=;�n?򅟲o~��W�ѣ���ڱt�<��-*���/��ޚ۳�����/�W��{׎����hq�BSO�9��?�|�%۰���<ۖ��٩�ʓ��܂Ul�	��֪�}� 4yĸg���L'v��=��f�N�������9 c�@��7x,�F�T3�-��A�&pL�n؍O���@��'�d� بO��+���u�ٟ6����p�uǚs�u�Nlv
�%P�W����[{��be�����Dd��e�2��s�F��mB+��d�X���i0����8/��oҀÝq;�`a���㊪4|npn��"�8?�؇th��8s�+	}X�݁*Ņ��J��ԡc2>썱_����PԐOY'46	�L�!Y��-���;͆S�yq]�ڴ�t��>g�R�j7���2�{t�Zt�K�W�{C����y��k� j
��c��9���{I�쐀 ��{�%��}oj2P��"^�	gz�5��y�B��b�͎%,���ym��S��kZ'�
�\���pZ��<�b�7IX�&��E�v����y���{�Y�&��l�1�N�"t�ѹDo:�����K8���S�@���`��s�bM-�qqg�W8/���Oq`o\�<�����+�mgelxF�ߐ�!�T��\Ҕ�R�!c�#Fy&��MEy,P����V�~Ka[Tvǚ�A�	���ty̽��!+3O��Ԝ���m&{����YV$�����K�=���I�������^f^�y֩s���� m���$e;0Y��si�*�(�MW���^�3�i�����Į�ݝM�F<���zb~ ��&�*���J�[��ic�V�ّA�����œ�TgNȉ�v��·��S.��(�oN�����`���L>�gk�Jc��ں��!��!wQ���������t��%�����wG�M�v��!�,d�E;i��ލ*�L�D��IW�KA����[�>���c��6�XLxM0�x����!������lvM�~�p��#�U�h3�+�/�LYC�r�=�&s��6nqL8Gx�X/�ň���o��繖r�
��CnO�����WD�#i��(�~����S���t^Z"�[�m+���#�y�˚�IWhi=񄦩�|N�y�H�dPR��nԶȘ��7�9�E�K�U���^g�AE�!�;hJ5FZ$ʟM����Ǥ���5d��Q�B�_�	Ew/��f����rA�R�L�~��x�T����&��������H v�R��$�~�eN���I >�µ8�,�*�O0���f6CK�~�'M c�-�^��!5O�.�l-�����#H�d�,��g�s�B��(KPВ�!��G=db��L�����Yг����L�w�8H�jW�}�gU�}�6x�������G^��K1��u���x[$���c�ggp�o��I�5���;�L6��ˤ�	�A\�Ϻ�-d��?�c��W�_׿ٵ!����X���"�s^���/�튧�vzT)�>��Erk��,���}�6�;E��m,x�\�H�_.�W��Mh�Ϥ͚��ɋFzO�0���喼7ˎL�O3b�<�p�l$�����$�p��ra"u��ˤ�sh�a�7<		OH��+@�Or�h�C�&��Do� ey�[�Տ`�u��+O}��^�_}Ξ�{��wqn�P��ж�ۇ?�I���h��;�������q���^�O����-{������������wZ��p�]��r}{ܫ�x�ֲ��N��{�~�oكf�G�Ny���[����G����/����?����o߹�\������к�����us�\����� ]⭗Ǉ�������X�yf���m+u����ū$ť2�V��yww��L��ߕж�p��� �=������n�/v��o�wW��O�p}�ُ�>�e=4��|,
8����f���<P��- B�,CI�=��V�җ�z����ww�~{W��6j���%��p��i�_���n�~��g��7�e�~W�|G�S�ˢٗ�SC��?Aidg���(���y���[	bL�*Kp��i��
³B�����@Nga_N[P�P�٢�m��I#�Y|�=������1V�b8�s�V�n��l7��/-�RV�@�%T87[QJ�Q턷	0�g4�[�W@L@8������hK��y/{ 6Z�i���p���&���AJ𗕨����O�I�`haH����7��-;��j�}ιûo~���#�IQIF��B�/�������� �� ��pC�H����lv7���~ӽ���VV���絨�I3	p7���{���P��_U���e�t�4z����Qf�3�f	Ѿ#h˳3�;���r�=)_g�dt��s'J�Y[����mc������ɕ�4�@�ܺ�%��=���s*)��|c��Naz9\2����vV)��'������{ʎ��%G���;]�LEk3���N���V�5UZ����E�ǜ��֠I�7��F�MZ~�wi��� 
Br��Rák�jp�'K�a/�?��~��w5*9Ív��� ���:�c1�(�N�,��&�'�4��T.��{��Ok:[�tv �=fG��l��|<�.˳icF�
w8���HQrn-'�}�x��C��yyY2~	�U}Ñ$A��9iv�deQ��{h�lM�Ѣ}JC�;)�A2�bq�n֒���+��{�.#9oC�v{�VR�R�2�ӌ;� �L��Z�������v����%}�y$dΡo ȨCW��}��1Y�����]� ��>�D_� �S�En�dr�R¡�4�C����!�@{��g1ι]I $F�3�qZsl)�8�ԃ�yA��H��e>&��[�H��,�	V�5��M���}���wW���~�X=8i���)�ɀ%�p��'�fTGH���+�dME��!��.��5C�����f�d-أ�{��a�g lT�h��"��*�aos�T��q�Ȑ�'����K��qz��,�1��h&��r�$�m�Z�(���/M�(F�A�x��?KJ�3�|
d�5� G��݃�bВ~���V�`z���A�s�-�qt��m�����}���땯���	DكNeό��Wy�?X*Ӝ
���(���n�yP���u�����ݫ�e	���t���n����-¹��"�饏}���%��8O:���G9�5U!w��SSeٱ�Q}.�G�������V�����tF_
��{���:��q
ٴh�B	�I�C��מ� CY	��*��*Y�@֭�8%�f�7*�5�Dq?�]Ά��ˡ�=��I��Ob���5ˌE`���F�L*ɬV��C���n\�$��uH��+�s����Q������߳���Y�N7�ָ��F����YD?	m%��ʆ������?�]*o���K>r�8K�ħMn�*�q��q�A|*�������̼;��h�R' �c���~�[��.c�� �Ї8�<<h|Q�`���ܼ��� �������D�\�����ٱ{�Mz�L�؇\��|4S�������P��~��
��+If?S��\���R�ɢ�S�XJs�����Np۟Ҟ-e/_*K��T�f����)p�T~�-J�X
t2����/xLq�ɾ\���|�|�ř��@�I�K"p���wu>K�)@�eA�W��2}D�أh��X}}g)��:�)�U��d�{�y�^���߃-%2��?���ę���$����.[�<��䄻��|sEO�3Y}J�\��[�1�{��o�m+�� ފ~5��8g� �c�T ��9��*[�����[R��hE%-	U��W|�'�~�Y����P�����B��.h���+��I�7�>>�A���������R�^|'�=�C3�0��-�{�t��.߫�cE�����$聼g\��oư���?��ѽ{^ٜ<w2>�	]\��uq���� xܷG�����n�y޶��0 ����;a�,$�/+fT$���x���tܴ�}ij`�j��d���H� �:&�?W���߼�J��k���Q_M�nE�A�Ϯ� �Ƃ|�ZY�g���ϱ�߅辶~w儕I6��O�����e����?sf�жxIcqrLj�%�a/e�ƿ����9�x�&�~�=z41���<�Z�#k^*�� �� ������Y:-���/'ҋ�%+��h�n·�C{�g����qS4,���S^����"�%ސ�gtJ��9���Zx���Ȫ��m|��E�XBp�< ����L	圝�����Y�7��c=\�N�Tc!��%�i����0H*J�ζ�(Y��3�S8�J��,1��r��^!h�@#Э�`�C��M�L��yO�贁�n.�+i�$���<u"Τ�J���#8R�_�����{
��L9��%iZ�Vq���A2O�PZ���ύ�mV_��+f��NG��c����]�G�D��QD	���g$2��Z&��x�B=e[7u�j�R����/��y�?T8A�U��cyrnh3��3|%Z��(�]S�?U�i?����x.���+}���I�����(C�r�;��D7^"ԞU}m�C�¡�}����Cw&U�ۏ=�������2�H@0�!3A�5-t�ha?�X��32��ȹGc�����%A.�wa9�-;Yzr� �����]	G\��7�h��)����3^�D㙎򸶿p�����')�G|�H�
�s�J�C^�g"�Z|Ne_�����S>���&2�<H��:� �I��1��i����7ЇJJ���Iq{����|�1j�i����jM9��3b0� �\���V�����EV�SР,�3�i�O� )�\J���LSOΕ�<f+5I�l�k�G�����UW����笞�L�x��=_j��4���yj-��r5d�*��A��>�}Be��ɒ��0��u�tӾe�r����g�=?�$���|���Ȍ�&P��y�~M"0d4����~�]$45's�W�)O�M�������q|��=z��~�{6��F��'����feNN|� w����YS�\��s� ӱ�J%�A;y�p�\J ��sθ��Ɂ2�,o�B(�L�|���
�/V�N��#�oDj�E��Ө�Pm�� 5��� �x"��|ϳ<��!�R�)z��c�=�^�r���Q6%�]�HY��;�����
k���~-y���9���5�����-׺���]�t��&%9�3D�����
��~�[��8~�G��!W���8�#�B�3�r��^X�\�
NS*a<^�
Y��N`!�#pf��D��l�]0ۧȊ�,��dأ�� �w�E��E]|>�$�p^��X��C������8���|����i���#��@�!�w�W>�����x�2l�O)��=����)�|^�E�S=X֡�=���"�����K�� �:�W��]n��R��l��{�^ø�k��������)�\�QZ�״�^ߣ�� �2xQ�s�:%��C6���	��@��4�N�'�-O��
Y�(=��z�`��˶r���=�$��Y�s虉Ǉ�E{�^�e_���g7 1��3�b�|�nd[����{ .�.^��+ZڀG��ۺ5����	}[�ǆ}��q�s��kE�JQM�P�� @�_�
T�#�Ah�Y.��פ�B�c�����ڪ����ڈ>֠oN�⾽�=��;�e�sn���W����L/>u��������(�c�v�ط�=�$�9������6��$��4h{������^�&I�����C��Kw��"�~��Λ?�9��������wןLa����W�h;u:��=8�w��i�B���|�	kf��%:� 8*S[�}{�ɃO�ܝ�^�_C{��⺸��}}�L��w�G�>�1�Nez<$Ŏ�l����C�"k%��wf��F_��4��v���-���\wj/����YPr��/NG����}}x��p�p+�^*JQ�B�B��vM/*�~A��߉�������[�c��:�g��B�z�yz���4�>%f��c���n�NrV2Hɧ6��Z��'��I���s���ҡ��
`��)=~>y���L��y�!��(�B���� �!���D���
xU�m�6.W��=�ж��52r<�>)5�a�	�-�q��hi��z��h������G���:T�o<PP=���׷8�\Ϸ;%��`�����yh #:Q���i��P�f4'+��f�e�Z8�"�����dt�}7�@ ���8��������N%�+��M��TDeId:[G8��f����y��)�^Jrb$�Ncѯ,A>�dl,�=@;'�(2�xo�i�%YY[w�0��	s��!�h��y�gb^a�n��_ȕY#�[P���R� s~,�!3���	�c�.'g��T�Mv����SU�@~^Sb�&/{�r0xj�,#�-�k2j���D$hfYY�p(tG��,�	��y����L�S<k��� T0q��M�t��J��3���,�� i�l_�M?+p�4��$:J����<��;J��q��k�g�����y���`.v>��8�/�����<��O�X�ε�od:�!�K��9�vs�c��A�jg���g�<�pB$��`	y�Ik�:��kgz��8�>�l�������{��pG^B���u�p�$�*�|��� ���=\��G�֦��TT�X�Q��\�xeI��Ą�\ ���p���8�ñ���D�r����w�w=�����D/�j�{�酖^	={
��l�����g��Zx��ErK��s}b��䩌SKbW"���K��T`K�99�g�k�Y[u�-��Pq`&-��Գp.�p,g��K�	�C_�C7(Ǌɹ��n�Av G���9�>�c9f�7�|�h�{�#t�,�]Pi� ��9?Yd�&ۄ<�Ξ_7�c�����}����#��5��M���+;�.�yԨ�B��ݞ��R�a �z�/�	A��񠀱f�!6=��F%|L�Ծ�:��؄n���A���2ƶ\���Φ��U����v�>6���'t�7����ݖ7�V&1�b��J�݂�6��Q�/�_3Y'�e}���ر�'������S�l�����ޭ���§���RR0�hc��W���2t�{A����u����x�ӓ�!�4>'� 7�*O0KB��]��R!?+^�M���g���&yzA��sƟ�h\�+���
�s����;-u:X���h]�;{����3�$ ����[3��/!�h�d5 .6��=�wܾ�J���?��.yE�W8�8}U���a'];WWɥӝ�u��`��*���ɹ"������ J�@=X�ux��Y��e��:Q>_��Tӹd}G��E .P0�����R�_2 ����9�:qz&?c*:s�����}!��� �Y��ϳ���{<�=�
`7d l�ۭ͂	�̱6T��9/�����'w�H�@rT�j�.1����X:��o/+!v
��r�?e )z��ҽ�l�=���S�
�:=�@�H+d�~�I�m�ւҺ�(���T�Xc�����`��~)�g�
��'}�JF8�� �z��K��G��R�O(ݣ�9kmqOOP����-��h&�v�:�I�*WY��tN$������"|��1�N1������3ݹ|]�A�dLDΗ����v�C�
��鈾�ߥ[O?g	�GO��.�+:�X�U�m�}�w����;?6 ������Z��T����s'��/2ԐI�;k?��SJn�79ǡ��2�fM�Y�{t����]\��uq�M�� �������.����/M�D�Sv���7�gYݬ2C���	�V`�C�6)��hM���`���1�!���ڿ����7�4-�?5N�7�_'��O�� 0wx%t���i��>�di�_LLe�%cbbeE����g����aK��y)�-֒ᛂ��(��1С���<sr��{�!��H��Q+ZaA��4��J�(�2���<���k���.���AC5��K#����-�b�xYsh�0
eĴ�p�('�9-N�#�wE�u���B�y�r��d^�q�;���̩L�����lX��=ӅE�;�\��E�1��*����+j�Ie�����	��Q��%/.�w��������j
A9�D�^���Xp����{@��%r)�d�s�p��T!��NW6�ܪ���Y����'��vKV�%����L-|7�-��j
t�_=h	х���z��7m���{�~&���Ϡ�_��gq>)2�	��{�o�����6Ÿ��uH!�ui1��J�"k���\�o2D9���WcS8�{kƥ;)�'�-&'�:��/]�A�	�B����R�>���[���<�rf���c�KZ�e	E�����<����,�DZ����G���F#s�/�9�$�X�P���|��BmE���`� �<T�2u�K����Tǆ�DwF�g���:9��~�gB������t����kY�A��`������y�Nj?�%�P�`�"��P#u*�H�,O��v�K-{�jٟ ��=8d��"�-��?��zPϡ?i-��@C<O�Q���%��?��@2�(��O�d2=����۽�y��:��;� ��@�AQ��lm	(��՝��.�Bd�{���Z�#>K%*i* R�<kIn̏�5;�@C�|5����C�%(t�DKp8�� p1��h�{�5��������?VB�W/���*�&�횙�e�9T;�\��I*ڛ[A-Z��$�+W��C���@U
��>�] �P�=u�r�׭�3��@�O�M �"��0����^\Ǳ����x�q�Q�,�X}3d��'{�?�Ϗ�s��, ��V�4�`P�-Ur��4���D�=3��)e���1� �!�YL�E;��C����Qj�q�:�JY�`'��o �t���I��c��he�VMN?�c�6 ����z�29�5pn�Ne�
����E�&�Zq�95�O��k��_ c����f���OjC"��鐱�
��tT����\E ��i5��v��J���'�7�#�R��<�����}�w�=�^�Q"_��<������Isމ3��As|D���X��x�?5����d���'���I(]lzI��ޡO�>bm�Z�M��F���{�-�:�g5��5�;�U�C� &��4�}}<�t�@>��Su�: ������Ƚ��˳Z)�v��F��]�<�#��Yr�rzd�ڬv��q���>�-ݯ�tj����XP���ber>�Z@������0,x�7�.��u���w]'B��� ����
���^J:g �g`+%���8�؃Л�R�d ��u�z̾��c��}QJ�!�P}a��S�N�"��@Nr{����!A%��ʜ9�K�ʙ�B��s���@f=#h��ya�5�3WR�3��g�S蝝�u8%d�gH����hiD�=����J�|��>W> ������O�� ���5���eK~�$��ˣ��Z��8`�k}��'�����¯h�tk�5/�7�BTW��X���T�f�	�Ә)��V0�������r�=�YZ��7hקՓ�?vG�}|2�@�ui�uO�>uxD�����G�A�D�pZ�9����6��ʗ�!�/L��y�3����{X/���v��7��/�~�?��Nɗ��*:���J�yl�{�����%�Z���v8�f3h���-��v�iks^h���^�g�<�ի�5��<���uq]\{�� ���z��?��?x�����/�nݓL�B�
`�)"d�l��*�������`�?���*L������mɁA���P�%x>З_�v�Ӻ%�U��?cQ��������k~��W����v�|�|�*=��+��7�\�P��}!��wv�x�]���9��%(�a��9�N�@���OlG��Z
����B��A���%��dX���y��L����%)����n=�R܀�eJ�|�s�,[<0B��m�'�z�fe+��\7[��%��X����CA'S�T�2��y`}��0���=�$;(��JgHA2��/Z$$��ܣ�y�gS�x��4&4���J�Qd|gG\����_RRa@E��"�x%�OK�D�og��Yg�9&��l�PR�_���5C�����k"sޏ�.�zV�r�����3�b��`Џ��ģ�5�DO��F��;1N���ǲ@�~y���o,�s�AT/�'�A�/��,0�����sj���z�3mh������Y���$��#���l$����U�p�UE�X���^^>��Q��v�cG��)�iz	�������9�����q���&���gD�Ԁ���3�襎�q7���Tr�kΈ�31�f��M2�cl��ا4�\�k�˗�܎!?�	Q~��q��M�'=��'>}��6�m�=;I�ZU�.�X0.��
pZ�E8.��7�W�� E�_	�L�}WC���D�{X�DY
��le�W�C��]��XW��ƅ����m�������2�(�hA`8�=vk<���,�2FY��;Yo��Q*�k��51�.cO� t��_tʞI�x��+d�V��&ٳwf<Pir�%�����3 mr��yڣ���L��jT�{���ξ>+zfc}���,5���vE	[��)/1�X��s.��]f:�k��y��$�1�0W['�s���x���q�F�U�^��g�N>FT�:ui���`p'Y��z��)�1+]�3'&ř�.
�䎾��t����������ʟ���b8m�}qV���S+�� �Ե�q�����b�/�;�{ɓ.i68����n��7&9����U�i-��Vr!�gO��|k#`��(�5�>������E��2����$��b�</�k6�B������1�g�1c<��=*ci�@�Dϛ���m.������5�]d��ր����g��R=��r~)8��D_zְ����(&߱*f�^�\yS�1��W�3݄h�:��;�f�����Ї�=�hr�|�N��|u�k C�hkY�zr�ӂg��j�@��V( r
��dc�%C}�Ov��h~������?���h��)p#@X�������G��:�-�>-��	z���%0E��5�4��ÅoaO&*8��,h=2xAb:E	P���B�����X�.��y ��NQ�p ,ӓT����Z�������/���;�9 ���������6أz���}I�TC���aA;���85{kT���;�O�^��3|�}z�ݮY��zw��t꠯=\���m��Oax����^�F��A9���2��>s|7���SOc(T���FQ��8�)d�gm�
*�u��t{���|9�¬��u�Vag+�B���)��;��>��i����3�i����E���F3��$����3B����ɪ��3��p̠�f���\V����`��g���Lg��]�}�����D�a&�e�֬��)�����_��/��K�6.�����~�E��@�MO�'��T_�;��Q�:�	:o��c(&S��$SH]C{�νk����b��8N��X����V�ڊ��q��M褴����@�Z��7���trr]Zx������RYҹ|�xM�'����mz��������[?'���#��6���+]s�՚�d���GW�㇏d�Zz��mj+iE��ˇ'�o}�wO���_?�6�{c<�y��|�G�⺸.��K�� @�=������������w�����U�7��F
3����fQ������;>�swo�C9Z���J]�g#N�>E�Ю̴�+:uZ_�/���~��Z�oC�[���a���`���JJ3�&i<�������*Ҟu��_�z��׾�mz��?�6��3�p�+Y�!Q����|p@'����O�9I����kǚ��ۄ<��j�rg���L�������}8�`P��P~�gj����D�������a,�� d{DY}dפ`3l��(�t�t�8���&X��U���r�h{@�g�_�a��b�FN�SL�*���y�ٹVJWq#�L1P�c9P�2��Q��3߬R�)�HB.��g�����P�҆�i����w��s�%F����!-��G��.L!dE���ƘOw��G7h�D��b&kʶ�n�i�D�?V���|O�$�K�zv"L�d�:���ߛHQ���mg������{{�D8$	��B0N�߰�q1�18�ȵu��ud�C�Z7|a��'�@	�g�R3�}8y0�0H�~V��e|a�e��g�x�g�AP	�<�&�l��72�e�=�`��3g�5�gZ�5S�D&����d��q+�v�o><��m�����}���%��s�s��n�~ �x&��t`��Ug<�c��Ó�a�p���?k��L�n�R���^�|v*��5&5�瞜=��\�̳�J�=��n��R�9��:�9�S��}]h2�6����$ܲ�z��#wGք�>�Sޤ��d�l�#��X��/�K��,yY� =�l��OBT���5��(��K��Z���k��Y~-2Ԡ�����u���5��4ú%����`�]��u�l����������zO�ѥ�H�cT?n���A����������ל�x�������ѓێ@���ڃ����K�����Uc>�4V;��3H�#�p��U����V9#���M�<s�rq�,:\��<d:���Ψ�q����=�a�z,{ٚ����E9V5Ǿȓn
�mKse�ڳ�tx5*�pv���E�/�c2�3Ӛ�8�2����>�l�e�!��*(�_:@DM��x,��:��H1y8��54�͙h�A�7�D��´��i�F���
���!��3e���)7՚o�3�w�y�]y�<�n�b����8�T ������K�
Zo��h�� sh5����^��kV|�.�z,Z�:�I�ϣj�N�n��'݌ڦߗWy̤:��ɰ��U�\��C��g���q9�S�A`ʺ�*Yv(?sU"P)>w,˪�8������.b��@�݁��A|^�"� ��d��T� ኔY��q��/Ȟ��q��3���>��9���yN��)�0%�RJZ�G�a7����s��RWy�g�x��}:{���s�����ɢ��m\�՗�K�Lo��������u�<������E����́�A
�
�נg ��W.*Vr�,t� �!�U�>�ω��65�
s�P����ƏMU��>ƿ���
����/���	�0�tB�o�S��i$x���|>�d-�V�Q;{�Z���.�#����Ѝ�U5�3M~�`�ۥ�Г����C��I��e3�27��ݲD��9�c6mt�tє������~� TC�@�)ZYC^��R��VPr�}@�	gI�Q��:D��A���.�L�?���d���� ��o7���>8���Dd�˰׳4پv�ױ�7�Ψ
�<�V�5�%	�J�����V8�g~�`�� y2����2*�ǻ�X���fϋ=n�^裀ףϵ�r+H߄\=L���| ���t<��,<?Υ�P���Ɋ��N����.Ia��h��frc̥��p�7��U+�V2�9 �ڦA���Чs��)h-Q<��a�v�G��_��v6���6��#o�0�v2}G��D�s ���E3�%����Pu��ޑ�E�b�*N� =�]�쓁T�Y�I��*Ǆ\	�l2����������0���zN�Ql���E��s³�Ǒ�%�=�&�����G-\"�&�GhIO�{m R��i����ч�Oy��a�SF�) ���ʲkd���:?������O^��B[�f[	�`e�zDx ��`?n�Da�Yb&'����GU�,���y"����[ܺz�*AL��o!ǚz,�W�c�s�y�W�l��L^�~͗��b�tV��R��+/�~��?��|_��"�d�s�֪�	���t4yo=��|(U�7C�~0��u-���&D�D6��X�q0������?���;=\o�V�����>���.���⺸~���� ,lڇ�����7?~�㷾��o�GeˢF]2f��K�`ce���%Qؠn��.���N��G��0Pi�F��|�c�,��g<*�s�?K;I��o�>/?��9�����F����
;vn?�4�}�9���{�������^��P��}8���Ua:\��R5�cuU�<��-��j�dv{>e5��^x� "-	�s�N���AY8G���w�)�[6|0e3��%}����K�xiil5k�;��l���+�p�g�p��D3�t��I��3u�pJ%��hM�@� �[	Q9��P�;-�3-��#��x�ry- Ms�c(Т�[�0�?dƅB�ksN��{�^|Z��4&�J=��֖ʥ4����Oq'K��,�}�M�,�������p�{8 ��.}_�b{&�P����T3��1�4�V��x�;B�<���:d��}�,P���L���N39s ����gY�'�(�*��^���ʻr5��2W-���/�ǰ�zx�O��K+zٷw��1�2c+�=�k� ��]�>3���m	��퓀�jM֌�H�gyp�KMbz'�8F�YTX��y��C����! ��!����S̀jA�L�xm��1:-�3���8c��������c/�Lv�C&ľG�W�s�|�z����z��5�>��߸CyM�f�S3Rf+e�z���` ?˖p�j堉��F�S����4��aCu'�~р��}���]��� f����O�φ��9�c|��~e�E�׬�.�<
��L�%�qѓ�r(�ٯ�� z�Q��޹����m�J�%U����]³)�ú��״~��,M|��� G�Gm���bN����DƠ���3�B���� L
x��Z���wȧZ�Wt5�uk��J�-��G�W=gg�	����)[�v����z��q�'��jH:�#Q��3�
�Ņ�+1�-�������>��R��b�<�}��� ���v���R$�\:rY����
��9Uf�+4=��Ǚ�4��b>��EϬ-䜎_ι�X��SZ��g�tԠ��KC�Ε6�3P��9��f�aC���u�u��	\����zقIK�I��d��#��v��	��1�(V';�Ł[K��)V�g��Ⱥ9}����y��h� g4�g!��\17�G�dw{Y����`��6P����s�R$�.Nz�j���Y�kP�Y�������	�!��jyK��x�Q��P5�)�*7�.vsTL0�}Q�9lY�l
��8��R��cH���_�ۢ�A�`��=б[�$������w���쀴@��Y0h7^�>�7uۣ�i�rƥ
b���I;�-�de�3�A ��	���gr�D��e�M+V��hp���ZSр���Y�U�^�Ȧ�z� , Ϗ�9���@=��@�f����5%���}F��Q@�cp�H�7ղ�]�"f�*����f�&�/���Z�"B��*=	�2�&���x�Ԍf����2}Q)v6[L���x��������6F����v�u���l4�x�*���57ݱ@w*N#hE2O�;�v�a��:
����"4 �Q�}�ؿ\|Dj�X E�QUǰ����P�V�w|�Y�pߎ�ظ��r�j1��"3���Z:иwׯ�71<���v��2fg%�e��,�ms2�{r��.����v
�R La����@3� `������#C�u�'�\��k-y@�6�ٲ��n��y�9]O���^+9$E\2w�vp:/6:k���*t����X��4!Vд��v�8;PZh�+H�|�]:����ؚ����.���9��Ô�w�����Flg:�u��u[�oP��&�P(_��{u��$������U]$«�ˠ�ْX�^��ZF(�v���!mV��_��l�W�Og��sS�=�xbYY� O@#���8��q�2����(��Q��Z���Mz7��J�� ��
@��ci�g����=)j�������3ڝppvO����iO�'�� O�����͐1���u=Ey���@�Y蠫�n��� |�����Zɹ{�/ҥK'��jk��a>��,�(�$��L�Cyxᅗ����3O�r[��t�KY��WS�ui}@
�P�����k��2�o9���=��݇C|P{}<V{�w��.�������� �Avf��ն��)o?:����&�w_԰VeQQQ��UV8��Ma�@�v�@��(�e:����f�A&bǸ(|�)~��q�'R�uZ۴���?��0f#�W��u�7���l.{�L�O���g��hఛC�`���|F�	���1�؀ҠJjB���U���8͓�^�Dɋ.�B�fdB��� S.b�P�!��p���.�5������	����j�n����9�\Aw6�E��b}����;�]���&��e�}���>�y��A`n����C��,s���9��3Ŋa@��^� �#����?�t���GO��E Ľk{���_����h�*����:&�S�ъ�O�� j�3Ӗk�M�^�Y�%Zm��p4�95�T�Җ���{���pp$�AW�Cii�����2�+�a�ͅ����"�ޞ�����o o7"�>��	I?c��3�%K�3�m�(^j * v�a?�p�W e#F���/)�snA/�����3�J�ry^`IFyG�y������i�zzV8�����@�q�y�Hec3�U0h>L�k )Al437k_c��N�!y%�I���T�l�C2@�G��9%��AN[w8��G������,)6N�Ղ���i��k�����<d*��lu�+�Z��y |� |�P�p*F��%XO���A�0�@w�n��tY����/���g���KrDi��������b�'	]��ëʸ2�N�G !t�BT��W
:,�9��7�@�iBKJ�D��<�";3-=?�G������[D �U�Ս~�U
� 9 ��Q��%	�������y��*��]��d0�<�)/��=�ayN;�ҊP oP&�ɢU8�&�`e��X��s�E��wo�����`��וǵ��Ӂg���>qhu��14 ������1${�#�M�2r������.^��Ȑ�`�N�]�<��!�+��9>Y`�P���v*.��}׵�gj��Y=��V ��4�g�+������9bQ�h��9�s՚e-2=��i=�L2�Y�#.E9��_T���͙޻���(��q��LGy�@{&�3����<������srb���4��H�-���Ł�i�-�(!�z�}gN�%8�afz�V�_�Bؐ��f*6_�#�$�W�"���n��^C51�ϝɰ���nYt���J�}�{;i}��I��U��`�*�f����G����%�@�c.�N	ڎ��Ӫ���J"#���~d N�{������!@~Mr�x���\���i@RΡeE�^B�א�����ez�f��C��������g��B���SD�h]�`�
�Q�;$`k�υ�E�4�̗��g���d1�"�j�=�P�/ L���X?p� X����.y�l{E�Q,;�sh
N�s�%*���[��4s��Jv~��yT�`~���l��ȸ�y �� �� �Wlg����3��@�9��Ux�u��n�I���=�8�JTA�g����~@j�G��Dŀrh)���XU?�T
�W�I� �MV#��|[Ƀ�4��
��Ԛ�8�-�����ӹ
�$`d����J1��*֙�  AVm���p��^K	�:�=��,�[��M2s-{���L�fY�'l"�:�K,SV�>����d^�U��M6*Sg��]"N���bo���.�L�zq�G�.�/@ᢣT���DO�V*ʬ�NM���Z͡�?�M�I�8L΀�l�,O�w��v�6j>n?od�ժ.��z��5�lj���)�&�.	\��)��di�Gժ��T�cN�Ր2�g�4��!���?��M�y�חhC�֧��%����z��by47�4grB�	/��NQ�j��:6�2_9�w�1�~���w�h�5������Y�*�� BЎ�"�=��ٍ���|�����h������fG��i|���a�����f�[!��Ϫ`:Tr�yϦ��f�Ad]9�=���O����k5�s�=�$�W��64�o�y�d��ds� ?Xb_��ã��h��ш��k�P@|�>�_��t�V���~���ك�>7�۞���
6����j��-j��t0��Q����oȐ&�i�h�9�9�p��yg���:]\��uq����Q�����=x�������?��ۗή�eÜ�� ]�Q����H��0`]�e��Ijlk�F#�U�u���ެ{و��&��k������?��++�O=}�Άp�ٌ��@��VP��,�@�T'��~rB�{��!5(��K@F�Pf�	,G
f�K�Qg���e���\��dj&�98�CI���i���uf�z���+I�1D"�e��L���Ʒer�L�	d�h閡`����J��V���P��B\��2����qc�����`�CO�S=�`ؚp%	���YKf��, o��1������K�-��y�\�uã->�T�����MPF������hb�~�.�*4i�A����	�
E���me����ip�$jؤ5Y�z*����m�j �ԫ3��|�q�lAд|�L��90�#A#-��c=K�c	��"?ю�g�3L�b��^E�(c��73� +�.��a�e�gdi�˶�,+�g�K�Q���� ���홮IB�ۻ�^FE6�w��_7����f\�X�Ep�Җ�0��^ťG�����X`�#�ɘ��N����ɡ}�6��e@7��0���sB���)��eOr�qt^�?Ӊ�b��(����m�UBȰ$ZT�l����m ,@ye�G�ٽǳ�v�ivƅF[%����s�f������0,{�ۘ����x�o�h�-�ӓ��X�n���h�3F�����S-%�NLSV%c�g��� ��"����&�J���s�Cw9/����Q�H�$��49K��V:*�xt�ƥ���b�$rg��k�9=����������hό Z��~���q��������/��t�9��������`{F�b�]��sV�V�TZE�k;2��r��E?���1���zd�K�Mv;{}
�Y�@�Yג�͝Xږ@�1��5���,Nv�N+q<3�c��vK܀�4+��ܲ@�Δ�8�	Zf����:�~������Q�[8�5���IARR�M�9u�8*�� H����ݰ��{�c�@-e�I��t����3:�c��T%�l;���w-Q��K=��Y�
?��7�5�ҝ���b=:x��E.�:�V�ǭIis5nu��I���h-7^xvF���R	�2�e��\'"+���J��STH�>���E�Y�L1�C"��ͱ=I6#y�"3>u�Pv2�����g��:������8��,�y���ێ��y�N^!Im)@�;y�Bp�r��;��,/��J&w1��=#g6F)��y�ܓA \�]Y;�oZ��r�8����|��ט�y1�j6}�:����V5��{7�h�.��"";��o��>Qpo �g�Ie��q5	-n0O�����R��!��A�=snr�v��%#���[�q�jAZ)����T�o^:��R���*���*�DO�-�n0_9�*?�>���Z�L~<���icR�� U�i�*H�\�7���bTW�磲�oC�uSOk�؈Tl�l����(
�� ��m�9��8��l����QY���#+�?��zp���3�`wNg� oc�Y'�Q]qB'Aft�5}r���rN�u҂2�%oy|��J�72m"�3ܐ�Y�j5�m��Gk���6[�����!�L�����S��e��l��rT�^�-�/�c��+%d�W]o"����=�,X�1�o�'�4��3+7���أ��9=l�27̸�?�����7v�� ?�l�.�q�}�:���٭"_��MiR������v�0f�&:Y�sǀ��1�k��;��mn�����x��#G\V����Y�Q�qj�ܝ���1����v������C�̺���Uq���^U���˴�ȹ�|w3��R]Ӂ��mSD{��n���*Y� Qq9W�����O�|T�J:��;�p� �]��&�P�X� f��wM
JYm�6�ލ�����y^�͞nw�6� 9���s��?a�J{�y±
ʁ�����% \E�{�������E2R�j,��{2z5s��>t�N�����>2o���-W�ޝ���E�)d�q�w  � m�β}��O^-�`���h]e Y�U6c\k����A];h-�4�z�����n;����
H1�D*�f���*䬷P#7���\� Őu�����o@����w<��e�Se�o�Tg>1汷N���F� ��P�u"�W�����e���B��*����ϗ���������m���O����6�a���:P��y��ՁV�!�Y�/�zR�N},,��W���?�/��^*s9 3��.���⺸~��k ������˿����ÿy~�\O��po� 	ڜ���*,�Iٓ��}�D��J�P�FW��Rde-݃�� ���w�r��.�%�����4��;S��#]�|u����8S  ���Q�[O(2��7Ci�|p�X83��\]�[r�����K� �\a?h�Ap(0�>2F�1U�T��s�|�@ ��P�F�2]p�a��yS�,`%��N�-/sN0ft�8�U���� K͂��)��p���ZLƝ�67ܫ� ;� @�)��i��f����H�rR��}h�$�"����eT �ѕLrpN7�%74b�ݔU7$���}����2��ڹ�	B)i�t`F��b�ŨϏ~�Ƌ�ч왅�J��o
������8�� ����s��UK��\��ݗ΍8�k�\Ѝ�5��뎚��@�I�]���u�j��v�:�Jy�2����ƶ�\0����bm9Ւ���EE|��J���s���˹��Z�	}U�O��
E�'�!�����_��^��Y�s�d��ΰ�w�$ �}�k�A�?0���2Ǫ4�妱R�utqi��ǎ�L[M�	�#V�*H�����}��|�YCS�9k՗IJ�[�nۈ2����<�࿟�r4���)QF����Y(���%�L)΋;HJ���r�S�3�i��Oj����� �� +8,�m�ʼڍ�NtΪء�@8z��܋Wz��c
��wj��>x�J���?�w��;��9@���2Ft�)BI��j^B�u��bҭ��o=�	}yͦ���~ۍE�z�M��F'wXu<���*�f[�nY��� �����$��@F=
�B�IVSO�1�
Ҽ�G���._�-� ze���� ]ze#��@??��x �\5��4,z0�{0^�lg��>��7o���+teZK&����Q��:���޻����ӽ�)���KP��ҺYPZ��V(s9����ʫ'ߘS@��F
�)�j�G K����2(9��JSW'^�@��������1����h_���q���3z��{�ν���Ǵ�T	&�6V�>&m;�9IA�&�i8oh���|je Q���#�����F�Z�%YՓ���2m�����t4~��d�[��<��o����wߡ��t:���ҙ�"���O9������Ui��_��M����r^����ljq�r0d������U�qtB����yU���
�і>�>��?z�>:?�����v�1�;ƞ�{V5p��1��b	4� d�.2({�u�B���^�m������*����p�iz��e�4��k�jT�Bv�!�/>��������O��p����S�d�k{������@�Z)�ݶIve΄乡2�Қ���&�1_k�a��kO^��o]�kG��n����u3�6��΃��g��{������jM��}����మ�5͕��(e~�;K�Г���B�I<�KJAv����h=u�}ٻ�ɠ�g�/�O=K�u%�,Bv�8[�L{c>~�)��/ߢ_l�|���y߈/��Μ2�y=g sW(4~��c � ��$v��D��x��Ֆ�e��
�y�_��:�q�������ݢ[���6
̱5�s����������?��伮�w��U�c| ���G��r�&3�� ������`$�Mp9z޷���TB�_����+c�_�v���~K  d.�'�z%��O��;曟�����F�b���ZA�|0gHȪ�N�^/�L����y5��Z���cO��J�I��k&+7������;dq.k��n�1)�����?z�>:{DC�юimܗ�gM�9�B[�ʊ�]���������L����6�Gع^iU�f�;��}�2��x�P��.��=}��|�]2�נmgӓ9ɼ��wo�g��g�t����嬽J�=�O�T���jG͉���� "�D�#ѳ\��s;W6&A����dm����'�}칫7�2`N���ܘ�Ӑu���C���c:�fz4Ξ$��#㑥���������@9_ɺ}�f�w�s��߁y)c�f~��:�g]lu:Ӎ�W��+w�&϶֊���n�,�;}(2�ݳ��1x����9� S:*�Q[��4�5 ��-����)"�|����Ӧ��A��.�٢��ve��z���[��x�)��0��@�{�6v�}z��+;Lv>����SҺ��d�i��c�[��g�G\ڭDq�I����X�b�,/'˅C�E��DW�1�K�!ƌ���:�LW�>=�
n��|��D>:�O>���x�+,�״���u�
��L�2V �����E��vn�kQ�1*�_3�� #+Y% ��&�$]���e�s���M�sy����m�T"&��������[�?�Ӄ�������ߤm֐����Ï��7Z�P������uj���~ˮv�ʈ�F���ܺ����5c@9'�n\:q>���W)(�\k�{��Mc����-�4�--�_��rI�I��y���[?��&;��������g�\|��Jt��f��h�+օ%c�C�>����_��/�y��[_{�h~8�/]�T�⺸.���W\�+ ��7rz�7��������'�v�/��s�����p�h�'C! @�l���{��}�X�9"
�Ӕ駞�c�$d�~�P�?���yvώ�(�]�?���EuL�5ݼq�?|K�1ؐ�Lj3<8����5SJU�Ձ��"/��=�Μ�%�W���������r���O�f�TG�a�O©dʼ@���(w��b�D0�{���ٻZ.���GlO7C�lj�'Y����9�UA��Y�22}q��4�b���@�R���{��U��ՠ�p�ۜ-N)H�����]3��M%�m�XG��ǤrO��w�d}�)yſ�X8��sScw�mZ����JB�xğ�Ep�F�"#�����я?A��#Q�u��tmg3���]�}��q��s&�z�Q��R�g�@Љ�ٔ��P�F��NXuE�2�iO)�\|; *��H�N�GQ�k��2���Η;q��'�1r�7���ƀf�MuZл��G ͍��7+E��T=Э�:Z+�V\Z��^��Ƚ$����z�;;�ge�XU~e-S���7zAƺ�*?/ 5U�'{/�Dz�ӶWz��fmN���m�\b_20�B�ۃ�)��-Xp�Y�C��<F���F9o��s T��D�3�{����H"|Ə_�|m��,+.�)U`,(�s�5u����i�� z�-g���|���0\���/JO��t�\�O�d�����9�g�1g�9�ȲKխ�l�)˚�OM�[:p�ǌq��a��8Ķ�n�}�:�W�5�i��I����u�Oﱵ����n��C�,�W�a��t�d��Y�ѫ��KT��r=� ZAn��I/J���.����^;SJ-�mxN6#�?���ѡ8�� Z�v�N�͊V�ӗoޥWnݥú�����o�ŝ�R�x�%�u26���mzm|����������S�n��3Y�
%�v��X���`-�˃��g>C�a�]s��n��mɄ'��l��ڪd+qV����d��z��o��*�>�B�s�@B=#V
�Ձs���W������`5�_����'����цs���3�&;�%���2MQ�Fǎ���W�@��q(h���P}Ry�f�ti����y�g._�/?�<][J&2;2ϊ�0 ��M~RVt��}��=$�?~�6��_�I���4YY�Yu�u�,��/>C��ҟ<G�k�~B���*�?״���I��R<8�>���ߠg�ޤ+�Zc` ����.O?��N �>�W�>�v���~�}����#>���إ/�v��Iu��C����@/`�'f�̹8�˳ȟ�Lh�5�L2�����>>'l��sG��KϾ@�8@pƁ�O>Z��2��_����Uz��[�ɴ������G�M����H"e���lM�N c����)�6ha @
W���� bW�Yf?cC\6��ڧ�;_�:��\��6���3,�?�ʟ�lg����c���_�MmU��G�п����o�((; �ƽY?:۞�̙,�;��0[om=ks
�� O��t?�L��Y���j�X$�5fpm��_���W��Ѭ���7�^*�zg��q��+��K_���D��>��?���H1���}�r�z�. ��n7[f2}{� �4��͢���(5r�Ҫ�Y�4(��Sv���/��ҫ��}m�MztN'�O�c��z���r�� �[��_~�槾@��L�����I��D���1�1O���WΪf�͜�*1�+�߸T.��t�Lo��et�3'u?��~U��Jpm��iC�1����5Jp�����L��v9�t�s�U9n^{��5����{�o��޼��m�fz2���WZN�l�@5]�y��E�e8l��?A��w���>̬V\B�3��;�^��;�~��^��x��`8�|�V	,^8P|��:�0��N���~�7�/��)m�^��ثs�r+�eyj@�?
�h�p��2�Ku;�=D �� ��J�Dpb�l�����[���_��)L��>�K��J�C���}~y�D�?}L���'c~����ƧR�m��s�r��ʘxj.' -y�R��sP|�Z�'�q�0u�r���2��i��#������]k5t�ݐ��T��ӑg�rۗ�v�߭�/Ry�K��O����uzg����1��,gb���A�Ղ�������j�P� ���. :�U�sG���g��RE�����X�͘ߕ���������|KW�M���k��,=�\x�~t����m�?�m�蝟���@�Z��|嘸�$_+=jk<�~u�CU�+l��&םp�3����U��k���+o̖Q]sK�_�E_~��q����m��*?bZ` �`�r��A���9��~��h��������=�GkA�l���b�l��*�$�hQ=V�Zc������|�����ib���2�ze�_��<=3ti���2�]x����V����鄞��E��V��Gп}�Gt���!�yꓵt���-��DŒ�������0�K�Үk��9���U�W3��^��}n����Ѝ��TG;>�xܩ��X�s|省F�.�����٦�>x���7�q�d��N+�Ζ-*&�܊V1�g��_�9l�HD ��S!���Ӑ{�է(��@Z�0��������A�D!{L������p�)��z���ז�UD�����}OU�+_�"�W)}S���6Kq�A��3o�*zc��|����o����F�<=j����ߝ<}��W_z�d|r0o)�rq]\������]@l�O��һ?x�A9}�tu~iǝ2%�]��6�P�|C���qJ��p�Bi/��2�^�[:�r���|�ï�7��k5  �u�Ͼ�߶*�A�������[���s}#9�M  �I�L��AЊ��Y�p ���75�S�+�|[� ���G�J6Gy��^� U��3Q�x���g��ǗZ�z8�ݩH���3�J�#u)��,��L����,�$z8]e��s���X�{Y {�>���by�b�Qk�m�P�����D�-i�d�`]#�]��[�yݱ}l��/o4�bWVgϤi�4u��_��@�������#�вNȄM���ۍܾ���q���:gpX5	1���s��٣���M����������n%۠k��g�X@�i�c������>#{)�L��e\XiZ�����S}�F���!`��j��f��,��,dv����x��p�o��.��"	8�CX�s�������hz8Z�r� ��E���q���R_�%�=��'QB�)�E2�4�Z�Tj������S磘O��������k�
�!���/2�?Z`1�m��2�- l���h%�e�"��\N�r?���s�u��"`�s֔�֚�7U��EH��:�	����Ci�4���� �&c���L*zl"�e���\A/k�0cY���= ��|%�)9��� ������3��η�L&@�;h�Zp��l@�3-�f��`_�/@C�<c2'��@��-��&h�w�?�@�� i�F���l���q���eQ��v�ʹ�����(��~O��x��e�|䭚
9pCޫ������*e�����j �?�x�K�>���-:���U{w�#[7��F�/I>"-���������>�ez��>��;?���iM���9�7Q�r��k/4>ˊT����!%3�L���KVKg���3��e�,��8��m��[�ܳ�í�OwV*�ٶ|��#�Vy����N��7��[/�wn�@���m��wߤv��B����Ink @��|��X8Ͳ�sV@J	�ّUGfGuu0���d�ݝ鈾���t���K��2R�f�t-=x���k�%���3�ƕ����{������[T��HF�d�I_���qFo�R�&k3�I�@�4�`�Zҿ����\NV�hc�8Hp|�襫��K_x���D�\V���803��4p� Z�z|�^x����G���Szp4I�h�@ەn�w�|�@�rbD��8_п�E���E�����҆�j �x���v�o?�%�^6�z̕(f����4n�9��4�S.==�ҍ��;W��o]�C����Oߡ�㍜��'	^�!횜�.��r�B�@	:��GK=U;M+����C�%k�AE��xi|���k���F����9��*FR�Í�
}��w�;���zHw~�������9��=�:��*0B�U�4�	,�\U9�cȶl'o7�JZ4���S�s�(�����6��W�v=����Cm� vZճ�6 �2�A��!g��N_[_�W��;�6?�?y��t�x��kO�aגV�P}#<&���A6�xu -9��/|��׵J���|��_�[���?�J�2�#�R�XÂ��$�����юn������n>O��'����=:��Y�}�W#A9k�0�ĳ͛�bgD�eѾG{�7�U�\y����=<��ݦW��1h��mC�si2�׿:k"v���:�Ϟ?�ҝr@�^�*}r~F����Ɛ}@�{��ca_��;gБ�� ��5-2��]��&�k��ǫ]9'��s/�'7�>:�I��)j�-HX�7���<����߽����g�ǟ~@���_�V�O����Bs���N{V�S@��WP�N�l]�fP4��y�d����a�|�5���恖�.8�9ھ�L� �J�f��@�i.��2-���E9Jӡ�X'�kR]L�`Q�Dg!�c�]�S��J ~�s[��ZD���Ttr��ݤ����!���<b�=ke���V�_"���DG�>�G�?��A����齳�o�#��H�5�e��ʑ�R;C�a;�f˓�T�S���*oH�s+U)�yWʲ�W��T"�x����_~��е�V�\�i'@�:�?�2�)�����[�>����g�����?zW��GGG�������Sq�c6���g �J�M@_�H�
Z����N*��dz��5������xz}H�����v�4�`�	�(҉T�s��f�E��-�7��k��|�l��?�1���}Zm0и�Ѭ�Qia���Td��<7�>|6T��D@Z�� ���B���<s,���D߼�]=<���  ��IDAT�1��#�,!UdHAR遴<�N�F��{tN�^���ߢwOҿ����A���"@�U��
�W���zE	}�v�-`���a���;�{e��sRIh�p���|�%z�\��s��u�}Oj�ߥ<TA�C�]���7nї�r����7�'}@��+z����L�$>��#a�j.����p�<����*u��)H��AU�P�W@�*|槂�K��"�������k�P�U�O8Q9C���WV�\X����.�ޛ�K������Oz
&!�B�Z�����v+^���9�O�v=|�g�is��<�<�G�v��僃aFw�|�hȋ�⺸.����  �Um��i���.����G�ƪg�#���\���p�,���Y���+%�N���Ɗ]��H�V0ޣ��������x���ҥ-=U��j=Jf���w�RA*&-��̝(�fZ��>Kt�!��<�z(�u��,�@��(�������s�p�S��n�WZ:��A�tI���u܇�M~6BT�b5
c�#C-��%�fP�=�����5�Cw|=�\k�S�k�@��%��E������WQ����m�K��=��gǖʁ��Td�G� 9M!�q	{�w���N@��ʧ Cr�G����hb;4@�����=�Q =xB(�X'3&p��*%n��]�*�����k��7�FSXkTp sr��� �t;h-��:ȳ0r#r� ���dqˀ�N�z_r�I���H 	9��h�QV���Z;�:v�����G��3@Б
��l��U<S�$:��ha_��P¸��[7--����9Z��C���{&)^�lH�2�f[ۊ~t��4%$�|��p�@Ҵ�Y�4Ap�E�`b-�͗1� hJ�p�s��<xn���V2�����<AJoY(��9�d�VʱH�γ�A?Q�������}#�H.�Y���5ޔi��@{c�P�l{��f` �L�(h�1e�y�v4�6z�w�}���{h6��}8�,+ӀW��T5C5@��EB���)PR����^<|a�v `��c�;���TtP
��ZMF7	ĳ�H&��|:�ѳ���qN�
`B1����^��e׹ؘk�O�s��9tUuNl�-J�hɖ׸���a~���~��'�~r�a�5���*���IvS�α���I{����s�SMIDI���s�k�0��� 5��>G�(Ø��
�O� Aؚ^��/�R��A��5)��ގ9���P9O!*�y 2���;�b�Y��������u�#7ߟO�m���N�Rߊ��Y�ܘ�d�8}��)�f�c3Qsgc`<��R{��.?Co���~z�KjZ���4�`h �-�;r	��:c	zD�v�h��{�A�e�:;�灞=w��-�Q�E	��U.��(�	젖���A�06�U�V�`gዛ���������}6��|a$=�e��h�2ZI��B�E���ݿnףsl�T��s�ɿ�ׄ���4Iņk�'h��~�)�6ф
dc*�3^N��9gX�c_�����y:��N�Λ4Z�H��伥�:*�~�wM�^��e찬uJ��`Rp 9P��5���t~y]��
/ᩩ+���U��d1J���	}80r}�8�]^�7���>�ە�̳-�J���$�U���DC^�s
ƣ�O=H�yo�����˳DWW7���ZKc���3��Q	�� ,s���H_o�>94ѷ���KǷ�{��>�2tڨM.�&Т�K��R3о�� �`@1�FT�k48�?2�G��������tf}�FS.�=Aj̾�J��ѫ��n"'3�Vd�ɇ����O�B?��=z��i��H�������g��7dq�W�Y%3�XV&����6Y��-�W3�<3Y���\�Ͱ -D����Z澃zRT~.P�)���K��ia��s��ަ�����������<��O�Qh���xX����F�W �}'+gl6���ȿ-�}k��>~�Vz��a���K�wk��g����`��{����%����W���	���������8�dX������\���( �ˍWW������V=*�έBV�l���+�3Y����R� ��{�g����gH�bT�,���9��%:u��,�>�?��m�����D�b��_��t,:X����(��VvP�k`��`,Fr;�K�U�ڹ˒YY?YPILE�jTo���Zҟ�MoR��j^�cy_^=CWolџ~����>���d�d�U�G�<����F)�O�g����^��̯���xl�]�|�ŝ�tu�8�΂T/`p",�M�ʹW��U�X����t]��7�ݢ{w��O��ܿ���o�&7^�`ա�u !�J�?�E����X���j�7��ߋ���7�v�2m����`�q�x)Q�eM%�^�N�Ϋ�A[����+�T˴}�y���w��4͟�0s�A��gXp�HBC����l���Dt@1�Bz`�=��9���`���-z��IZc��1kR)x�<f_��&�Q (˿�0�6�k��e�׎��k�gY�<�~0�뾕�Ƽ�1^i���\oL��]�/Ue�N�7��]���Y�Z�Fz*��˛'hi��3UB��ܩ~��R�4<i��Fڼ�<��<���o����ӏޣ�q�W��g- ��좡�(��Ki0x���`� Vwc��D�7�. Z�L���:����f��\�n�K��9��*@����v�E�6;���(�\:��rX��[/�O����ϩͺ4�<i	�*L7�T�����#H{M�oP��z�-�����f���|`./oГg�9l�*A�d~��R:m_�청�W�i���i=�k�~��5���C��[t/oꞜ3�x3�)8U���@�x���t�0�=�z�w;9��$������9�c�����F��6�ߵ�viiqq���R��ػ��W:r���#�$JI.
h�h�2�A;]��ŧ#��N(�\�}Hh�`|3u����Зז�p�����������ׯ @��gM��[�,���o�y�܋P;�)"���ìO����ʸP��O�@0�6�f����K��)�G�D��&��MУ,8z��<�Z�R�!/��d���W
�1(J5�$8؀��Ǆ��<��L��\�ϩ��2_@+KY]|�7��)TZHP_�`��}��*�Y�ME�z���>C��a(9�k�`�d��"Q���g��3A�ģ�����<c����T��  E�� P��܏ԑ��M�h��{�^|��ήJ��>@up[�W�3����xCzIU�~%�eY�0d	e���D��e<d΀JWΩ:$�g�Mq�@��_;�q{���`�Oպ�˾�7=QɆpxҰ������?��; 3(��W� v��A�KV��4mz��Z9�~��G�K�-�3he�C㋍�{*�4F� X8��Wrc�X�\ɳ������+���G2D��碮�:�J�q��)X��@��eNà/9_Ҟ�Vq��W(C	9C�
b�֎e�(U`%�%ut���*�-�J	��@��u�^�������:�F�<��tY@Eȕ�ۅ���|I`�4B�3e��}�xƐ�<��[��l� ^I[-�j>-��p/Yۼ_]g�|�J������u��c<�������Z��2�^�a�C鿛����Z?S�e�eOpڶ�����wSb��@�,�ײ�V!V�I�d0��)H��I���t6,���ñ{���A/`'ZK���ܧ4��~lCy��1R����l����y�=R����ǐ�Q���C��ӄW6�O��<) F��TXq*�g���w2��W!�$����u�G�����fcz:��9�t����9��|\J�fE[z���Ul(#�٨�d��Y����q r	�8�������N��臟�K�$d[A�8���q�&T0���-%�m�m�k�+��c {Գ��1�8�9���h�]�o^�F�=�uCFTc�^�괱V"yMFr�Ȃ�z��9+�L��wtn�H�w����ߢ��{��<��nչ�����u��J��87������cYU�? X�v�om����OHFN��_��]��zK�nLWIJ�l�4������r>��k��������i�W~��h{�w ��7F�Rh��r�#S	Aִi� ѥ�H/��,�
�.��@=Wn ڀ;�g�����J�������{�]������w�o�ޖ==�����{� R}��.�\�֊��	𨏮G�5\����a�d��5���=q�ff_�(�M#M8�YX�䖬�t��စtTi�LF�J�zFgi�~��S�����ޛ�ӃIu���%��4 ��@F�ysZE�v���ɰ$�n�,�W��8`���[t�Y�v��A��wI�������`�H�|��Տ>��ί/��������������-���8�s�h4]ZB�Q��� �>�λ��1 4.�x8cp!��[z��=s���$7Ӄ�VX#]vv��-6V�m���:�=�%:~�Iz�����/��l� �F6Y��0Tl7�m�T-����3�]��>�gVo��}��5:7^����H8�i�gQ�>!%�-��� �Z�
l%�'����
�����O�~��sz8֌dnGp��(�n��&�F���a@I�,��K�N�eBl��h��~�d�3h�3�e�*�Y�J=��d�#Q��%�ݲ9'g�vy�zzz�4���\�%}ɕ���P�:|"�sꉲ�澈g���&�i��j�yc}�^9y�;��> |�5
��9E�*���a_D��/}FO
�����I~�⓴��[���w��;��Q{�7 H7��եD�Q�Bm��ե:�F�(�6�I�8���z�]���8iU�`>ݐ��CB�ڪ�?뵭�o.�=ɓ�v3zf�A'.����&����Do��,k��Z�raR�������s*`X�J��"d�?�����-zj딵h��<�F��&�X�* Q@XRI��r�`�h[���s��~k�*����������ƑT���J�������������['F���4i�����ｰr��߼@��L���\�b^����vHS�Bu�:H�å�HP��¬��Y�_���[?��C�i�wT_���z�_/@5���4'�!��{i�&`l*�-�[腭�lߞz�����Ni:Sm~�K��stѪi�9Tx�V�!���K�L^���V��C�N�yhe��ɐ�������B=�����]�Vb� �q4�G�>��a�g��Е�-i�!�H}*XZ�%ؗ�Ţ���ܥ����.L�κHVb�4���'.�N���;�pe�e�Ur��4�Z) TH�om����S+T66ӱ������f��u�.o�zZ�s�mx�Z���A�B�%�~ �?)@��Ȳ��:.N�h����Go�N!̮�{��n���X���0/yU�P��:^�,*}��jfd���$'�������4���~���J�Ⱦ�����|.��)`pҜ��},��ؒ��@F������I*��wXu���DѮ��Z֗g�-����z|=�_��� H'�d�����ŭ��>���Q7?��1M[��u1nD�zs�5��oMQ�gKp�S�8w�q4$kR�2h .�Q%��e0UP���9T�,�$��� �߿|��+Xf}��>"����nd��w���綣��6�8+S����������`��I�0�Ygg�\Ԣ����4.���o�k5T4�V2��L���6x��N�JԦ����w�<C��}3CÜMC6W�݀0C�q-ˌ2��pA�{O�G������0��|�Z�JT�#3fu,���ggbA�#��q$���� �3��? X�>�����@�N1���"�wN�
4��0@?f݋�m���*���Y�Dn�(�3~x,l�����Z1��jb��j49T��9P��}������Z�u��(��s��?�`~oY��������\�ƚ_릩>oc�0�pzl� q���=����Q���� �1�P2L�����|+�R�a8b���9TO��V֣/�7�Xr�Ё�,`�*@ Tpt�R�lܒ�Q{8j��+�?Su`̫���?���fʣ�ʟ�Yھ�-t���|���%&GݷM;��}�����d����x2',C6'8�TviCk�9��U�R�/�\���I^kpv\D޷R�)yW��l@9{��m�~x#D+^GF���z�Eq ����f��7A�Ö��e4�*�c<��@!��O�\T���I�A��Q@I������C��@9��Yj	�Nn5�a���0��{��c%�B�����t�e��CP��"Q*t���ynLN�� �5@��ga��5$�^��؃h��&��rF��S�
�*���r���} lSKЪ��CH��Z�3YJ#k#ko�ʱ��RJ�R53V禱̢�P��v���F��w�Y ���G K*-+ϒ�7�V��渇h�4C7�1u�0ѫ�����|�T�j:s���	ЊC�RA
�x��ى����,
�ri�g��ha��?��!�4*�9�9�(K�K�e����od�	x���V�AL�p^������r3!n|�{\ a⿤�Np-�7]������}�F��{���/~D���6�f�_���K���q^��M`�Qi�ɴ�f!w��D� �$��$��Xާ�]=K�6�����9('I��z�j!^���\Z�Y��� �|���k��߹�������'ڟ(D�VY6�V�/hB��� �W8g��֝��yM��]���矐Վ�G�����&X�\�?�9&�L�@�@��L�L,} �9���C;��~�}��v+Ѿe�02V�Y��P�Y�~d:�	>+�܎#�vf��Mb#���v~���:=s�u��|f�����>�c�X=���Ѐ�X��le�h���m!~��4y��e�G� U*�U R�"
m�V~�*)���t�j\��B'ɔ�I�Ysۇ=�ƥ�t<��jhO��%Osd6~J��چ�좎��r����r�i���i:F����9ōV�E̥91v�\�z�A1�5��-]�X�@N	Х���C�0�q�ۅL7;y��{��9Z�j�t��k��u������s-�JPX�f��l���='z��MJ?�^O�t7�g���G;P��W�j
x�8��no��qF��qF_�r�aLKyn;yNߺt�NOV���A��������L�k�|�g��$X�r����o��/��է��z�>��s��@g�6�eA��-v"��=��#;nK� ^�yj4���H,�:Z�2m;�߽�$�i��y�t�k+�*�RZ�P��E���<,�n�<�!Xܧ���}���G�I.%M�:P�O�Zɑ��m�D����u���}L���omA*h+�q�WL�����n��0��d��7]�L_6�-cH����%�Y��	̈��|�H���J��ޡ�|*e�����U����-��qE��D�}���C�3�z���Z�)��.g�X���ۧ�����S��$d��� ���3&�a�X�5MRj��*�K���y�'ן����ߣ���-�19 "��2�n�[/xT6��7Mp ���m%شz��y�k�>_Y٤뙯���7�n��� i�K�8D�����~�~�2�]��\��0��;C�ޔ~:�GI3�����4�K������Wl
e�T>W�.��D�s��b��F���'������!M����0]F�>�c��i_'�Ƚ��B�M�d�2�����\z�����;�=�?V>9K��>��h�6��N5�d�6��#^PF
XV/g����O��������&ͦS�����h-#�P�ܑ�$�aà��1��%�(�۬����p���O��J/m�Xߛ7Z����ձ#��k�NHJ�W�Qk�+�]�[2�d!��v��+�N҅c;��#�x���B��7�==�wSl��g-P?"�Ëy�77�P;M��ߣ��F*sX��zg]a����χɳk��T壀��#K��4�P�b�F��?{zoNO��D�׷�N��̽ǔkF���26��*uB�-%`�L��2ec<�o�x���ߧ�6'tT�I#�\�v����� (�ne�1=�^lr�x��t,�@|ڒZ`_Aʥ����o�,k�31{�1��yv����V��,ڳďf ���_+�[�r;�Rᾶ��)/�?��:��+��"�)8F#vl�M���Tw�J-#:�5��������+��hE��y^����O�tx����~��@�z|=�_��G�_;  ��/�=�o��~�����;o��M�R��>�F�*��J#_.�Mc��:iFejF������ʞ,5^!�����ב�G������@�_u�_����BF����<'��T�-����DJ�`~ufY�:$x ��Rk�`�����E�(NP�Ϙ�a.#���؈ɂ��2t'?��͂l�J��Q��[�M�d�%(m��F�F�Q�� �{$���+22xA��X#�Z+��5�M4��*Gf��Ɲ��2�=*7�Q�_��?����d�z�F[єl�-3�c߹R�Q �pUAr*ʢ�h!x���%��}� ��.�� ��n�� ����
��%�#�z����D Z���e\��}*g�ў����[d�C�Z_��Y@Ц����9J>�����{z��o(=�@}�7�Iǽ��E�z	�U�2;�@�)�%�N��4U�= 3�>����`#�+Th���g!`��7�a����അ��F��'�Ll�ƒ��2Ϫ��>Z����a8�0b>��o��L�P�}0ǝ~�ny�����g���XӤ�^��%�Y2{���?��#{��%��΍��h�A����g�r���:�N0�e��	�*�~ќnU`3%���[!e���� ��@��|6b+U	�3����s��5�GV>�ȍk�AF+�O/�}��5��4�T#{���p�D��,�>�t!e��Q��O60�\t��	9�� 1t�[����0�T�u|zF�ڷ��v (� ̀.ɜ�Cy�kT��P8nh�unt�lh�	��Sx�fp�z�܉%�BP�A{�d3�g�T���y�? ��@��8� �
 ��-y �V���<պU{�)|�M�o���ء;� ��W?�ѷn�H;q�NA>�s�k�ƀFZ��GTζV2i:���Ž�p���Nї�������c��*Z���'NL�
t�#h�چ0����<��J62�����q#k`k�J[1��F����O/5=g���j���o?�"��~��(�J��Q�*�����@&���͐a8jN5�����dK���g���:��ޯVzwڈ�D/M���Uh
Ady�����Μ�M��˷��z�fm��mz;��/Vx%��*��s�ݤ�c��#�46 �I��������v�IZ�Ϟ�s���(�,A����9�Ϯ�_��/Кh��񓴟_���#ڛ@�"Z��&����LFכE^q��h=�c�;��x�����z����pW{r�z&��?�s�c�r�MdhBw��'�Dr��L߸�,���?��z�!��1��0z��|��UAU����IisA*�������<���ǔf�@Ұ�
hT��d���TP2:Q���;����hH2w�m����{�)}�@�ngnN����5�W����g g -��k�88���vc��'�o��nP�=��atX��Ѽ��9R��F�l/E+	�m��3϶�˷��/~�=�.�R��N���U�9U�!zFiU�r�OV�>������>�������`F�0�=�쀴2?�C��3=���>�����=�	��իO����O�[m�0t#�1�Ӫrĺ2��.*]2Z�u��E$��t���-mv-}��(>�I9c�?)�"�e����?��S�kЩ��l�2K���ѩ�Mzr~�vo�O���d�ιt+<E�=t�nq��B�c�!�����zj7�	��K�k���Aw
�@�[_�M)����J c *��&�-�A����H/\}�>��]�8��5���gpI�刽#gی�ER�#.&��&�s�@e���矤�+��J�(��]��4����9Σ��e����������:��g�@�`<�#M�ly�VF�L�xT;� �[t�
<T]�A?O?M�wNJ�>hy��(��s���Re��2ь� @����q��y�����M��ۣ{�_l n���?z�G�T*O��K �=i��6�*J�W�
0zz�4=�y���]���L��a��N*ۀj���!`X�ia������ҵ'��kߗ��������h$���۵�]�?n$i0\lh
��>� k�sv�of��W��k[��^t� ��kH������Joҵ�^҄"mC�J���h�^�~����-�f����*0D��=Z ֬:������j���WZɺ��g��ٳ4zx(�`l�xf�G�L���g��G,[i$v�H�z�,}q���d�D^v�D�[�@ŧR+��*[� @������6��<w�έoS�ZBX4�nmQ�}�h�=*�'t؏�k�H}�q6���={�&�~��W�W��Ƹ�D+?i��6`�C����|���[;�w�r�Q�|��� ��\Q#���YW1|@ɏ��q�iF���յ�i8&���gv���x�ppћQ=�<	FVk@�eP�K;�h���<��4$=6^O��|j�����^�;�#6Mzz|=�_������� �W̊���֩_�W��}�_�w���nGgg��F���W~l������h�}O�Ӕ����!D�2׌5�Am�ރݰ��������[SQ�!eퟩ?_�v���k_��|T�N��{�>�yw,Jj�ϖ�𦸐���pdL�Q;�f�J��R�����Op��A3��|h�`���:+��#%����g�4�d�a��l���#���X\y2ݾ�F�X�R��p|%E?��(
���,�'���VM4��N�����)�ќ�v�m�~2�T�s�B ��M�y��7�$>9�T�Е3[@���@������+��X_S,�HT�d�`S��$N�a`�Bd��Obe�U/�g��A�R�����88��n��Gu<�AV90�������}<e����ؓ+̸��w	r"Kؿ�����<`H_8��k����n��y�YTZP���5�N����r6�6J� �m���+��c<�)~=BU��j�Q��gZ�o�l�؉�e%�Gp(�����р��l��m�0$���k��5i��=�LMq������~S��T�=5�:X$<�}�YHBIc�%*"h��0�@�`� ��F���G���]�H�B���S�A[���Rs��)y�B��G������&�.-,�����jK���ز��������@L3d[_S�p�E���t#/�D����XElQ1�m�� �P���T�g��x�@�����8č��{�=KNs
:�`(:ӊ����gK�"�@p'H*c/����@(�=���)��D����`��d��>�С�&���2��	��Uޛ�$��LY
3�>Z������ ;��@QPC�mG�%���{z��5�
PJ��\f �L,`L;��;*�-��'�&Hye�#�Z��'��_���\�yw�R��'�@��z�#��|�����P^�}P�iƙR��<��/��:-̓�x6��;w:�j?�����F��J�NB�ٻ��;�ړ�G��L�dB�P�J�Vh���u��� ^�J�7�8-�z÷N^��k�t8;Ԁ@]~zy�qF�IW��u�Ŵ�A�Ʋ�I�v��1�]X���^��������!:g/�Ò�>�T���a���K�GʪZ&�$�15t|/ҫ���e.�����	�9[��,�����Z���˜!�T���q��߻q�4���z��Kr�u����FyK�,����ח??N.�:Y��_�A��Z�J�8qH{��j���zz-�xXm�JS��^�i>���'_������KlK[�����E[�!�H�uʻ��Ie�d4#�Ǔ��]�v��K�h{�H����q�}��*=�`���B��>7��ʋ-	��<��._��?�Rj���NrI��ւ�亝��J}�v�
�H�r�t1�1� ��aO������ك=ɂ��)�uTg�d��Gu(?�n"�z�!c�~  �Gtj%���/�����_��>j֙d��R����)�.�{���sH�wR#��D���tmk��C�hF_��_F�ӿ`�#c�(���B^��<�q�پu���w^�ny$O���3h�+4�ME�:I]2���Z��M�3>ѱ��~��gi�7Z�q�`��� ��H&6�?-L���I�n$+��>C_ܽCo��$�,p�?�������E�C�,@UR}��XO���2����?�*��<��r��M�x4&���ʒ��O�ҵ��������H���7�y����8i�;�_�z�Ұ���x�FЪӼ��〸T�!����淞�8E�׉fs᥽�N7� �)g�9��S���i�U�idܭ���'�"�x�����Դ5��G�����&��Z���LXUӉ��;2�[��|ޞ�zVt�6�m�i�Л�W��!� %����|���Ng\�c��^����7�rѴ�i�& ��-g\Gǀ�*�Θp�%����,V~}� �A���o^�N{�w����:տiY�8K��d&r�{�;�s�J��4�d=&
h�����-h&;�T��>��%B�,Y;Sckƪj�V��*:]�S2�rO����~��M��q����(�:`HTfܮ����@ �۴ ��U�$���d>߾�,��Oߤ�k!n��:@/~*vU���;�iE彴L��Lg���=u�<M�$�#��ֵ����s��-UtEo'�h�HO�y]���Kt�J��D�� Z%s��"�A����K�`�k/�B�h%;;��������-��|�4���LI�.��l��˙�J���5�����Z�+y�N����ܡ��}z��Ajӑ�<���h�	��".:=���g���G�'�5Jk�P���!��8���VE��2 #£����ݽ#���J� $D�s��n���ӊ8�{��W�8æ[�pRہm��}�'Ⱥ���VM�5���b�:�֋߼�0�|�e���E �=�_���ׯ�~�  f@̰�WVv����._��ur�����N�E<�|-�?hjs����so�U�ES�*G
�C � )eZ�jYPh���oL�܀��u��P�_]�  _�_9r�_�Z8��g���O�����]so�^�|f��b!�ۘ����g� ���{NQǵ`cU�G![���2�QK��֮��g�Ԣ/7��JIi}���>�2��%	��*/�$(�����6�ft��kC?���U�U�D}�������	F�+ǆ�YM	D�%iƦ=ȃ IГ([�E�G���R�ЮJ��lƒq��\����#�
�~"Z��z�K(�����3��s��]�`eLu���q_hgH_������6�=��̪�T)�F��X��c��c/���w������e�k��sa�{�ܤ�� �5G��C��9p��&��o�����]�`XY~}�f��x �:;de����-F�H��캑�6S�*Z����J0
�qh��ʲ>��/����s�g�xR�]=E+��r���L�  ���:�W�h��pt"��i���Ih ���X���m)��s�q��?�6�{/[m�����
��וk�ʂ����U��ݎV�0�"�?��Rqd��[�u?k�0���;H�����@/x�����J)߲�;2���qiEd�B�ܪ�Zc�ظ��� J���qyp�������+i�_��k�"P�� h�=�3P���5�Y��uF�p�{ کu����dsa͊3� �zo= �PˤO��Ѐ׫,?�4�= OԘ\���l�t�]Z�  �����&��n�mT�1�״�e��%�A�L�k�P�E�(�t6t�%�x�d��W��5�
'�;<�y� ٹ��]��tk�][ߡq����i� U�L�( �������7%T���z^&VU��=�z�&��ۯ�l�$ ���Y����jSFoL���*She,�}�=Y���tli&c-޵6v�>�Ͽ����/)1����9gE��xA�������h��G4Gq�{5��B�n}���������9�_�(O�������\��dq���%�����[;�L���R�����Z�T鼴y�~y�6��,Ӕ�W�ՙ��:�.x�g�@�:��hM�I���� ��B�k��;��dk�ro Z��_9#� ?ί��	�~��^�M���t�I ��܀�5��T���Ĺ�}ؠ=x���m�-}����Hp\J�K_�(��lQSx6d�fl�^���g|V����Z'R`e�H�&kt��/������D�wp����@��ƚ�J����^��뙍�ta{�f{��8Q�F�5�WTۚ�IN��J��m4%zT�cC��s��'��O~�=:\����Ij���] Xy�BC��|V�kI�|���F��SOS�7���$:��DV�<8(�������hӲF��V#�H���"��8E�����%�}i�R�E1e�i�MQgt�}Yk^�������^|�:���u��3���(c���`���MZ�_M�>%d������>�[�=�u��j�m\�ld��$�9���τ Y��Ǵfd���g�^{���CƩYS�
^!1T �J��~֋�g51��)h�ʹI�?s���/=A��͏h>�Fw��s�	e��� ��R�L�-�l� 6(˹K�:��_���@*t�<k�.���ia�0C2����IJ��6g�
?���|߯_�N��ԏ��8��$�c��"o�G�XC�޲L����@�u9��Vj���W�����ߙژk�&�)�Q
Ptt�I/ZA#��$[�t�ĩ�����i�{@����"���+�2�Ϥ���N�2o5����F��.�;��A���ۥ�^E�p�8Y�9~��j`����yeti(e�yL��>Ϟ�H�>x���#A�
Dㆁ���s��[�D�a?:����wne���m��>���@{W��%�$�a�U�"l"[��x�$&=��FW7N��{���(Z�?�P��G_?���^�/cQ�AҶ"����St㤶a�s6Am8[q�Z�P��*�]�|e��Ó&@4�Kq�m�K��8ӭv��r�r����!���n�M�Zɔ1u�+m]X\���\ʺ�T ����B��}�U�,�o���o�Œ

���"�:u�>��.�w@U0��D�R��qJV%Ò��i�����m`}�L?��ݺA��\�BI������m�6�ap{
_"��h�����_��8^�z��{�{t���p��i����#���_���t�q����h�%�Y4=����>�UgM��\7��т���>~��H &)��=���Ãy���׉8�3H>�'�j@S���}R� /HR��[��Zve�Qu�.������,aS�}&y�QFaqz���;���<�y~�'�����z|=����� �/�M״���ݟ�6�N�XT.�;ev����w�b*p��G���䯐�����>��u�"�B���� ����Bj�3���y�;�Կ���_�������������\a�L�ZV�#*A�������Қ�����5�f�V�A��d$��0fS4=��Ȍ�b���ʱz�v���&���6b	l�1� /[��(:a��G���7�!��������
�["F��T���
r�p�(�ʴNN��KG�e�}o��z-�2����C�[��4/ڢ�+�oncs��6p��a�e��`Eӄ}>W�9I�а/զj�P�'�(����b�� �+�z����UF���^���2��8-������(�T�ѫ����2�1S57��¥YT��z��H�,ᬓ;a������3\�*AL�it���#�8���}��<�Ie�	lټc��C�!�����H �b�q���Y�������G�ʂ�pS�Or��AlJN��{^�u�`P}�Q�s(�H Fi�>TN��8�T���� �z�A?���(%)����e;�(l��ƺӒ��zZ��L�>��ٮ�ա��Zf:C,kqF}�T�/Q�����Ñ�-S�j	�3���eC���Ϛap5��<�����`�q��9�pnPJ59h����7ΐy�V9�t��4�w�-? |?��@���~���^��@@���*Y_1/G���-rSѳ���|]}r��m��i��0՞c�T&E�N�t�^ԓ�Dm3p��,	C���
#�d�7Ƴ���.�#ߩ��A(�����@�T�j�^(S�d6ʉ}��6�4(��b3�󾧶5r��@�sd�q����2=�s�&�ʘH%�qŦ)�}p�B?�ؒ+@J-�$�뜺O��DX�k'�>��Z�����p\��%�MV�^h �"pe�/��m���	d��# Ա�΀�+1Z�=�^ѽ;�5�G�7�]�zO�6O�;�?��X�u1M�*@2������	z�͑+,俾s��F𫷊<��?��pg��S�I���L�W�W m�^�,�K����ݛ�s�K�r�?Ƕz˪�:�.��MC�Z�d�&p�o��@C���rl�z.���y�iF]�"㿂Cg��s�/xYG&9�s������|���C�7QQ�g���b�<���Q߅���f����JRP����TP��M3.�,��oS�'].<�O ���s�������7�Bz�j�� �M��V-�[�uȸ���E�I{�nӄ^�|���C�G4���V�P��ݺ���67-\.Q�e��m���pY�fDWV��~�%�[�>�hv���
#
O�Oc^.��7*����K�.S3�*S��P�����0��\͗�����,�y[�N[��BS ���mz����	���qh� ^��`M�e��AX��@9v鷞}�Z&����P��L��Q*�`��i�X�uなUi�Mn����F�d������<��y�mN���e^]^ݤ�Uɶ�>��{Cp���t{��U*�#��(e�5P%-�2��c��eޏv?���i�$�?�P�,��U4�J����+а��B�+��S���7'�}b(z��^W����n=�Z�Sa���r���6Nҏ>z�>�S�5z��p��~	�E�sgAG�D E0}�9^�'��ͧ�a0�}Wۤ$ۊPXk�����^G�+�jqh��,�3��8��3g.���~���y�����9͙o$��EhEA��]����y�/e}�8���T��X�����[ Zξ�T�a��b�J;]���A�����Ƕ���v{��)RZ���+� �Rc~�TtC5�{K���0�������'i)����T:kρV@�����
�tW�E؋8��˭��
������u�"���lc����������'Gח��#R ��4�K��R�)|�e\?`:r�[4p����kA�{`�y� 2}�e�42�z�s�/�_�C{�M�Ӄ�$������cP�U M +2o�Ϟ:+ ����;���ӑ��G֊��'�;C�2_�
�)�nNWN����o�A8�@��U�Pg��<*�����a�M�����+]���_`�(�]u� *��\�4��]��R*�P�1�"�j�@�I���xf�<=x��T-R^V|�_�����ɗ1�sQ^e�e��͈��mۀ��\ѫ�E���z��lJǳ}]���ӑ>_����ባ@qF{{�h�]�k����#4�u}Ͽ��e��@�Ŝ�����U���n�aʋ2�ܜA��ͷ���֗4��k����?��g�;��ԍ�z|=�_��_q��  ڬ��Nw'����-�Ҭ}�+3�z�gf�x8=�>kfq�TY��JP��H�*�|�p��g\.�#���������B��0����+�-�Y�������&� �g:SZ�DE0W�M.b�`v�%	��&A����8������V\8��K%[���+&��7�UM��7*gN	��xI�~�Ć���_���x|����y�c���d���,KM-�Ƴ7�IZ�e�=C�zN	�Sq4�S��(aJOo����]u�ȑ2�Z��*�4�W��+�c"WVj�{�K	>���hk6�Ű�T 	������8ؚ�~��O_���
��7k2�TH�v��~Jh�LF"_�����W���C���,��[(s�Z�
^+ip
A�Bf\���~W�mώ:L����h�GF�kytuh8G�l�ux8_�l@��r�
��0��G�r��d��,� Q��9z�xP�d�)֧Ҥfr+iԲ���bʵ���*�t`T6�(�jb*඲�G�U��;����z�6�|CK87��=�mF^D/RB�	�
+��f��7�f������I�z�#��%J,㕡;M�]-�*�^��ȝyJ`��ƌ��dM��&߯R .<ȝ�~���>�H~�
�/��Kt쵌�����;�!������w�N�ㅮ��nP����+4T��2n{�ٚ��fN�H*N��� 	���\���O:-@&�>|&�Z �	0��p�z0| �P���ZF�J�<���/�Ω�.:]�>G�01�j4Թ@Ȫ��m�m6��-t�M)M���"�4�h ���/+��.`�h8G�X��"�Q���`�+��%����$Z�={�<�Y?tv������2��WT7�A�C�2Nԕ���M�i��g���>K=�C�q*�[v��]�c&P:���=,�36�i� n~�xK�:��RƖ%I+A0�v��:�k ��2�[�??j��8�h#�Ɖ�t��45P�z�r�y:��CO���s ��:��u��ǖ橓��]*�e�ۖ��t����i�)�؎Rc Ed��mG��/oЩvI����<����rY_���D�'*Y�aK�z{�K!��7.^�L�h�y����F�%�G�<h�F��^R�y[�k�����%)�������?������5�V���+pIvs�hT[����Ü�������ty��w~��W}rz'�l��[�y��� 00���4�	c��|������
�����G ��p!�\�n�K��Á^����+�R���L�c/����
��������Ӱj.l�<4�Z~yOZ�����ٳ��w��,�9��U�C��mFʣ�mh�{�-����%�N��ti�N��Ҥ��ט��;�OR����\���k&�d�yI������~�~��	�?��wԊ��
�һݣ2��vW��J{RM��p��d��/��s?���ao
��<��(E���'�k*`9�L��ie���	�|l�~��S�'*�Z��U@����2Y��SR���c[ڛ�ׯ�|�y(`��(��@� �{�N��������4�Ԅn��7>��`�O.��3�F07eQ	�[�d4a��3�_�i&t�䙼��ү���k�p�����S{��|/�ϨYBI��蠣�;g�ΧoӬM�������_�|I'�hr6���*�W�xl�6���� Y��8���Z�۱Wd� ��~)��VI@��1y�Y�g��ѩ�*݋hz����@�䔵5�����*��#z)˼�`�>[�������
����־?�E�{T*�a��3��n�<O��M'��%�_M
�WS5�"ב�����
�bp�V޷�+���:�Ix��� �.�� �a^��S�CU�P>���,T�Y�_x"�Ϳ�wM�LR�	K�l>b�V�F����CŢ�A�6ʲ��?u�VFc����lTJAV���T{��{�ZZ(?}��V)k����Sg�/?�w�L���t�١�4���{�XS��M&�i����t&��e�̕�L�6ax��k�N��ϧ�h�&S���&�)���u�d������И��9������_&/����ma�ۦ��k�w��1�B�6X��j;�
hh`wCg��.zy J2[^�[����X&4
Z���x��:�q�U�C�Y�\o0�Z����M�כ��$s��g���>]\�T[܀��R�͙����<�}
\Q(������7�c�#��.W���������=��� �Tiz����]@&�'�g=�7;\p���,T�:�{���ݗ��,���iz|=�_������ �zG9{~��~��/~x�`9�j��(�0Px��#L��T�82��Q�M�`���{���l�>|H��b~�8D^��k?�G9oVGz��,���G-��
�k��F�F�����^��BV
��Z
�h(t+�	}-�g�F���4G����\(���
TP�H����K�Sv�W�7�8F,�C�K�>j;��E�ܓ������P�9����16jy����ɳ䪥nT(�ݝP��w�2��0Z��H% G�f���K��Q����%�V����Z�j�D�g��X)�Ɍ8�$��4���}&^��9J��`	'�8�T	oA:�`2��`Q�l�5�Q䡲��*����+�V�eњ
>P��g8x��x	�r]�Q��BH��x��=��S��{�+��6�S�Oz����fE�u6X0�r�5e�<`T��7�2��i]�A�/0��kNAy�*gm�(�z:�\�٭3��I�8�a��P���\4fh�u ��^����G��Xr'%7�S���K�78&G�������ʝ�C*`K������2q��;�(�GY�ɑ�#�A�jd�%�
�Aͺ�?K���8�� �`�p�
E�G���~�-JXF�Ń�T%���$:�Ee8�<���-�*=��Q�\-t�w��
��P� �#�$u�M��eM�S^�ZPP�U㴩�_�C~��A��w��DY��K֜�}�.��Tt�؎���-�Mh���ّzg�B�ైwé������u���G��E��+��l���ւ�(a�K@5!��:W� ɦA� >Y?�Gu��l	���2�d�@���
rJ���F&�a��{�;���G#v�':7^���̴48XC�m�7rt�_W�@�-���F�	�xxãd���?�o+��Ol��/�~ ����mo�2MSd�����U�&�#vR�'ѕ�۴��|���H�{9����?�#m���~Q��߷mf��Ȫ�p��K�r��+'N�k�@��aG����dW+���y_*�XʕG�?�;��zj���ن�g[�
��Y�4�c�d)�h�lK�&ʄ4tQ	�i,�����C��H�!�i��2l>M@C�3^�m�:�F>�|�NE.��g�	�§���r�JT���\��W���BU�%�y�q�,��f���x�ER�{�K��(��3A�vyu�d瀝�0��p����z�"��=�Dl<��A7��YG�XO��dRd`�9�˫z����N^��|t��'Y�PRYG ��sE�9C�0$9Y�$���L�ֶh6;TW���\;⬇>�;eXp�@)�����j:2�T���^Z��Ƕ���ib�=Z�W[i(ھ�s���W��|�:�y-�9}������zD[��u�R�d���h�=�P��hC$�Q�xE,Y�V[�q����3���J�k/�E2
Cr]���� K����#8`�[?�4�w-����WU�zn���v��� �Dy�S�����g�Q@MЦ`��P�sɴ&��g�P�#��=Ū�N"�i~�$����h�[%ġ�"�SU����oW*v�p�(8f/@����weNt��&���s��d�d�����_�A�����(H��i�+޼x�[#g��;�^�e� �k�g 6G�5ػ�nv�%��~���&�f��i�����e��Akߩ�#zN��,�����f0�
\�bq����y
��L;c���C�X�������u�=o�
��ǀj�3Dr ��Z��B�q�3m���:XԶ�*�%��@��z)o�m��Mр)Z}�h!����qZ��^ƜyH����|���T��I�������<W�Fך[7p�W��ynf���5�p��}�����b�V@�ݕQ��Z���Ϳ�3���3��(��b�n�EEPJ��!�_���W��z�_��� ���*��OЏ��/�p�g^�G�"`L��3#���;��e>(���Gr����u��ә�g���Y�f��DrO*�w𭡏�lE�)Y袤^M�k{s�$}����1��>��.�w�T���mDU��w��	B5�����m���b'�M=��an-$B�i�`I0�"UP��pE���ڃ�t �lo�cr��%X�TW�1�� u�������)�y�⸑3�s�>֋�^C�"_�'ZM��W幪�j��BϏu��|�P���.͸
@��*$�k�EC��K^�>Q��ꐊC��V�m����^�5��0ｽ�P�|Ihl�������p��'��o�N/��j�,�[���?���a��|���ܹ�9�����}�@9������X���n?S�̒�j
�/� �b6���]��������/���g���z���'kkk�_������+�_w �_?�������?��pe��^?ی�k"#�QrΘ��
�l;�L��|Jk��G��=Eo!+�έ0e���џ�������~_�FU؂)�5���G��s�P��W̑��y����	Y ��������O���u��os«��!�pst��
��쀦l�(L� �]
͈
��OE��>��&5c)�#�.�_��%�}I�Q"�]�;����L��٭��|\QX����{p�ٶ!
�}u̸������?Zrgx����ߑ�(�
�.$���l���(�%��@B��Q��e����TZ��kFűcD֤��i�8ܓ��7�֖�4�g�V~����T*��
�l��%�_�O����Ȝ�����=,���Eի.�]����޲�l=�m]�Ukh�_�]C�b���@I`V�z�l�p�{P'U�nl~@6��Y����2���Qj%R��$��۳9*�#Uc�+��`����\��@kY�6��d���p� /��>�j}�������Ab�-uք��x,�D{�w���"��0R�S�� Z*��ihmm�;���C	Io�|�*�ֳ���3�+���wg`��2��>ʟ�L��M`W I�M]���HR�V�8�,�y�ŀ��~��p/^�
OZvz�@|�|%���
��R|��K�z2��}�1Y���hXI�8�9��)/z� ��M۫�la)�g*��2���������X*p9�e�<������!#c匨i��1��J#�S��˫�l��`�����"��H�� �%� �����T�Y[�8g���-��G��`��ȫ��uˎ��kj�g!F��*[0�`�k�1��܍��Q���f_�g��h�2��7����C�Ne�[��.^��|ز�k@��k�"�yAm�>�rZ�D��D7Ϟ�zw/��^�c+M5��]%��q%����$�]��h&������\9����&�����8�g2��R�sȰ�+�:����Mje��u�<}������Ƙ�5��X��Q�):����g��C{s�Uxk�-H��f�$Z�3�|l����x�qg�M��2�4X0�%]݅����щ0�f!簣��:4�v+�o���v� ���.6��g2=&`m����9p62;��]=y����$�����֭q�P�at|��P�2ϫ�|}��isЉ4���>��t�cCe-�����0{�ɱ+؞�L�E�r��s���e5��q@5�/E�
ث������ d~usi����&a$��ނ�:���-g�q�������-�@/*�R��e�f%�=��hvڥl��I��0i]�k�v-�l�a��&�ߞס�^�,˿y���͹�<H������M�
P��=�f�W�	�q�J��f�Z��5䌾`6���mz��=�ҫ����U!��<D'3�m�X�[����lSJ�J)����W�����7Y+�P
t�p��(�w: n�暵�l+  (n��qem�~���<g��`-��sPl�Bl�*�Ϥ�1����
���Ӯ#��d�ny�;T�0^����f��GE���siѴ@�}�{�9^�|`,����D�,��{P��m c����4Ú����4ϲ�5�TK�E'��J��݉Ђ,�nU�S����]*`�����q���'胇w����F�W��a����"�w�|~��ⴓ ,�t\u#�&˃�ۃ7�3>��Q�:$|U��]� ���.���;t��'Yޒ�L��JL__�#��1��{�r���mH[���ώ���t�6�u
|�X*������3�'
8�u�bE�3〮������F>���A量�겡�P L1!���E��0}�d����4�E�K�:=B����M�J�~�j]8��!���I��q�EZq�[ p|����<���: �5y��Y�t�bf�CX_�Z^�iB��M2�v���Ҁ!N1���>F�?�o焮s+8cu��e�2=L�[��C�}���o��*h�j��a�|�GDO��@˳�z!�oؿ;�bcL���]b)K�V<�%�j�ס�W���}��z�v�W�r�K��D׽��ߐ��EO
���Xv�i;���sK�္ ڔ��5,-j]_��5fۓ�ㄼ���������"�F��A��[�%:�t���{��rXm�'`�T���Ǚ�����|�ǙW�_^���Ei��1���j�#5.�u�AW~l*�I�wRM&�� �6H��߼�q��ڽC���u\��AR��G�e���TQ���3Ku5$V�r�~�c�w�C��S�$˫��ُ�{�J��V�}ad~3��M7g�%�J�$�=ܽG�EnЛO������r @>]7���� aM/�=�K/�CI�Y�h-I�%Q�T�S��#|�	VH��g}�oi?=\~��_�������������_xy-� &�{!������z|}��� |F�>�hiw��>���l�SkG���c3�����ߡ��s=v�E%
r���`aa�H��.�Dv������7�6�o�gT��#�uX���  s��ё[Ժ��[��
b�$eO���#�5���ͳ����`-Whp��qG���=8�%2�)�o|�f[lC��Vw���<�GuȮ�oPMQ�=wa�ʓSrgI��"���g�A��Z�KK��N=
�xJ�G��<Y����T{C�+���`��Q/
�gujF�10�[�wn�yo��*S����>�F�)��P��zQ�}I����{v��3X�=��lŪ7���>��}�{�^�BO���� ��<=���D�uw%;2�2��^U�]��2��� ��J{�'h���5�{UN'��]in��@�w1��(�E�L��p�鳢EȜ�8���XcA��9.�߷�7Mݣ����
gU*����X��l;��;FT�64m�)NA�-u�lн齅����p�������@Vr��`Li�QOW�0v��?x5�f�5ȠP�o�ՇR��P� ��6g{�YP ���"q���k`���#vֵ�2�cI�?�<��'�ޚ�k��@��8�Ǖ�0��B8� ��N34�X��n��~w���8��s	�.�>3�3˜	��6�d!4��έ�']�+�l��ݦjiQr	p06�����c_+�ಠr��T亀�����Dl����
g��x{��j'�lc ("a�dL�w���U8DJ[���c��H���N	2��K���
�MMa9���Uw'�{u�`z�8:���A��1�~�lV<±!r���T��s� F)}�����e�;�4��o���-H���Vv��HA@/���(�+G�0��r��z�S���uδ� 8w<ֵ�:Y����pd�Ԙ��de��'	-)�n��y;ֈ��`��qD�
��Ԛ^�5Z��f��	d����Dj�F�b��I����	��N��˴*%�����t�f��<��(ф�tRZq=84�4&W���1ˊ/t��t1uʟQV\�i����m�����������B�s�F9��K0�+g!���^ܦ�>H�RoG�r{c對v��r�����b��m��B��'h���B�+ǚ1}�m2	\�w�l}V�^�E>��%� ߏ����z;��M�3�KϠ�F��M�ewU����Nu�P�̃�25G�h�&�üV|��y���Ï�pl�L�������ʙ�����F�%�y�g���˙��	us�U�6�����*6��M0Y�@�����4���w�k��.�b�+/�$i���h�ޝ��(�"���Uz���0ݏ��ji���W"�y�N�t�ȿ�cZ ���f��^�XyF[dN����O$�Q0�r�zl�-g��=�����v޳���t�H��"��z�D#M�6���g���y�;au�� �:;�(�M}�6�H ���������S���lz4�F�h4��'?����|�K9��S��*��ڱ�A_@��P�)�ls���Ѵ�+��t��s�H��U�ezRZ��t(��Z���fcc{��@N˚��'i�x��2��_��-��Y>N����1}�{�.(:��s�!����qn����3�E�v@ JB� �V~�.�|;�4��K5��9����ίl�r^��V���Z���O�4W'a/�^J0�Oe�&��8+-t�l
=	
�ڈҴT��1��y�z
��a�UϾ��r�-����ak�DKY�����ո�{U	Ci[��G�J ԧ^��a��.�ݢ��fUwRɄ�A��F����:�����Z�{A��`zN��L�?��X�ޟFAʢm4m���:ݞݥ�Q��k,���دW�k�<p`qV2��ҽ?��J�;���>?h��.@�*U BE��r���UB��Lp�&�]��Y�玤�L��e���з�П?�0��F�YĹ3��p_�+mi(c���F���W�8�<�~|}���C]Gɤϻ�/Ů*_�{�\��Ln�T;���/4�#X:�:�M���m���A�
��ڨ>���yU���[_n�A"��sz��%������6����`�� ����)GO>nl����~�#�x�?���ے����� ЀN�"E�!W4C����HI����9+��q��9��3��<%т@x�����t�}���ު��0�ȼMj̙�>u��~}_ݪ4�a�M���� �sz#ͬ�h���	��^xF���DJ���_^����A�Ǹ���M#��k"mR���l �Ǽ2��$���hM1��0�I(At�$2�yۅ˻��S'匉Uɶ���h-W�`�u%Q�?��2�:�[��Q첝����&�}יEj�+��'ٹ0����� 	�dn�b�5����"nXmǴ�i�1(�j�J��6��Cr��H@���}���`,� �E񂏯&8���P���B�+�����ȩt����od|�M�C��I��T�]'X��o��~�W���=0�_C���7�<���|���ȑ#��K�o@��P�U0bt.$�D�s�Z�4�ש�ͳ�5��E;_z5�~xm9���,˲d�l���t��W����,��u�:s��~��q ������r�B�+�����blGԩ�_T�@85�c����i���r�i�0Q-�p��WwD�	"t���2�����v����|��}:��Q����d��"���=�Zp�/�@j��?D?B�$w�TZ[}��(� ���Of��d�+C染��5��i�X�K�3pg"P��Ƚ~�d����.LU��2@)�z@n�6�L� �p.q	Em�k4s���35`m��K���k�P�?zQhk�FpnD��(d�T�-�'2���\w�"3�[3B����z0G�/�����y(�ө(�`[,]S�����@���g�x�L�ދM8����THk�;� s����Y<�z��Н[p6�g�4���Ʃ2��jo �d�X(�zl���#J�9=�tKTJS�S�kɨ%h��JlZ��I�=}V�Z�����S�-W5h5bB�Eq8C��2nF���`J���r��j��U�Z�Tц�UYG�p���a�V�� s��~9���Xz>S*%��=Ak �Q%�L���l�����"�A֞"x/�*��sD�N�.��y�<F��ˍ�N��`����lk���uK�zB�GPV��+/�s���Eɝ�	2�� �)�����} 3"�w�_chi5C����߫��-����n�׀	�ѵD:�Br�/�� zSG�� '����Q�Q�%z/��t�d�v�߅�F�a5�� `\�,�$2V�ȥx��
�C�2��cޖ[�$v��;�4��	���d�4�	���?��/<V8�|ݭ�^[��(�'G����^��@%Yz�.�e��.�p����" ���w��	ń*�a.9dTjf3@��O(I�o��e<�V�FM�?��9ő�\�L�� [Rr���P��"m�fc��_$掮P��&T���iу����[��&�4Ū8{�f�����YӡG�vH�tc<�uˉb��{ߺ��F�E+��:5�:v`�C.Z	�F�5�8�[���q�:������A����>eZ+�Y��ۚrV�����xu���?>���h�"��){E2VD�D^�gǡ��j?���f>��qy�ޔ��B�s��:�"�?g��_�)���������,���*B���Ӊ�����vB��S�-�y-=�K�3���.u���`
Pr�,t��j�84佫�9Kk4�	(�����1��]s(��k�j�:�'���@���:��[�X�p���#S>��Kt�pB���3�΃�d���C�r>A�i7�L�+]Ji�ĥ�]�kW���J����zk�8A����w�.)�@cS�æIZ-�Ҁ�2��Oo�3h�켯�qK��M��Mi�U��\Σ���L�	���4ھM����y�?��d7q\��+�p 5���P]]��B�+���
�k���6F�:�V׻��{ʳL�ʿ�h�F.��id�o���� 	�
Lb�
X i�l��!8��43����U	��]C[̀f:*G�������JABy�*7�`��[�цٚy���k�Q�����o�g�;�E��f�OuD�
,��T)u�����Ǥ��P2�/\��������R����$)�H"�u�}���4x�<p�:��,dA.�=N$��-� ��R��糣��
��y��� �D\šѳ3�|�la/�l`;��ϟ���'o�[���cP�iH�A[�ip���ː��-�T6Y�5�W�C!z����d��pۉ���e�DH��g/YY�WO�M�T�����E���y�3a���g�{׹���9ͤ	V�:J�"`Gi@ߩ���6&��%

�>5����x��ù�����^TWQ�Z�KyB�.����Z�.���(�z^��U�5�Bë�������l$�&?�,�3a@���K��d���ld�8h9G���@�U�~�k�i�,��;{�F��@#͂�Ւ�Ŕ&=�@���t��4�9�yd�ܳ�D�^��+aHl�!�,Kc�h9�f���we�Bd7+�� i��9�,K�V�)�t._�pK-g�rբ���׏�t��7�� ��h�d�`0�1*��KA���y�7��?�;ɬ�,6W��a0Co�6*P4�g���"� �L��e�����C
x����vT%���/:����tV�D�}c�uD�/�/����WUJ�\Z���+{5��y̘�?�]�R �4�:F��^ ��(om@�y����N��ӎ�}�]��oZ^���O���U#��bFE����g?��
�kޣq�wo����MY<��L�}Ϫw��7�Ϥ���Oe��y���dl�7���R]��JA���·4�h��ᅃUzb�)�'�p %�3�5ρ�O� ��{HRF��Kw�%�dF"��ҳ�����ߘ-β��zI����n[�UE�RD�'���
�z��qe����7������0�W�5�df��"�a����
�m\"����ӛ���o(g[�d|��ˠ ����FC0�іڼ��n1/��/h�"Y��YY�ߜgZ�5x��rS��;�F�viv>���� '.���,�{�ٚ����8$k6�|�C�i��}4b� ?��1�t(9���h��t�͎ҡ�|�ν�b�� #o�ή������U��
�V%]?���5��S��f�K�"��j��?Y&��:���EٳAeݺ���:��:��z���^�|A��Y��V��KM�F���die�J^�%�y#�Й��u�:s�k׏ ���y�6�5���0��:{?d�\X�!V�.x��nL�3+�%�E�aN��ZL���JB� �3�U��8���#�%��7��[�˪Y�X��^�c�rXl!�0�E���?.�B#��ظ�,��p�m�g� ��LA�׶S�)���gKu�����o���zV
ooh�3�~�;͈��<A6���A��iA(�E�Cꀆ�Q�@L��Oo��1��9��F�}dt�yiHJ��� F��}�k�~Y,�7Uq�D��KA md-�F�L��Ҕ�F5� �kH�9��<��y:Z�by�ʂh.ٿN �����kSae�ʺ"�����>k֘��El�0��nB�z4?'K+�	�#��}��\;ZN�T�V=�X!A��)pC�b(�]*�=��&�hYY8����0�R�-�
���>.8q(�S|��o�K��ܽ���T� N[��:���F�{]"���E^@0�J\���1������\�� 0Q��:����?�d
2 J��Zp{?2u���Y�Qn4��h�����[u�������,qz �w��PLdÈ��޽L��m}9�^�/�G�)����cПk<" ��l��v�e�
D��n2 _�G������
�o�׷'P�D�@Y��D>�T��މu.�
"��5�NR��A�7��b�Λבֿ��ϐ����$�K �b�##C/8RZ���T<�l]��	Uu��@C�<��C��,t� {(�	���m�0�d ,v/�M�� ��qBxV"����`g-r�q�N��
 @���;��9�u�,z�Y�S�=tN�X��V]uoQ������=2D�x���lTw x��j��3�R i�n������o������T�J�$K���q�����t���nU�G
,�H+Z�7�&j��r��WW�=������ .ݤ���eg������U�v���,#u�3����O��-kr���8�듺�CЬ-Ekt�O$FBf&緺~������$�.zoH;VIF̖T��آө�]��Km.���s]�v�3� ����3�8������D����=�{紆�w♍9��5� &��ܵ�B��)��*����V+�Y��Ll�I;�lHv��_�m�S-�ά�
��7�Cp�ۧ�ү4'��!Rڳ���:&�E�ug�����x9o�x���;�[���D��$-�B	�,�q��M��Q?�佶�S��NT+i�ܢF��,���-�,`��2��ҴQ� F�﹃8?oeiY�rM��ҩ�b��Kψ��O޻��k2�T��-Ύ;l���u�τ~��[pB�3@Z3(����$/AW���������u��k����5k���$��n6���j̑߈S��c[���s�r���܆i_d��
�ड़���~�|V9�gRJD��3��S��8����ܳ�Ou[�l�d�����p2��sZ�iey��l.�n�JX���jciΠI�R���D��.�+���t��-�@J��=K�4�j4C�1 ���{ �C�ó��m�й�k�͌��>��'��1ۇ�78������
�b�����n줡���U�l�tQ��n�0�X��+��&�9t^SeX��N�b��T���*�[S�H�|	�`Y�h����ʲ8��XU�j�2}��VV��_�A8�K������6�N�dy4�Ly��i|3 C��})Y`L�L&0Hpe�LC!���F7j��Z׃����f�v}o|#I�*XPVuE2��"9+s�G-����y����n�ɮM��G�˔���jfP�������.��3�^�:6|%�Q���lG��:�))I��5�wg��F�>S�.�*�C��J�.M�\���F�rM���+�M�yp���%�!��kk7���U�F+IX5�52���9�k��N�$8����O,��&Dv3oHQ�¥��w�jO��@/�3P�45>i�GT/��B+���,MF��.��sPE�ͭO���+﴿��G��W�����KK�^�fj��P�E�Q+L� ��WUځ>�
�ߙn%��S���L��II���Hf�'��c'k�d��w����s�a�����V��2�+���Q�-���w���K�BB U����c�`���%���T�$M2�G��&L�=��i�ZQ>�^��`�
����b�y�T�i��L�T:�3s��^z:�=f���h����op����~��$�z�� �D�d<����⣞��	���M��k���*$�Dk���-�ڳ�Պ����`���;�G���oZ�FA�f�T�~����K׷S�3�Y��6z��g�����fTڰb퐀�#�j�OX�e���l��Y_@�*���� 9晴���Q����/�%.gG{N7A�\g�3יk��q �Yg�5G������oc��ÛotM�/g�?�]�q����*����O?D��P�E��pd0�X�*�Lq1gn�gYx��;����;M3YK}���ٙ�f��Ư6F 0�ƕV����b�S2�.ij��^��y5�~S'�O1�o���`�P�HG�Q�Y��Z��y��e�1l ��˪��	��:�F�P
B9�����iJ�Dvo=�y����z/�[ ��V�H�Tdߠ_ul�ˌ�`�G?q��f�@�k�`h"����-�<�@X�������_����Ř�s��`}=�/`[A�@aT%Hu1Sl���=ѳ���#xB���j�ս�L��#d�M�ڮ�C��\���U?A:�\h�TO�q�x�jC�6�3b�`�[f�K�.8����8�|)~�c���x��;�� -������h����T�?�T5x�R)��s�x;�|��G�\�?��:�����y[��;}�	{����^}���x���ѳ����ܖ@wjD##�����R���Ś���bVW�
<ĕ�B_5�-���2��r� p�@�
���Mh\[񛊟xP���o1�~<�=#_�m�k�[�CrT��d��W���y����(*c7̩*{���zՍ�0?'Z
a/<;�~�>�.�� �&{g�>І-%2lb�[xW�� �a���|�A������А� ̒mP� �Q^^x�����k�j:��s��^��,,؞5I3�Pl�Sr
�|uK˖Tڂ`l�e�|̘�@5��L7�C�G�Z���ڸ�rCZwޓ��<;&�?�4"2%��z�<�xF!Պ~�]I��J@1U�r�ı����������ʃ��	x�n,д�z���b��W[Uk�\�j|��"������1�Λ���B��!�1�),좟^�@�r�L�s��k��'J@��޼�m���soէP�C�d-f����`G�+o$���8?������l+�P颕`�x0�R����Ī
��E�%8��9�E�t��ܹd����ϊ:'��&p�0�W֨�R�^�S%�u=�p	�i
�L�M�4Od FiE�Ʋl�dW��0��F�l�����ʧ4P�Œ|�#���	 �1��qXI��d��J���$L�8��X!ˡ=�	����q�����j�����^Zt汴#�tV�L2vVɀ����a2o�,\St;�f��8�7cBi�O��NW��3�ͪ�s�H��x��s�m|�Z5��`��P�kƽ�� ��mF�ws��kT�4jC��jQ����oY�P�e�f0}oN��K�$�O�ge��J�J'��ʊ���Z�Lè�A�et�>�i�6i/i��Fi�1�^ɪ��47�p��.jO�r�Py�GL��'�F�s����e!��J��
Ќ�F ����J/)��͙�z&*p�d󊅞F˦�1X�% L�*FG��ZZ���c\�Y�u�_C�q�1����;�!l8ú�~�X-�l�WB��h�S�Y��	�%��2ǾW]���Z�W�L7,K�z�R���yj���P�MEkZ�E�͊���vA|(3K���E�)����!d�I�)NB��)a�!�&����0��oT�i	z�2�`nM) ,W�F5���M��-��8?w�lC��AV��\�F��4�q��=��g�4pj��U>����y�X��Q�ζ�I��(i2E��<6�&gQ�ȥ�@���Yޓ���ZZ�/�HП�<:�H?�s;̟��{�!#U�V�peς��K��p�K$T>U��i�r�dTK��Nu�p �e%m`S2�qV�%�4F��,,[��<$`Al_c�8c��ѫ��!�f���fIZ:>
_D�u��:�l��1R��[{���x�bg��J��)ǧ7:����wV��f�-d �IV"��oM| }��=l�6��&�0�/��+����k�M�|��74��|E�e��^K{�h��A�|g�X���J���^��|`��E�,E�aKe4o/@ +�)ڌ�oeę9�u���S��!v��U�Z���q����Nغ�Wћ��S��c�k��&�L��*%TQ%M��%�I�����*tif�Q��p�L�^�W����
W���z8��$zJʕV�r�2�2��B�F�5Z�Aڍ���P@��M;QV�i���=^����ᦧ��J�H ��y�F2$t�ki��K?��K��eU	z��Mz����V�n-�f;��G���wl-��T��*My2p��{���I��	���e��@р���p]�mN�WZ��s����@������
(|���)�n(�G[@��d���#���7+uEآh�����-,V �J96��'_����>�S�X�)-Z���+���Z�]�~��4� >��Y����[�o6�T��>���9
`Q�͐�&)�F��d~�z�C3^���y�����4�es�<��d��~��?ٯ�.M��� ���\g�3���c� ��t{v����_�����}���{{7Fq��h�dA��A�&�>Y tY:�r�0m�9����Lp�R\�,s�9m_!U��S����ۮ�_�������v�%�f��"�EE���_�xA֕�DGZ�Oik�8]��o��p� ����HJ�A�2�Jg�l}���e�b#�/z��\�,��y���� �����F�I�nM	�&<FEqѨBѪR����18pG��ݲ<̈p'��%�e�5Hj�����P@=x
��iۃ�d�x�+|�(3���FJve	��+�у)�Nwr���3H��7/��N��LA˗�5��G�9a�8q܍c�u��(�U8߃+%z��ʒ5�ج߅�P�� #���Y&sD�����b]g$�I�Wz��ġ�U��:"m��Z`�̈��3�&I� �Rֽ���8���W��e�������tF9M�ĸ�*J�	�T=Ã(m�L��e��<�Y�,P��ր����Vk������j��z�� ����7V{j.YB����G���t�F�Ѯ�?:�
x����c�'Su�`����q)K�hl*e:���|�-�s���O���'����A��U�Qq�HYYz������b0~�҄�1���_-�C ��L������l}����|����{�Z?��88B�Mt��j��_H�����Q��7/-<�䟵���n�<�OH p�{,��1��u>���\g�h씵��P�:������
�Z���5�� 3SYԢ�y���	�y�Q��R&�p9vmC[o�p�Y9xQ��|�Q�Zּ�f���������ABW@��Q����p0��ȠjO]BD�f0��-t8*�������oX�H%C�N��Z���aQθ8g�K��d������PB3i�f옓��cz��#t��	ꦑ��]�/<�v�^2�n�x�j�c��ǆ3�`��-d��˩�*�
�F>Bи�K���AV�� ���	��T�/���<�C���2�l@��6N��eS�����3�>d�L��"�%��0D����qΞ=4:z���e~��^��3�|o1s�;v%��'R�U����e�w6 �|��>�c:v�$���k���E��	�w�~z�ϕ�bL;���	^�\y0Y"|��U��Q3��-y��"Wߵ����9��p8�F�6�������j���vfc��q���#�����|6�]����ϥ]�Wi{�A�Q/9���@2<���I`U�����[f�����Xm??�%���:  �L-��wQ�*T4>c���K��8P��=�)�:��N^��_;DǏ���{2]]p�9�/��|�N�~[�ȍ�ݵ@�ȑǟ���>��;-]��h� ��ڙ%��������f��kV,�N�MG-k�<Z l.b�ǳL^;���!��]p�9���D�.ϭ��x�'n��e�,�h�e~��lKs�fv�r���$���Xx��n��KÉ�E��Q�G�G�b M*���	5����ky�^z��XߐLԷ���|�Χ�=����}� ���k8Х��Q�Pc��`A��]�M/�:&�?T�PqX�е	�m��s��%��&�fè.�W���g;�ZZ[� ܖ�Lhk�i��O��~�9{i����f]�	�q4�n��0�s�`g��8pȥ����U�b~*��Y y&���˙G�W��!�i��Fh�����ޙ2a�1���ݠmβ�gl��g��=��!���	ZZ��� �TM8�"�'�M����L��'�oBü�+I�Nk:���A�KI�d��cB����VEF����Y�s&y��+8G��+�J����'Ā:�Z��nF)h��! 5
�pK��f�0�M��D����d:#Z=�Eu@H�6?��{%���P�L�̓O@�!�zϑQ�y@^nz#�SG�G#ڻo%���y9���P�=( ��E�к��+��(�/��.4�i�ύ���v����AT@�3�.�ߑ��N�ݣ�\�э�9����.�G�ƻ���u:q�$�����2�}�~d��[�}��7�Ok�i��p�G9{}4Ш�"�]�E�c������ڪ3gWomT�Z����<���7���%��ɲ���K�J��4����p,��͍m�ѳ��G��V��l﬋L�  �K�n��c���6.S�2иrJ����i��4p. 2&�Mv2 ��%��ܷ�j��|��DC���3������vM��~��=&Aⵕ]t�Y�2}��|��U�e�h`�'�$�X/te Sr�R�o�[ƺ�TGP�].E̦Tx��̯Y���;�Z��k�>
++ת_��R�a�Yǘ8NoxY��={v�E��VW'Y.ni�n��F�8�'�!�M�������a-M��\	�3�ok�P'5�:��5۽��v��%C2���ʳ����"G'�5:���W^~���whii��t���g�Z^���R��g80���eR�����b��d[C{�K���>Sw����6s�K�[���z�����~��(�Aѳ%x��`��ŦJI��Y֫^<~�.=�BZ�d�V�dv�5�ԶKfK����Dm���i��1=����9�.��RY���F-�)�}�?z��Cϕ��zQ?���I���+h�s"�9/R�����p��<�6�t�X^�c���lI�7pIQy�!c�1@��C���a��ş������m�İA�*��3י��u�Z�~�  f@���V�V��#���_[���~�i��m�.�Z��г�P)�>�L��ݯm��ݓݙ!v4���r.��{��_�
f�(g���/>�h8�ӥ���Z���d�\�,��U~*Z���5���CL	�?6����8F�r�?�d<���67$�W�^:��;UM�4$�C���dH�B߷��Ƣ\[�,A�5��V�nCP���8�1��a����f�TNRLp��
��d�q"�Q�6��p_�
��wd��z!2��yaH���Zƍ�
�X�wWm���9�	��k�������3��K��F��C ܁�����܁!����(@���ma�삡�KPA���#��Yf��3�=���q���6�G�`J�o?��6E��/�#sv��rer�g�&�δ��K0�b����0G�j������:3�* aш*)L/�s�T�Jq\�e����L�H�A/8���T�7i���O�ecR�5�?�V�x	x�X8m�wf��;M��✊A,��>xf�i{�[�%��.�|���q%��u���;�PhG�k%!i1���Q�謝A)X�ٯ'g�+�ל�P���,F�k�Ui���n�60�,í�� O�n��J~�tM$�s	$;�>V�l#s�3��"$.�NC��A	GK1���G�95��gZ�\ּt��<��B6kS*\��1��xz��ک�Q� G7��(�g�#3�Y��F85|A�U�-Q��~/�����Z	��+�|��.{�`�s�����՚��/�Mk��(�����&�c��
;�m%�A�ʋ�\u�b�[�;hV���O�S8T8���j�ʢ��~QQ�Je�y�J hYd5��J��V������̦³&R���@[J=ھYz�V�	D�MWK��u�=��/�tg��l��yF���-��e��M�����h2�lu?U�:J���ː3��$dU�ਲ`��J�6lY���ه�t�V��2դ\ ���E�ޚE)=����;�|��7gRf\b8liiyB�}������lwt�m�8���A����N�^���V��gS�P�HH2 ��p~|O+}�U���d8Y��>�,*Swo����׬�l�s�#��O�������5Ư���9g�������o��ͣ4��h4l�u�6Z�L�M9K��8t}�I�u_��[�[H��3v$�g H+�z�KF�<�٧��� �'ǫf��{σ���O��Ǝ�N�1�_[[�w��b���>�m�M��3Z��(ٟIKKVtS;���mT^��ɀ��'aQO�>(�P��I���x��r�&���Y�E|�x�9;���W��n���9��I����׳�4�w\z!}�K�B�٩L�3��J��@N�Y���E;-2:����(����w�\���	�up���<��Կ��x�t����cO<K���:�ră��A*�������� ݶ��i<V�>hJVl���(�pU�����'+�l�d�0q�;��Ǚ�i
B�3����Eni��^��#��"�����^z�f��hK�[�Q~�Yg������r;�����$�� �r=Ug,�wL��d 芊�� 3y�.-�+���6���o�����J>w����?J��W,
��05�w�
}�����=�~�-/3 ��[�:��P��� З�����T1�Tt�Z�Y5h���A�ՙ��,�T���m���z�����L��+�e4��}k��_�z��/����gj���䏬3�W��|W�r$E�H�p��u?�Wz�*��eBh�a���r�����u�#W�ҁ�_���z�fy���'i+Ù�\2��;�q����o�w��'�pm�L�Hb�<��B��d�5)�c朸��	*{�koCh�]�`���`��O��z~%�4l�1oީ���7,��>Aw�� �<�#��|[��p4���^������{G�y'�;�ʟ��OH��@�����,]�inK�ʊ +" �>ה�8��!�{��a�N�(�z��KS��Ό���uߙ�n��?@;;s���k®���%z׻/��}�S� ���â�d�ћT+뭌:A���Q�"��^����G�{�1Yn4&�23�S�T�V�g�vM�����w?i�,��[�K���r�
NR?W~]۵L��OЧ?�q:q� ��^�$g�Sט.��a��,;�_G �,y\�8�a;�o��Ӧ�vK«�ǆ�ʼ̍�B'�N����e�M7�HϿp���s��'_x�^_t}�����ik�I�6�UbDE�Z$f�~˴m��S
p<��ta�I���V�wd~�����0��q@����D�̼!�c:|x�n����*���G��5������s��t�֩��6ub_�P�_���y��`,4[�U�D{�b8�Dr���� ��D�V�@ q��YFLg���Ǟ�i�k�J�`�������f]�t��{i}�H���=�����B}&��E���в&y�:T
i�W�02���Q�th�B�%Y��Z��mH^a 6H����lo)��m~��Љ<��N�w��S^HU[4r/��-E"t(݋�K�絻��k��{i׾�	����+������oѷp��ov�n��_�xH�ԋ=g�̷�K��?�G��y�Z�ח�\���  ��������,�ZO-u�\p�ֈ�Sæ99�L6���3י��u��/\?�
 r�������ӥ��v��Y&(�)x��~�:��N���x����=R��{}��{
NR7��ᢂ�2v%���*��fY(_FK�t�[~�ML�`�L�P,�V�.Q<�F��CV֔Q�]7���q��+�t�x~�4��,X�0gΫ[�Jd%�^��Uv�u��{�5���sϵh�@�I�&?t	N�*8��΃̞�^�>�o��@�3ߐxn\�Kl? @#��wӜ�a!��9GО�>� ��"�."��ں��?�C��HA�4V^�{1���>��+UCz�"��6��a0Fl�2j�X��ƚ�R�4����>�`�9R�@����Ld��y��Ɨ�r�S�+3.�"?ÃT��s���J�nM���c��U�<������ǂں���hX;*�	�p��Ye�R���l\�Pݻ��؋CmсUt�cD��){aʰgy`(^8bQ�t�JP�������q��a��r�� ~�>˫#�zά�t^�^sb���k�% ��"5��;���}(�BV|�!)M��zb� ?:���9��9����=�C9�dk�d�:��?������<޳�ʞ������/MX��mE9���k���n��7h�AN����
��tN����̠��ɖd,�~cu�
�E��J�p^�<����Hd�V��dY?�G&~�n�������KŀT�σ<5��BW �ƃ��T���������V�C� �0�TT��
���
<�A3b�'�w�$�Ĭ�{ ՁӬ�^3P)@�a:�g�����+�kx|��6Wq���^���ѱ� ��kLEnuÕҲ�.��c�*
��_��Q��j0�?���|�u�Ȳ 9��W�dRyV��1zK+�D�=���_<v�w�vf��%��G�����[ ���e��:q�?����O��w��>�	��:!A�!��s#`��t!�>��&���Ix����;=c��;ʺZ��u�
���|��;��hg>��d*e};����E�<��lu@앶������Mg�t�ݏ�#�=C�}�c����%wK��sc7�w\��� $��d4R��J��BY��8�:)]@��k��1W�@�9^Xl _j��,�4g@r���׏ѵ��F�����%㴃����W^=I�����KΣ���w��iuޠ���'ZZ��5����4�Z�������#�S��ϭ�Rց\_��66�l�H����z���λ��S���7���E��'�-z���陧_�O~���O�������C/�%�`�Zٰ����fPl����,S�<�:�Sjs~���}����]*w��1�5�������\G�>�*W��1H9�H��3��y�Ez���H_��e0��9J+�W�ъ0E/$�O8 "xT��
B3�G��n���m<�1ܳM<@5�d���8��wf���cz饣t͵����;4�O��z�~���t�z��W�g��>���g>�Ӵ�}�F�Ҳz3��n>�����\���Jl��;�L�WC�)|y���@f��hl�4�7��3T�%	�q;�y���n��~���Gi6�%3���"������ks����_��?����?G'��k��{��j=��$x��}���0V��/H�	�5���p�~̽�+e\t0ӵ�f�l�F��nD/�z�n����WN�ܕ�F`�lrgӎ�����[�_���h4ɳ��<hi���;��\ ���-S{�K��I���xN�U��G�7h�A�Xdtg����L��D=�t󽙯L�4�f�* B[�Y����������L�רBof$N��y�8�]�.���4�ׂ�u���6A���?�dV�;���HA{&��z�mI`1��Nt۵7���r@" �<�ic�=*�@��'<@O��}�c?E��ډsi��o��j�G��x<�0/�b�/�S��R�7S�M���s�n(%εѢ��x���3ӈ����2m�����[l��K;�@��t���]Ow�� }�K�J�	�g�����{�Kit|�;�o���E}�ևa�8��^=�(��g6��RY7�1w�D�m�?����hg'���D'f},���٦��&=��������G>�^��/��ۇdLR� �WNkQ^�l�H&���!�	UA*{�[����-$�w�
���* Kr;�VA�,b0�4�߹���`�&_zS���j��3�3��7�C=����~�����
F�'��9���K�7T��dm�g�-�T��m.�qЈ�Q�{Ͷg},��
��|S  �=��|�9��{hg;�g3�� |XA�4�e��/f:�����}�c�k���f֥��[���Ln���bP��:�Op���$���Ȃ����
�HT��>� �$�?����u��FO>�|֗Uw��:}G�o'�>���ӳ/�g�Կ�Yz�{�A۳�<nD�r?����M�ym0�'M�̿"At��SE��Ԛ,x�Ϛ4�� �`4<����1��>詧^���|?;��m�:��������˯|�.��b��>I�Ia�-��"�gH��T@cKd5x��~t�%��U&�'?�6���g�'����� V�lX�/�98p��<�Ε��4�䳇����K���ޙ:�m"9�F_Z�RuY�3��F>SC����/}���o�9�xX� �܌�����r�l�?�g�y�������#/e�-�.Y%�Πi
��u��F�!�v�y�2{��;�
�n��ᘃ�w �m�U7`s�蒷de���b��g�3י���#�  ��Y�M�~���C�G�ͥm�"�ٰS��1�L֘�"�^Cǳ!��ɣ�ge�N|�)r��.�Q���f��?.x�-�B���p�{>��5
O�f	���D�;�E���͸5e)v\&n&�kN�x����p�����;��vLI�r�&D�������E�Ί� Ӄ4�FO��0�2�T�ȱ��B�� �G�p	��{D$W���"��/�J%�1�1"'��fj;I�7�N���wS1��F>"-cT�}�\+�hS���D>W({kFh��C�����
$$[��"QqR�+�`=N�dUJ M�N�)p.��J�^y�<
���T�{��L�Vt�H����L�-��>��%��}D&�8XK@*d����c� ��zC<Wh�X�]�M9�c
(��w�9�@s%��o�b���ġ B!�]�5xP��Xh�vx�-%P���>F��Q���E9Fp��r}&�i�=��sXm�e6��ޓ�gϪO%���N�,/�
������$Ī����k}:���������`�}'�~0�;9�j!�GrP�����3��>�Ev �}�^�/Hp�%�N����j���ϩρ�{�2�/����>T�Ig T�+�D��`)��>���OKY:e٥e�|f����n�u��`7$��N�t�x��<��G(�)�Wo�Y��'h6OS���y#���Hp��KV��T����p2.��6`���Tp
 ���͑�WmB���L43Zc���������
�����M��GdG4ڲ��sA[�8�*f�68��p��
�F*__�%
M�*j�N��k�Z����G��B�J]�'�C�9 ��ϥE��W��AT΂�WL�4ɦD#,�]���:�ԉ�;��c.���c���k��'P7�5��w���{��K��D;}C����q�(]���3M�M�ٹ�y�}�qi����M�q���)� �X��9́���s�7�V�����8r����z�І��I��فЈ���s02�Z�6�7�q8�~���>B�n�|��F�	��Z��^mOa��Q&40�1(�P��& �Ъ�z���A+s��9���ƚu=�ȳtӍ����W�<��^���C��c�_�v���^8H��������o�xp%X��uP���Z�[y���\^`/�J���k2����B"�IM��3	��o�t�u7�3O���1.3́�N�`�RE4�����}�[7ҩ�-��y7��N�aN���fTt)އA�����W�)��-��d`T�	u���&?*<��<*�i&R��������mnv٦dOzc�x;uv'�Z gj;��i��տ��.�Տ�{�Q��NA�T��M�	��h�[���$���џ"W�@%���P=(�!ZU�}��������ڋ�X�KH�i�UXN�}#�[o��^}�E���?Oӝ)M��e��5&�U/�.	�Y*-�"lѰ0|��Q��A��/Ӕ��L����*��|�L��O�d�y���	���?�[j������6��$|����z��-��7���Q_ L'��t���d����z��hD��FA�}�Ir�	MR@K��[R��{Wwy�=�2]����y�s�$��FT~��t\%��R���/���_��t�����0Tc$y��0v��3��uE�Dh�u��dJ�r�ϙ�-���=ˮ�d������H�=�B�[�I���V�������♧^���������h)��@h&���'{�J%.�˽��\u=m��,�rN�M���W�f�r�����	�Тo")�s���������|�&|Ԁ*�|T�R�@k:I�"���6�w�]4��i������d�Z��f���$��{ �&��$�|:� �M�Jf�$��>��eA-�l�ww�W�G�	�t�=���
���$�g�wRҟ��'e�� Jf�+/���������D��M���#:����dz�����R%�ė����)�O��`A��7�u'M�1eK��蛁���ι�}���5��3�p��{54V,�Mƪ����H���H�'������ܚ|&G����r��1\�)�(�� �;`�i��E��&XRz�FHo����3�Ҙg�+2/�+�+���ݐ0hE[D����赙&��9�A��M_��g���8��Yd~�j�Q|��Ǚ�9�WT�vm��k	Wx������W�����4�L�)�S��T/dٶ�����7�F?x�0M���y��@��κ�������� =�«t���c��9�V4"j�Ugb�lt|��~jի���mW�?��J�G
$6�)�=�LN
@���y;�M��֕yﶥ���Y��I[S���gH�W.���u�o�{t��:}��+��]�@z�����|a�M��1E��m���/��`��j�\�b���,|9w3b���=Dw����T�G����&�u�d������������_޽4�v��F����^�&<3`�
�O)U>�|й1����k�;��ɒ���*���(6�ۍ���s���v�coл����CXW�w)s�EDB�U�hT6�(�<=)���o����'��7]���(˙�ĕ�MmU�2�s�@9����T�:�w�m��l��w�L>��oS�1k�Z���|�s�(���Bj���������K����
Љ N���+��&�~k�5���R���u�:s����׏ �4}/�ml���u�m��k}0�7m��8�,�@Mp#�;���9/�:�ȱs��E������ɘ���+s���)+��Q��ڴ�u*��?K�	A��X�1rd�U�PU*�QJ�dfA���fm~ߋ/>N��s+�wN!��f��6�`s(� �_ZH�8j��#h3�N��2�d%%��z���:�0��ߜ!u��`hN8����A��1'�iJ?ޑ* EEX�&�@9nP#�~�
}��Y_#ũR��;��P�U�(�g�)�d�aΡz���Os,����|��=���ϥ2C��,��T�& 5�xEsv��'MKp�����-���/����U�P�k�j����`�~�������b(_���8�uW=���S��b(��T��E߀/��K3��+�s1+�	�hqn�e
VŢ�+-"#�̯:y�l�����}!x�)y��GY���@�Ӿ�۞�y��tK�݃g�j|�@6x���Wu}�-�aӢ=���)P;�*����iU4�sڃ�\���|P�Yc�T� 蠮�P6�p��[����>�E0 Jm`�?F����4 ��=!۟t�̉�XF^�5���Q�m	|�e����j�K��r>U�_T�������Rѻ/��0�@��;=�L�࿍�?���A��k*�%��v�OcEv������}����ѫj�{D��P�F���yD���[)i�:MԂ�3hl���`w �i���M���s��GiMЖ�*�5L�n����U <(n�h�A�1E;����3������ߘ�0 'U���
����I�A�0�V˩�d�De@��R�d��AV��.�7!�V�{q���W�|�>1�E��8L���*N�2׶m�W�)o_��T���()%�$:&�z	t�u��㏿,�J��c����)j�o{'��ij%�1d��bK�=�:�ǿ�;������y`Z�QR9�7� �8�C,��I)�|mb2��@�QV��1;-�Pm;������톾��k���M�K�nRg%�&"�"�/������K@��;n}���=�>���4�`��!ߓ�C� К\�&w@4pb������y@����O��y����H���e�w�]��ى�e�[�h�ǅ���;M�HpOxr����7��苴{m(�		4��U�6|vFKVL�*gé��Ơ���L��' ���'u|20��W�{��S��|�mGv��翇vT�%�ͨ��}n�#����hyeDx����g����3�d�`��Q�Кm��϶�j���ޚ�1X"����Y V��8���p��&��W������J���F)J����!�����A<\}��i��/Ѕg�����ir��4�=�}LoQޏ e��R�)��z�s�\J ��������n}�fӼ�S�M޿�OW��y�n�Die���/�x����?��ߕ��vhaO�Ƥ4p�	S�YOr����݂���Q�׶�[��bߔ
�dbe��+70�p����:|d�v8��^��5�1�#(����c�8�k���}������L�;�����'��a�5	ϵGfn����殻Ȟ��haCЈIe��!*r�*m�{�e�����|���� ��8H�7S
��eNI�?ƽh�o~�Z�_��ߢ���)�Z�Y�}t�KE��	(��H]���#�0y+���5y�ZfY���	��� �,��9q�򫮾��x�e����"�V>G"��q�~���Y���m:���o��
��?��<�-!ʁ�/7$��2�s�k��X6��A0BG��E�A�����c ��hW׍��p# �vsFO��(-�2-Ι���D�T���kʙ�'�'.y/�-��[�7���s���3�'�E|j�f�E?C9r�
��2��l١�?��W!.���cg�7�Z���;�{��q�͈���o�j�o��c��$�h0�/������whue(@AiA�Zi�	�O��ƴ��1�ekA��i�!<�.ī~o��;�@h��m�R����U��6lbW'c�ik��Ws��V��}V֞}�E��;铟��<�m�xE%���&�y�F��t���ً��N5�ɿ�C�;��γ$ �d1�����,��ۖ���|��,���W�4vMV�U=˔��ͼK��������s������ڦ��}�6��󼅗[E%�Y �����[�Y�����nm��l���,�.���m��K>��Z��ސA@"��U4S��I`�)*�ô�R�u��^~���ﯤ?��_��k���K��E7��&ʞ@(p� ��(Aa�JF����#��Ѫ@Ik�������_�*�=�r�48ΕM"	�m$���}4��4=�[-����i�1���R_\�v�&��=��T�"�{_�(��ۯ�kP�A� Ӷ����V%�mй���x�n���,��D�`3蕟�Ϟ,nF�WT�����d����+�w��+
�TQ@-Mc��,��
�zr���_k��WUQݎ/؀���U�^[��z����W�'�����}���v&�'�x��~��Y�( )���'���c�"��B�)���y�i�q{�;n����������=�F��q�'&*1��^TO���g��&�20gJǏ��6N��絭�3eޤ�"3��Fr�Zy�p�iY��sz��!�b���J!f�}��O��my��n��֕K�x�j�ǥ������ZqX���\g�3׏��-* ��~s����K_�9��S���Y�b��uf�\��R>�H�AvY���=��k�����,��b)����G�A��g���;�4�L�3Oݗ���O�rڵ{w�_�$���Ⳑ�a���������iG�[�t�}����=��m 6����:"JҼE��*�I����N���_��%6G�<`��Q�W��m����k�?�s�2�"��`���<Kϑ���3�	��"��J5�*��	�"�`�)hp�7��TE�4�2����)%4���0���ms�ù|�Y��j��v�<����FC�@W�˯2�Q��~j�^q ٴ��|� ���� C3��>XK9�ѝx�c����m!-Q(�}r�)����ĔjͶ���IX�Ps�f*,8|�={h���t3_y����e�%����wm��1X ͟��SKֹ-��@�E1+���	}	���	ٹ����`'�yWp���� ����BS-N�C�,j͔-y=�%CԖM��z�s�2�� �d����A�8S��m֤�gS�x-����L��K���c�����S6k댟{��iU�h9c�hc�\ ����i{�}� B�# ���uJ<֨�i}�xUk�6�� �B�5�<�����)4�m*	�D��^�T���J�o�<Yf���%��Ԓ߇��vɰ0�JJe"U|���t$��Tm��dw�������.�r&d=�o+/���+ܶ�c��%^;�B�!��u|�o����K?����mJ�P��p~�9o����g?w��~�{=J�U 	�ձ T ��@4��E
��)��h�d7�F(��:k��q�Jg� �G���g��:ɸ���|�p�H�w{�[���Ӛ���d��O(�G ��?�B0.F�1����h�q�4�b�!ۯrV$����&��C�\�cL�Iz����<K�ygސ�͙Lg���%���h=*PI�]���|H�������'���ୀ"?O�tE��I�sYĶ$9�*;X`=��EO���f�!Ӌu��֬7�y������+hc}�:N�cgZ%H0�Ϛ�,��^J ��� ;s�wM��lCW}�f:����M(ӫ�d�~�r!H@�u~C~C*Ϩu9%D�7�X�Jkk+�u�ܑ�9�y��� ˆq�u�8�l�C���f&oq L�y���́�9}���ї�׈�r�h%�ށ28֡�C�zN(N����(��>�U2�V3,�����2[��ڛ�gj%�y��h��[�k��=wx�8�?o�N�=g�w�X�"��Mo�}�2�N�錁趢�$���>m.u;0�H�S�x� 2]�P��H�c.��߹F�;O3�q��42�_Y��s@.i��`�\�w���y���7�z���i6�=F�}��)�5 ]2>�@ם\=��A�UL��Ū\�*!*kt�8�x���N��W�)��@X��q6�$ ��4ū��Q�:p
�t��)�ۿ�g��Ch�3>a��~�:�� �)�"Y�<�ܥL��iH�SU��[�h ���b��C�2����Ut��)i���&��y�ۜV�7�x��.he,^�Y�\���2�\����^������ޕ�϶�4s�ʬ���]�\X�{����`����%ߑ�^�ЅY?�R��ܓ�]u�m4��4�{6���33ɻ6	�1Γ��,��V>�;��ԘY�׿~-���vyϖ� �b�?��xX��O��U|��l8C��j8�KX�8�[nS�zQ���,�^ e꺏{�9)Cκgz�?��/�!�#�H�O��KQ�r;S)˃�vCǏ����o����e�tJ�70�.M�L��a�v=�����F ���Q�:�b�O,�6d�� �3�,嗟�ƙ���������[�9尃gK���f�������_�t�7�m���l�
`z��ZC���V�[�65؏�j�X�,i ^��� @�8Ӂ����Ǥ���F��GQ�ݤ	B�������m���y��LmO�������O� �b[�y�J����J�i�����kA|�W�Z���x�5@'�֘�*r`�h���~�^|�ڙj`u����:�uZ�uo(�1��Ɣ�b��{���=����;���O�=?{K�$�kVs�^7.S�g��y3T/�o�ךJ�Y8��>-���`���n��wNg�bcB����t�Ⱥ�c����d�7Aԕ�8cޞ?��k�@��-��!}�[����o�d$4�]�kI��R.�y5�� ��oc�E��
NHS29�3nCc��F��%��O<Kw1mf��f}޷>�krR]3X��1o���mU�����_��韮�����1��I���_��sp�m m3ݗR�W��(ak$�TI ��J{7��V�<�u���<૿{;�:9��dۀ���e�8�o g<�J�,?j��y�~c\s��t���A�qS�p��N�w[ 	$�i��S��	I����5"/��q�oS��1 �؉��+�'����s�{7
Z)�~�vR�#����i�N�w�-��?��,����3��Ly�h�)��*`"�hi�}�R��N��N'�)��TX������k0��-�������c���ᱬ�=�����s�$��`ѥޫF������^]K������8��w���}�'��v��E���)x�����결C\�¾�{�6�,�������%?g3/���i�"!�C��H�$���K�%�G�<ק;tpg�f���us���:��Eq�ۚ�ڰ^6�>���w�޳�[��������3י��u��W�7 �����>��уϜ?NϏ}���v�k�7� 8�$h�b`0]O��;q��~ޛ���?�G��T@����9oC'�STHE�W̧�̬���-��߿����}��Bێ;y\m�^��Vʪ �ݑ��ќ��=�����ۮ�
';�����-l� ������
��
2�K��4�ߪ������-�hX�γ"gY��u��Don�d��n�R�<����%`��]��2�-s��ќu���!!N0�̸�M/�e��H(����T��'�]ٻ�� 	-��=�͙ KЗ�
�H��p!��؃�ќ��` HB�0��Ѓ9�Z�^�s�����襱�x�
�{|'�Un ��\�G�ɲ���&���������0V/�m��` |���Ap�R5\�Q���,��s��Rj0'Ptw�ݸ��f��9h@�P범`>��	����(�bT,dc�o4�z)�thS�ց�4��FY�՘|+���f��T��0����@U�dk��EGL��m���t���<��d;�B�VA��c���������]|���vF�&��0nqb��Z�F�^]���	�T�i�Le9Mc|�x�9���(憒{4��&mBe�����ǋ��؀MdAN̡)� Q�����מR9� �8M�l'�M�T�I_@02Ġk/4Tͫ5i�����?��3\U�	&���Y@r����̝�l-�/�D^:����%僝U"�Єd� ���� w�tS��':�[Ā�l��r?�ur��xo���W�z&k~�Ʀ�^ܧ	Ut���lq��;���e���i��,.T��٭ͷ���u�+.V9	�z.U�*R,�Ǧz�0b���E���/ƠRAs������ `��&�Q+U�P��3'P��x��X�LӁ]B�*�߲�)R��JO���e���]Iy�)\�hm%Pa�=�~h���,�G��Y��yh�ۑn��>q���;��;ʿ[a�^~
;��<6g��LfB�����%�������ǟ�_:��t��+Zλ�E��6a6�,�����-!XJNs*�8�-�'�*�jV�T6�zRd�nC�|�7����{_��S�4�uҞ���|�j��j^�%:$x���v
�yr���������˿�+���<7�yZƑ�������<�<�y���ΣL�}��f�<���g���.n#�RI��;WR��]y��t���y��%�{hw��8�,���&����|8��zД��!���A�箇�>�.�n�^ [3|�:�����Ė��o��V:E�����Lc��7�9Hf<��I潓v������_�d��i.�LO{I3!5{��P���Y�d��i;��]}�fեc��ʛ�dWzi�����e�7:d��m_"�y����9��� �7���W����w$�#Y�Q�00��Ȼ��G��y<8KI�ێ���<���t�U7ѧ?��L��[�m.��;�XE>~(�pi_��֌*@3?a�\V���Nʠ�h2oL�^s������L��<�eR�����ޛ>Y��ay�}�UU�=����`APA���`�!K"mK�v���>�R��,��I�"!Ԁ � �`�����{��jy�޻�����<��7�S_����r�Y�����j�3ݒ�֚���v0p�+�q�*}��M��-���3�r��Z�Z�z����#X5�u�2�jA>�-�Lx�܂,3�L�m�6��οCo\��淖q�ʖd��n�9C
�L�=�U>�<9k���3ڬ��O����g����\�cM;����*�k�3���]E�L�����/��(6R�x��[��o� 0��{ٷ�ؙ�7�����[�v~6�ٺ��J�k��*|�7�|oU4K�i��F�Ĳ��w߻B�y���|����������Vή���W���� R6�I���W���Q����\�U��.��u\Of�)��&G�\/��w�F�t����E1]�?�ٹ'k�S5��?���������:qb&�w0�g�gẼΣTpȘ�:�b�:M|��%�[�Y���fc$�ys�P8�t|1���k�ꪙ�R��M^�pʍe���T��>-o5��N�<p(U`�YE��,�	���A\��� 9� Ճ7f$�m5��,�\g�Ae�;��>;
�`��մ�?l��p�A�V��v.N�o��sW�6�j���3pbO��ö���{��H/���ĳws�ڰ�0��w��[��c6� SV�y�
��U��U�}�*u H�9ṙ���H �`q.RUioN?�ɛ��Ԯ�p r�m����Z���ͧ���6�F��j�}�@������>��gک�K;�
^��9ɪV�ǶhL��d̂���?8@��̹�S�٪@լY��읭�g�}i�Zk���QP؎ɼc)�����'��^c[�����{�w�������ϿN������P�"�ٸmVK�Ǌ�A�S���,/���0y��*�e�� k�/�`ڙ|N�\�whtx�l
����s?�%�*k�?����`A�/�,�C���z-�ɀ�u����4��b�Q� ��fT�A[T����AմʁG�y�fKa~:�cR�y��rcAQf��<��_�s�/5�5jk�v�x~'m�US�l)a���::�n������6]����ڒ�Z�<��o�no�(@�!k%M�3��y������II}xY*Ì�DC"�VF�_�V�����Gmn���^o�۟HEh�y�`�+�e4�S���.������vnY_������/��5�_���y�/����`{�	�_r&�X�͂����~H�a>� � �)�U?x���[t�-�<i��1��]�/>���9�z��EU��\�{R�O��#*���S���{���{����k��S�ҧ���m�`��|<��|���_�3>��ضf���t��k�����۽f�5��Pj.K��9]��I�䐌�����Uے�\f@R�?z�٘Mx�͔��h�vu�H
N����ViA�e�Z/l���?w����Hݢ�����u��o\?w ��7�n��*is��n�oj�"����)��SsTdw�ha��(��b�߯k���?�4�z$)���	��$�\YV���� ^���A^˃=:srM�]�n�x�'����L�����;�2klz4e`�y���h�)R�)�?�뿤�/�Mڬoб㫴^J�E�?�"d����F���E ��{�>��jc]�H����n'Q@�=������Ϻ��'���}����2��AA&(Ӏ� A��s�ם��I�^8��n̾��B����gmL��m<(�R� �Dp������@��Ɓn��(��X 8��
;;fQ�>z��?�XB��@?N	3�uDp:��ѻ�5���qX���O ����w�F�C�/�������z�v�is&c, M$+s�'��؃z�@Z�e�>D�d	�J�,uʫ����}V��su�}:B����������}������E_s.ʥ���y���-����!���^��˜��t$���G��vƞ#��d����FeI�,?���j%Q�[Q� ���t{�gcgăz�Ʉ��3����={�s9Z�ԟ��F�^��b<$�h�Na��p���u�����f2�;�dd�  �����pCe�wB`�7��ݠ1瓠u}>;\���Y�r.joK#0"�+�J�=���-0c\�K�����O�R����
�I�j��}�o͂��Gy��������3}���������U��L;���0I~�b`8�Ώ)�O��yoߡ����:�3�D���d��l�Ȣ����ҍ�#��Ƙ��~ڿ�r��3�]W�>��y�7��ݟ�t�35�4`�<���g�����A���
�y�,sQm K��Q���m�YJl��{�:����0v�)/�����;G؁��o�;�wp(�����m�q��v{��$,0�d[g�p�o-��p9�ΐ鹿z��'��ƴT0W�^%�Xu+�.��%�U�*�$|Bu�=PU8��Ae�X_f������`ξ�(%J9�/�t�'i��T�����Y�h]����ƹ��;�#���p�6Ҭ?�p��Ԟ/5��yI�Ҭ���٫��
[ҶaM��#]|�}Z�S�=fw��O��mWk�~�Q���F��`�(�_q��3��/�W��i��AoU�G�J,Rm�A&q2��G�XL��C���7Hbb����ۧ�;�}��Jm�Ł ��3�M97LW&HZ�i�v��\��6���7�7ߢ��;F�y�s��Ж%�mV�(z$Y��n�)�*F��_�s��rF0;�s^H@�����~���nz��*�J���$�d�ek�WLL������?�)��׿f�L1$���`��x�O����.�s5}S�Ց.�':��^y�<�?��H��*"�Ҫn*2��49W����\�9?J�hny������ds��~���?�'�^���e�ߙ���\�"mF+W�g�ø@�6Vk�i!%��gP�w���d~�@D�+�kk�Y�*�ju����D�?�c��|F�l$�.����d|��D~� �c]܎D|O�]Y�����w�z�V+�t!%��������&3;��!��`�!'Q�Ll7����������v% ����W]���k��j�;l�)�Pe����D.���v�%��klm�o|�?I�w./��6���8�X%rK�|�mO1Pl�x���?��ߠ�����I��O�C��-�\��菪[�#L:m�=0d%��R����>]h�nkT��ǵ��^	g��������������[_��S �tJ
d+5�;����4��M^�[����U��i�Z�!я��&-��\�t_�:3l�}�AE[d@�J~���?�	xc�һ�������'�g��-D-C[r�8�͸=!?��H���J^�N�/n���M�#~�u������C� �Z��>3e[d�f�#��hǨ�&؇�Ze���o|�����)��X�WYyJ��ӕ����{Z�q����_����!l�-!e@D���D/��%Y�bm�x\����1J�D1N��]�4=�+���g�ɹ7/���f0�6trW���س��h��07�ѥ;��V���q��S������-e3k:ł����ҕ˻����3�J0,�f� �fC���UQ��7㌖������/���I*4��e�������}�S-��Ә:n��KTqB�ۙ��eVD��P6����`�������b� ��*�j �!tgdH��ܱpfY��.^�B~x����̍�	"n�*T��N���_�}Z�m1DHq-� �,�e-�n.��6���5�)�ϕnx����`"�����N�a��z��L_��/Rm��`�+n��gf�Aq~Z�?7~�/x�������uMd����9����(��#T�~�7i|�O�]�=���~J_�S�f��s�� UI�����U^t�h�(J�d�ג��K��9N��Cz���w>J>��s߃����J� ���ՕT��u�z�ӟ�{o�A��+���)���|i����>���%�W(��聃�ˊm2��>��5��7R�?������:R�1|�|��M ��u>u��bvrq���qO��_j�m_�s��}ݾn_�w��N���֚M��.�2�zD!��!d��1n�iFI�_��C�.�cw�-2"��0��v$E�!���x6���O�@�vpH�ܔ��Az�����w^H��q���G�λ��ﾟΜ��[s�g�`��O�>�Z�y�-�t���{�f\4Ŝ���4J���8��w����h!Hd�M�Q6$�V���v�7ޤM+ܯ
z �Z'E	˜R8գ?m�LOD}���bN����%�ช@\�d�����2XO��sX��eݗW6�% k8�$�d7B`I�D}F1�~�˔�Z*��g�iPξ<�^R'�ܣ˪��$�S-P�*
��Ef/7�����e�<3�r��Խ��՗�����p�����ຍ���P�ޫ+����X��L�n���=Ba�4U��1�g;��m��೉��D��5���ܡ�l�=����0��#�������#Y��-��U�ͺ����@�ﵕ�H�a9�F��@��2�uY��[�u�������(�i��u��AOokD �Tk8aN���5;���Xr��Qi�Kt#K��4�kA�_k��W=��^$_��f�D?y�����h�v���;L�|��c=f��}�L�S�_W{��п��ޙ4C�{/V�z��D��=-�`�l�Y�fz�ʨB��������X�J���1m���g����Q�ֲ�������6=�wF,�X�����F�p��F����zl����
E]����L$?;:6���G�A+ټ��:o�<+aDa�&�������ꄐO����n��&��-z7W�W}� ����>���iTE	���͎�cF�|&�n�;�D�T��;q~�$g��
G`��N�&k��~-��o��`c ����v܀�������
	�Fz�?�}�\%�	k����w��2
�ި��f����ʫ�%�\0��� I |H[W����p�,ݪ=v��ͺ�߼�:]����A�ߐ��IQy�F�sBu�G�U
(tJ��?�PT`�Z2jΝ�,AvZJfu�L�S�J����e��:�j�}������{��W��]�=�S.�8Q�x�5tqB�Q��6h���X�%�-{��xSB��y����}�O@�x&�(�F��ڇNV�q�n��9L�<.;Y�8��Y�@�!����N�y�1b'��r������]{�B��G��Y>�Ӄ������9]�|M漼���Hmn�����O���b�A"��h吃���m��gI������\WX�N���ܚ��������]��,Gd�
 ��?>�L�H�R��?�}:8\K�{&lv.��Y��H��"С؈�������#-6���'��O?`��P�jxR�����E�4���L�g��~���2�9P�6�w~����9p�Y�<����d����n��U��.gm�Yx�߼�}��&������NtF&�N����җة�̳���3�������Lo�A�j�WnJk�T k->���sܪիm8#�og�s[2|�O�h�zC?��K�+����h�4���+�g:.���H�3i��^&��l�~E*��-� �b��DVL_i����@��Z�sK�y�"�j
Y�o�I��-=4[�-G�'\Mq����{@?n�{��h��W����x݆��xM�p�6G�JH��
n��
 ���:e�����Wۺ$i'�I�m����+E���gx��5�d���M��usE�N̤r� �!���Q9���`�Ϻj�]� F����|���W��S�A���_��uS#P�3.�=r��c{H��.�=�7^|����/P�&�\�i!|��vS�U}J���; `�ΪM62V�NM�#�B)�W ��T}#��xN��j{��ʖ�Jǒ�  MIB�ǪÍ�g���jg���7�W��g�~X[4̍���5*��
K��d&n�g�^�v�e�J�q�`;8��@r�����e�-���Qe,��l�b��*�\@�پ�`����4�n��!�՚^�"}�+�������W_�3�26�!؂�"Ϩ�������k��,�~"�H�vpV�����e0&�O�ʅ� �[F&�G��o�N o�WF�og�O�߿���_!-	c�R��X����g�@�)�G�4��O��Zf�����2�4ߦ���Ґ2S:�>Y�t:K�O ժM�t*���")��Û��@�Ͱ.EtD��ꆨ��:�����!�nG�*�l�e� -&�r���x��7ߧ��I�~��R��$玫�p���|����lź4W/b0�W�;�������yL��
2U�?��!=��u:�_6Ў70�&�Y��~Pdx��K�0Og�}�*a,󊵤P�FJ��MP�{2���<Z6�r6!q������"�گ|���|��#�1�.�'t�9LF� D�_d�C�N�c��euz�O��M�PV�?��`C�d�(�m1^?ܣ�o]�'N����(���to��`Va U2�	bT*8�>��X���C�K��ܥ��J�3t���&c��'hk{�f��%k��:���ݺ�!�ߺB{{6�]
@�6;w�Z��Kސ��:�$'3[s��@�� �L��l�\b����zI/_�B���D�Y�K�*0�Q�K�������#�[u~r��hH������u��ۯ�; �!H���'ݱ8�n�^mH�,8#��l����%r��h����\����g���a���GO�r֞��~_es�&���r�Ċ��0r2KK�����l&�P�fE�.ޠ.�$�p�u��-)_&=��t��^3(��3[D�+�Ď�.TFu�sf.[?��i�)!8�9������@(&Eu�E?��>��ڥ�����Q3M��0FpA�#
E(��)V�>���
x���^�IROz�%�`�xP]��|}`�=�h�șDL@�{�|���1G����K�3�sJb��-��kߓ۟Ǥr"KF�c��Y��u]5țsr���u겸K��F��1�"�i��W�l��r�J�|Ś��X�ޮ�$tK���Y����7x ��wa�� �:�5q����`�iG[w1�H�+�}A��-H&�l]O3�'�d��bR�9U�|Nx�J�{ 
_��c����r��Z�A�G�c���:�/�����@8�h����.P4�n�� U�7 "Ψ�H����M�!� �F���c���Y�����Hf��3@>�2��|�l�L�9տ-�\����r��fFx%�A�ya�}���g� Sy?w7��F2jI�� �U��4ޟ� ���#��5��R���DV2�i������o���A�8�Js�Wc>GnWH�w�I
�H�9u����ԏ{rS�X���չ���L>k)X�Qt�/�V�q5hթ��e�W&4���j�g�������?��2\ '$�Ӝ.@E� ;�b�ϼ��;f��6�T�N�AN�2�J��w�M����'ϱ�M��j��oy�<�L�_]���=�(ټ��eӍ19��y���t�'��^���j�Oҙ�c�=0Y�U�)�e���`�º��K���ͥ��Q�3�jﰎefk  ����z��d��`9���ާ����d�K	�!Y���X�9#�A�����Ñ��X�d�gQ� �$8���o]�
cp� $g��L�z��SV�+i�Nd�5i�b�,��"��ܹ�p�Q��* `Qc.�ۢ
Ɲ�dm��V�t��17�??nT��`������4 ���c�D�03q��>��������+�0E������so�g�}��i@
M:�xh�&6SM��y��%��u�D�� ���w�q�Ktsw���N�����q�nYY܊���zB#d� �d�5�ތ]�z��ϭƟ�Qg,�m?	J�`����6�U��$�xT�q{�s���b2����$�,A�VݰC�x����2Y�  x�9�jЏ�{��o���W��!=��ӱa`2&����鯶G�Μy�c�R���I�R�>[Β�7k�v���W%�Ń�W �s�H�����DU˘&��=��YW���ʦ��uz�������$Y�9l[rA�V��ds/%l�dC��d0�jХ�J@U���~ދ�Y�pHz�2�T5��w����9�}��7�üf�2���ކ��!W��!���)Yk'�`	e�~e��3j	����e��Tm�Jg�d~����]��j����+���	X�l�&�;w��z�9���19G��8"?XCj3��Z1F��z)M'�S@�H1�e޼��T���=\��F��!n +y<�xfI[�,L>r&!����|�����=�-�2n�D��	O̲^���{�͌3;.}��*{L4
l�m-��O?�ڄ��v�엉	k<��g���h�>�]����3wž�` �,�6[�]#tHv������DZ���Kf㋗L���������o_�Fi�T{�j��n�/Y6r��lK��}q��6�����3���1�ŃW0m��O��co���H{(�L�N/��cZe&fA�����<TZ�L�$��Fw�i]�7E�&�+L�f\��n�s{&T]�zC "~�O3�e�C��-`����/��uS�$��H2��jIՊm�?���\�*/s��>��" �l����<o�Lz܎�A��^}�"�����ಂ'���K�+���{�{?t	71��>� ࣵSQe� `�eE���zeO@~Y�hi�.�=#�׳�벺�<�mR��˯%m?���pUE���'3�	��@CF�ddg����-I'���2�|H�l1���z�����Y��V*JM�R���#��*�u��m�^���7ߕ`9��+tx�#�G�4���$0X�R�3��3���We��^�D>q��W_=��(X�+7�n�ۦ�Ks�Mޗe��"s�*=[lw\lvP�VEi� ;��a��(e������C&[����i�ڐ)�y;����,�N���w��Va&��BtZ'��_��:ݱ���t�Ԍ��r$4�T{?�4' S��{Fi�SE���Ǖڌ�ȭ���0ޤ���v�x^Tщژ�g#d0���hM�_yU��ӝ{M���(3mo�Vw�^7Y����k��m�K=nD	�]�TB�2�}Q�&�끎Փt���r��6��n>r�n_��������� �S��V��n���_�|�/޻|X��y<U��L�����Q��
Iq>e���*�]i��_^x�~�O�l�AJɜ�ʀE�.ʢ5)��� �(SȉhJ3�]��g�)�ܛp��d�n� ��a]����@�I��"��F���Q/'��?-}�z�
/1�)/J�9����@u����rE�]~�v5��"G�j��4�K�Ρ��hOn\�HK�ޱY�x�P8.#�E��U­��#��L(F�Ŕ1�!У\>hk��o>u堗�La�f�DLȎ3#���z�@�.M��܈J�V̮s��X�J�àC �����F�X�����a�˺tk�������P^a(L�q�uEIo8$����?�ȳt�v6왡4}on&��� �:�1�aQ��|=�(��R7���$s*�&g�# m�xNMAw9��>��ѝ(ZB_ײ�3[�.��}�c`�ZR/{V�E&܈�r(�������ڽ��Y�x�\I���dR�;0�R�w�C�q����� �$;K�In��v��f�Cc���Ԕ��m�n|[�5Up�n/�T�. ^�Χ3l<k����?eY%��i�� ���G"�*�p ���Kd�FVsl`��zЗ�v��y�'��g��c�A�2���kY[� +eD67�j�l:)��=�u��k����͠v@;oF]�L �Y0�;�a�O���~;CzE�a�1�^��2�1�jN<[W�M2��0���� ��4���W���׶���>�C�|AN�W�	���]5�jY �=��B�ȵ	 +ݍ���Y|��B�Sw;����d�H�=�L�1D�b�9��P�����y�>w[o󟡚E����'z���u�d]�GAL��q3L���+\�k�@��`S��zBu�?�c���x��'�ٕ������JB�S5�~B����������P��g�fI����m%��	�=��(K0h	5���2ЕK7(�4ΩA"(��$�� �G=c�Qe˔h����"�UW����P1�r���T�i�Yf\&xn*� ���$�(�q9�v�&�����v�|� �y:�9U+uUg=�N|�� T��@=�zq� -�zs)}�9�&�����V���^�G��s�c총���Km!v�}��q8x�<;�iY�8��p@V��bzNE �3�H2��J|�w�yl_h@H�\
y�ᝠ�����an���> ͞><\�!g��Y�ZL��Q���w��/x�;`E~Kީ�=/<�7-s��|�z�n�+��skg����@�GBi�}M�K�ӶW�^ C�F�Q.�t�)���影�#�o[n�>9�{г��W3�.]�����o�eY ������z�}��;zݴs��(�._�G:%�p�e��;aÑώ�%���iP�3��u���E��E��'䌶�}��Hgt(�g�NT��ʎ�ٕt︪�4�K��I��6���%-�t��o�G�#Y�T]�ګ��:��&Mb0����s����E�G[oh�D�%�%i ��d �*no9��C+I6�N��������ץL�8�K���I�bq%���@�vz	l"����R�IB��i�>E�0���U����A����%�C�2��`&�)�ު>$��F\���L�PR����R��*�.�/=:��[Κ�n-&t>�6E��ZpL��6��՛���]���������|4:W��q���_�;�< �<�g%�bG�.��H�9�~d�`vS�d�Y  � /�����.O$��0���ꪶSɮ/�����{Ҏt��E@jO��$�S{�[����k�d�ٌ�hSe�h`��Y��J�S���N�"I���7��Uƪ�����3�B�ʢ*�xw�n���P����i�窚n�7���ԫ���}*��H׏2ȜGk�
p�����ލkK���fi	#�B3�(�.&��@ـh�R��|D�K��%�����b`v;s5|� ��#@ڣWb�/&�7�T�oh�[ѥv��-���������0��2(����aQ,Y����z  ��IDAT�&�J�I�����'�����8<�j~bК����1d=�xrYg�!lRZ�Y�LE��֞5 �6�7�:��}[G^�nk�kxx86=h�N�4р�dc�UVi<
oOu2��W��&A�1z�-Ki�����vo������1�,x���r��;y�o.
��{��>(�pF�P��Y��>�g��L�C՟�1�.��YO���+>z���7������/U�7��Yn��0{t-��DW����]��ǟj˼����3>���~]�s�dL���$�oӞ��>G��,Fg�3���̡�$��_KZa�	ܛ鹈?BQ��(��0wU��S��IU�ؖ������j����zsy����
�n�z�>�^��h�B���xg:�������3�'���X�M�]���u��}�7��; �����ŭ���?�t�¹K���m�X�ab�R1�5������f(�1�^�o��&,���y��Ǟ��^c��f�֋������=���J�*;�"�;�$��J酨c�iV��J�A�����_��Q��#��*�Rz1ͥܛf���g�����Q���}^����W^�K	�]���m��AbGw���̆���Lߛ(C�w��wT"8(��__���P"����j�y
ŤS�)�&�ˣ+���¸���E��Z����B�"��MΕ`/g���@�/]��6�����u��L�<3g�ޫ��g�z���p��k�s2F8S�l�H^A6�oLW1@v<�\`@t�Ha��&�*�x|�ԍo��nm�p8X��b=�t�Ϩf�ҨJ��?P¨��H_'�D=�����Q:�e�DB�IR4��;#ŗ�7Rr����)Ց�JM�or�ґ�� @8�]f��O>����F�z5�����N�����|�|���[���B��
#�b�S�$��hہ����O�Bm߫����?K�P��Vo#���)e;h��pP�<��H)���j�����d�,4�;:o�T��7�Q|O�0|�	n�~Tn1 R;ú�˴/b�Q��o�� >z?�����v�j`˜��=�Z�����Vr~��B�RE�2�?5c��8�3]I��%ӝC�y�f��^jp�����ݞ���@�?�4���I�XC8Px0R�w�=A�bИ;? �j�~���2���u����ƫ=?B&=�E�d���|���&�?" ��Q%����A|�P�1�wu����=:���Oi1��$dst����N�6i���p&;��_��k)R�$kūJ�(t �Ś��JR~YW��%f��<���I2��)����s��Sϋ�&�G��s����f	aQr���Bpz�Ax)h��@G�B*���אU��g8`���{�M���f�;N���u���;�����#ȕQ����!��d���y9m�� y	8��<����|�VȾ�V�`r��0�o�?]L6^rr��<�y;����,����3��U���P���"k���,����!�co2�Yp{���fi4�Y[�������7~n���u�(���k�H���G'N���� 4O�;�س�(Q�,J��n��:;��"���@e��A;��%(�ϕ���A�i� �^��xy>WJ�OJ�9T��#UdT��5�w��uiQ�&���_T��J)�]�K��l��Q�lԠ�U�H=����8m�\�+;<��ՁeY���|��S&:No�=2�D7��8�+�SHf�\��m�d�IՔ�F�7h�=���j=��;�]�h���2ڕդ��<��a����t����ԯ�	|൬ т�Q�@��Ř�:�m_0 ��5�2ge��+��[���6_r��~�`�6�'s�c�l����Q	 ��6�i�U���,*�3؄�a����-4���zC�ڒ�jq��j7�x�I�K�:�dmf�gƟy�7o\׶�X�Y{�z�r��݃�;����Q��!t�L�M6
�E��y����XNq��� ^_�su�Q�-J�{J�w<�ݽ:[:����о��Md��<�U��! p?ª�u59�Z�¿6�������~��Ơ���?Ƭ����=���:i��]��G��kV�>&��������y*�;A�+Q��l�v6����tx�g�>��G�[x�h?�a_qU�pWɮ��1y ���g0���Jr��D��[��ZU�p���#��`ߡ� l��U+`�����U������g�+�7���g�ylY�A������H6UB�"dd'�@'m���7˪�_X���z���؟g@�1�ꭋ���{����hr+c^ I�^�y$� ��d G�� O�\a9��>9��f�x���#�#i	�%�U�)��b���)'	���ߥS�N�s�f�V��N���t3��]�?���Q�r�Ƴ�X�V����k�Z���⺑��ٗ�m�t/�|��6�c2��RhC*��N�����i祷-����@�ΰ���5�i4w�=_�~M������$�����zӅ��=��Ok�Y��<ܢ�H;�ߥ/�q'k����E��E}�VU�����-Vr[NA��^#����:ʸ7��u�C�*���f�Mw��R� �� ��r9�����>�7���L�����+t��^�A�irUڪA�� ��H�Q`v"��Rn������;_�����N�Ji~���-�"X���������^?� �*��lo6���������<����Y�;�>�h����Òu�:��|�}��'i�Y*ғo�4�*E5�|o)ɔ���ܾ�,5�:BPF��6�g�iu �@����O�0ٜ̐1͸ ���G�z6���ګta<h���ב�ؔ�6?�y�J%�䊾gH��0˘'�i�����;�%�HaC.ut���Q��=�gb�h���N�>�<�*�c)!�L��Ȃr6������`x��ͱ����{uZ�<{�-�2
���3U�?m7'�9�O��N
�P�-��@�AD��NG3< ��:e{u���BC!�EW��`�5�� u��@'��ɔ���д�q�f]��ޙۍ��H8ua����?1�����~w���+O����A��_����C�/�4��B�����sG�R��)Q��Sɪ��eO���Yr�w��IY�(r ���U3�wx �F����{'ӑ��ۈ0��_ա��|8��&W╗v7�K@
y���m6@��J�bMb�V��#z	r!u�꽊�e&=��:C�@�UC���$YZNhjĹHpV����ث"�9���>��a8i਋�^�D2�4{��c��\��]i윯�G�]"�H�̠Ag�D�̓�W{2����ѩ��sE9S�ΐؙ�'88���T�P GzG�2���]��"T������ͫ�=��|�?�~�'�:9��GxoW�Q�r4��8}�x��s�Y.KLe�q:'Q��,|�j������n��<n�g�!���~J� f�k�5M.�q���x��C��GC搨��9��1� �у&�k��[+;_�iN�W�r-�V�tikQ����X]/E��Zi2>���y�)o(c.�)�s*��P���a���t��������um�{�g�>�C�x�����V��V�5��(��WB�b��8������F�1���͡�˱���QA��k\��'�t$�5��MeA�*�V�j�H�D_�d�t:BW�i�|>����m`����aՂ3��̼�+����e�җy_���8���������(hy��T�_�i�����tb�كG��I�'��HKV@3��6��_c@����o�]�f[��]a����|{��*@kV�_���1��P� �hO J��&W�CF2f`Q�"`~�҂{]�t� ���Ї������X��*�a0��l��O��ˎ��r��]r�^{�]JGx ��j���<� ��W2����ޞ�|� Y�c��P�`OGhV��Φ7P͇��L ����^��s���UӰ�P�g�/��v��e�5�9f�����E��@����ȷ��Vx@PY� 0�Ž�Y�?����v�[�|�JK5��=��B(Z��o��azg_ih�r��E�����V�HIύ�`���y�1��p9�:��S����&�MS��X@_�?B ���\_2��.���l��^�Nl���fsx�<�S*�����=E ��\L����{�玃XB)*��I��*�������w?s���>�H*a��Vd�������Q�,�W?�w'*܃&6I�}H�	δ�)&�	�
n��VJ:g�5���/��;�`N�р�b����d��r�~�*�ݯ�Uš�5�mƄ>�6�d6:��g�WM)��U�$)%]��ús|��ѯ#.�`�s�1W؎��_���t�؎�H6`��ucz�H�\�G��/�'#"���؄������2K՗�����C�x��JU�5�Xu*IG��,�UTc�R��y�a�ר��޶M��cS�P�� fl�֕���ki�R\O���/�,�mM2T'-Sղ��)p�ym�
I��:�� @
��.+*�|tz��0暔�1�P������|�"k�#|s6�X�jz��,��T4�4_d��76�8�Nz���y�VJ��l�k���ۚ˼+�.Z���k��X5�%������ِ�k�{�}�B�9Ϡ�ⶌ�z�J�n9#`:-����T+m���UWV�0��27����~$������s�lu?B�� ��S?s\�3��t�VJwJ}2��-�ݭl��`n}�p�]�����vN�v��l��#���U{^���M�肝!yPt)x\I��3U�R����Ht'�W�`�>7|F�~�"i$$�T~�J zM���>rmk��~�m�9(�p�i�g�����ܮJ�0�'^��>�Y.i}י37��1��oK�Ѻ}ݾn_���u�\ �A6�Q�r��-�p����n�_Y�6e<��#
�	F{r6?�ج���0�~��Wn\�c�w�w>@���5HϮ�)��l} !(�<c2�����y �S��R�
�eܓ+��I8��Y�9꺐;�}ֵ.�K�æ��);/}��zp��$}���.e���fB5k�Q�TVʇ$��w8L��]�*}v���`AwpP����1�����8�RQը�{'�tܳ�1��}M?��ږ)h�E����n���yI��"S.2�uϠl¹oA�u��;� ��=����L�|�����;���l@'����?c�{�"О�!
f�/}�Xu��&�$���L�"<J�{�o�ї���[�Q-�r��J%�7Qb��6/�u�������*e�%���g��n\V��9/t���hT�OV���j?()��ؘ<��v�I�����*]�,���v�W�����2<}]�X�yX�믍�f�F��giKB�ṝѣlX3a��W�� �8c���(ʾ��U�Rdʐ �0��0X� �iP��@kT����%�G����C�Ed$ (% ����]0 ��!��Gu^۝)[koOb�F45~���y5� B�>V� ���g�G׊��:�q�1O&∩L���s'����ç��K�F[9_1>���П_]��Ɵ:y���
�8��x�x�,��7u�#�[]H;�F*�FP!�9�L¨�	'g�8�A8���	29��_M�(���@.#�s28)}lF|��9l����� FJ\=�1��1=_�s�8x
H������T�O��y;s.g��H���W!w��LY����t�6ѿ����.�;~�-��y����3�s�5Qm�]��%+�36��	����#�d��l=���'�,��A������>rD	dȯ�e����?�=s\����h8�1�p�`�>�b�g����X}a��im��y��=����s�_P�g�`�X'#6II�ݗ��z��*������򯌻ĥ+c�@WZ9��H#���e���3��H����Pi�Va���qj��Â��JC�\]m��D���y�2\>ĿBp�ȧ���s�=M��h��4=߱�3�g
:�� '�j&�d�8�b%xɫz�{��f��p��*A �7�����w�E��Qs������bo��׬ҬZ�t���j����%+U}+[樜�9��,�H�cǶh{{�v�F�<�Y�/��r�����?�V�� �=����h�8���+�����`��T�=�__�$=o��d]��Y�gN���6�fS���f,���	�~)��CV�����q�	"�0�k(Y~�,�M��ٌ��Q�&��A�5��`���#��q�]<����`_<�J���` �"����ڴ^ׁ����i{7o_8$�/G;+�fJ�%y�g2���:�i�0x�����@de��|�^��b�&�j�;C��VF�%���r�ꪇ�y�aY+� �jO��e��ƻs��kΪ���K��}�; ����b&{z��w��$�Ԕ�T�D�����ίUF���lpMg�J������pJ��vJ�X�Z��tQe�V���<�@P&�LV�$ϴZ���*�g���W̌�s���%AȬA����d��&��a�ޙb�a{@����;�@�&t�d�%W������3���l����h��&�6����j>�����3'%у�u�U���Ku�z�7]}J��� ����N>7�*�_Kw5���F�
�T@&*��Z2Z
�Mc�2�Y���8q�f�4��T�)��ۨ��ή7`�)l�^'֌\_����U�X'۬����ݠ���7��@�3���B��E*V"�ee�&?���L��I���NϞ��$dƉ4�^wt��@Z|}3Zo�p߽wI�)ΔW�yڴ�8w������rd����ᇝn\���%G�E:]l4>(>�a*��zw�/����'�x��� ݆������� ���o&7ex<�[3����Iv�j���,���<���-f{Yj����(��G�7�z��֢��t��R�����|���F��YE`<�{��;���'5��ASCv�Fn�������QՉ�&u�Y�0z�?��_��k�1  �6���w��5Jr��ʪ�.���^���:���t��1�jsf���up�&�M
zN�]�VTF[���
	�%����;�_����Q�I����#�YR^AZ3p+��8��(�F#�o���Tq>�JF N?fY��`Q9Q��� ������cl�ӧO�h6�2�}R ��Q|��}ݾn_G���
 � ���ry�ͷ�<����r<Er2̡벌"S��\Sf[=G�U3�7�7}��{RR�w?H��ZY�����M�%U�E���b�^)FI��i�����?�&�Eσe��/m�eՈ��%I;:�b�Ƶ�K�Ѝ��,J˄��L!�y�L'�g�����1�L��������$@[:�=E�/#H@SǸ�צ�N�1zs^�psc��9J�-�R�����t��;����x0&�֨;	Ϭ�9�%d��P$���3�	� �D� B�"~0�ݐ�m3~��n��r�K
�(�5�B��r���6�W9�Q'"a��9�,��z�b���D��E�zQG�2��+���A�i������G�V���*] 4|}(���`wϳ��7�_N���)�ds�4F���#��
h�Q�����K�&��)uC��)�7��-�FN_(�Y�c���Q ��ut����d%��|���@#� �秙� t�J�C���<J�� @P��x�5�Sǅ�Zw�fuJ!���o�/�������=�Ä�G0��z��a�	N�c���ͪAӝ��� a�fe��FvH��_� u�@�p�oB9�HM�e 1۵p �x��~g��Nz�7^}$���t����!RCwA��i��K�V"��c�nR�=�y4�ۜȲr:6�0Z訑��2��y�@��?���@�0�����=ڲ�N�d`5��>>�-`v��u�|q:�F��C���.��B��5�r1A�ȱ�F�Z���kPZ�����J"/ju��(�� +D�et��
T�'E��G��Gi�߸?/�`h�%�d�ku���8#��sם�%���"�X��8��S�	 ��9��(�i�m�*0&Ͷ`��v����$��"|���%��ŝM��=$����$��JX�/*�5徬m�z���3��B��k���K5�Z��?�Lv�s��U��O2��c�>@3��c@d<6�H��qF�  �����)u��AA6�TA8������@O=~?���y:l��i�Y�5璺{v�v��;]�c3q>`�ku�g-,=�������g�H����Y�@2vN�]p�о�6#	��z�A�n�9\j�- �y�,��cs���ns���ؾ�_�D��C��e�Ѫ�\�{lh�_H�^מ:T�V��S�5���c@���"�k�\��w�y��]ߧ����D�x�����<�:�����3���j#21K#a~����YbߡV�+����c��р��#�5�:^��̰��8H�u�g��Ir
�U�����晄Ol�q����TT ��=JRg9t���<l/3}���U�8ql���NfrVjЛ�P�{����u#�F3	�k0zv琋�C����?�p�?Q����7��()��\�g��k��3���x�*��E[��c7Y�]�^#C���ު�(lr��(Enr��kI����Q�hc�����;J�s4߁�E���Gvv��X���ښ�N�Ȅ��[�LO?��fo[Ya�}���QP��es�@zq��S�i�5 kuvlcS�.�7�o_���Ͽu��쐓?�pL�g��qҞ�CMV	��ٓ����ễe^��� s��=$�,._8#D�������(i���%����	-��<����Z�7_,���m�~}�J�"+P��������A�m~'Ξ�����t���Zh��	��j������>>��b<�?�Y����Mg�l��rFk�
M��Iz�o�j���S5r4��n��p(�T?���4����O�.�;��W�σ�;X���.�ө-��0���g��eA�d�r�·<#rxȚ};O٣�I���Z�%��[8[y��d�QX��Y��-�����U�J�j�'��V8E����(��a�Ƙ8]k�+:�(�ӡɁ{�=Eo�} m^7����KeWi]@ �s�A���ܽ6g��V��|�6����ܢ���Vu���b�u� ����^t�a#Si�$ �!�6�$WWI�k
ش���'��5�r�$�>�ڎr8�x�����eڬ�4�@��g���mf��u�,��G
;u���݁$*ػr�����RfM�.],��e�}�^z�'o�9Y	�J�%'���}r�72��x�V�M
`H���p��N��2���;W�,W�}�ܰw�.���3V�� 4\�c� p�w���vNn�]n:� eߗ>k��{����>F�%���I~r{�4T�W�<�@{��ѿx�,�\['����Th��<Y?2~X J1���G�l|�W���
Yr����+Ŋ�����R���_�RԳ��M�4��������W{��>Iۖ\��
?V
��'��r;|>�Ɍ�&�A��/��iՒYB�M�gyY�m��� }�ʇl������J��{�θj約��Z��lz�X�KP�¿K���$����,�yv��;gO�;i��!Ό�n_������o�~� �j��2����3�g|v9[o��:�.�:�p�@�'�H�e{z_�d����D��M��p����V��1$���!�PQZ][�p���u�&�WMVT�ս2�j�d�͝Ѝ� � J(�Gj�7�a#=���Ht���{�^��;3Z�%sމӾ�x�(mV�g�pD@}5�����+�3�����;"�Jn�K؊�8.�[;�4������#8�����)�PJ>>�����{ăæU+)襷S(F�,���#cΪ�kvp1���s�:��#SJ��d�Sf��"Y}(7Kl�+_4��#4'w�"�Z�ȁ1b�̩�,�JJ�(`�Y�(�P�r�qO��k�m½}�k��"v��CJ�:`l�g�%y �{4����C�E���ĉ���	*���@/�Mn��T��o]��zʃ6H3�U����[�Wo���d]f,�|`����ʚ�12_z^�0h���y�*��S��n�s��C?�"^::�b�d,ܯ���Y�x��A0���%Ψ/)J��I��|
��F���	�f��`�j�B)w�q i#��hAD��Æ$?O�|q�[��n��b��j�55$�?� ����� P����@	Ŏ<'����.l/�;��4���e��l�s�ĠB�Q5�!������췯�=?Oˋ�&�4��l��|@BP�G������p��1G&=d\w>���ftIy?�Їp�z��SS�a�� .���V�O�ѐ������]� �%�C��2��>��E�,�{d+!�g���*x�;/ļ������8�p�Nk��;�$KE��4=.�V�v��:t	����O���G�Ӑ����(u�]mO
*���'�J�C ��b:M��%	�?F���v���ť8��!�1�i�}n�q17c���6_�sG�g�d�?��#t��Ľ^Mso��fR8l������Н��ƃT�9�)4�m ~�\����H�~�.���{� H�o�,A�@����u`�,�i���"��֌>����pI��Z���MΚ�^����̒
H�����X��Wy�͠��������Hc��K�҅si�,�&���8�eT�8+�jd(J�q�Ӳ=�V�y�-�gݟ����}�|�lTز�R��dR� 	�N�C�}���7�jel�)9�+sT�r�B����m/�/(�ɷ��9�y�>C��:5���u�o���?%v�����l[�)�@}��}|�B߀�YE�����L=�/Y=@�i�h�ܧg�y�ν�����3��9 ��珸r�f�k�Ve�ݍ�t`���D��z=�d������ԪfY��jCS畮L�Νbt�X�NEmȜ���/�D*}ׇy۷3���wЅ��R^�i\�5��-L^���}-����QT�b���c;[��ktՔ_���g��w��������[�j:L5�,�1�J/\�E=eF�k��pj3/L��=$���y=ir-��hy6� �}�׻���6�f�s�'��ud��k{Xd��<�lv��T�gD����E���S;�W��ez��~K@T�ڋ(`��&�UD���*�8`ɲ�zU�Xf
{聻鮳�E��<�M�V.Z�7l��(��!��T�R:�FKhC�����h�io�^���tǙ�t��]Z��׍��5���8ڂ��$H��X,�n���d>��������ǟ~��C�*&��uD��wN�<U�eI�S�,�ۺ.�U��f�;3�Z�T�䧲$�V;w�jI?~�|���FUx1:�S6z����c�f"?s�vNk2�H�:I6����|?�z�K���Kb���h>	�w�I��� ����<A�_�&�D��<���<i��m�̘�����[�;?�u�6�y�ǃ�K�{F@Y���F^s)�=Ⱦ!b�mc�����F�*?��I�cJ����Xә�'�ë7h�d��v�x�1r�q�fP�~ӵ���S�;����7�`�:�ȼ`(���њ8����@sAU4T��MA�,�_��?e �lU/X���_�2�޿�#��@�����E���p�u�R;km�ڃo���X��1�:u�����7���3r;HA��ue�q�'�$�QW"��sEQ���@�\�Y�2�&�F=���=�@;{��d�,�l:(����Z�{2Z&ѥ��\# ���X7?s� B�<W/��j[�~�!��#��q"�Q��Df���z����
�R�Et�uc �=r_۶�3m�z$�s�ˬ���G������o�xլ}�˿�v���rEϯZ�G}lJ�ɪ\:h&k�9)�G6�n�}�j;�(�	��>�x٧>�8�v���ԆT���s<��>�<��
a$�d�)�R��7�AaW
��3O?�zW��#��Q�}L�2�a��w$�?�H��_Q��~O蛒+�nv�!pF��Q���۰g�fE^�����$�%���&�����=A��>�d�88[M�o*�}{EAi#���e����bF��K
ʁ~�\�[�|�\@��i6fc����Wޣ77�α��W�]�hy�@�ÿ�z�VP^2J�[�����������?=���[[;7v:MG6��u��}ݾ��ϻ 3�y*����w{{����g��MYφB��48wz�;�g��U����Q2��1��뗩���cO�f�jBr�ޝ�"V�b�a5�v���5�� �����٦�`�rOp,��eJR�����e©�_]�`Tsjqi�7n]��w����h��@B��U8+ȝ1^6�Ό�G�RB�S���ݿf�+�<��'��]�Hp���(-��GP��ϖ��>�qЗќ�9�2�s�:����� ���+���gk���(�O��A�=wFt�L���C>v� �s�"7b���b��9�z��s��h�H�͡HO�~/��a�k�
�C�RV��8���;�;���(�/�}�N�ł#S�[�D�9����Pr:���R���o�쑍iB�oJ��h��*�Ѱm��A�Vy"/�W�J�g�h52�l ��s$C�Qt?q&��?Sx�ߖ��{�q=;��:��V��a< �S�����YG��ߥ�[�&����.I�4ċ��|��?K\o�x��(d.!o���{j'-�=�1�e����o�����±&%������J��0:H�7@s}�ԃ�ng�I�WN��q���xF�xb�m��(H`��@��sc��٩���H)v5�O��4�@Ɯ��x��Y�]f�dh'��.:��3�c�F�=9ʻ�3�4�F�.����C�/ԱHtt�P��بt]��ԝ?�z�=R�)LϞ��jzT�j6Lߣ ���P�m '\֡������ l�?�Cϫ�oQܾ�p\���bw�~6C��*�9d�w ���zJ�+*zr��Ǵ�D��ѫ��7��ڟ �6m}U;^����oc��� �Yz %Qu�fs0��9}�����o_j�S�x�|~��v<Kv)��L.�yk(tk�`���X� Y�d�{_�<�B5��cQ�h�S��e&�����8cd�9�4��d�A��y�/��S��޽Ҿ>PY�1��-:�{��{F"���ǳd��8۹�o1���~�|�����Ī�r3jg�<��9����d%��#�d��;QM���uM��#t�����f&�t sUv��Tu�8c%���^��9{�u�A���fI�t�K����AhtT@s�9w������|��M�	pP~#��Q�`I��df,�-}���Ʒ���lrξm��*�v/�\OŖβ�8+���KQ`����G��~�>�®c�Y+�ġ�e�k?Z��b��+��k���B6w�������4{��Y�����}Cc;h����F��(H�#�!V����|���y�L���E_�_m�Ju�ZU^�Wk=��쩐��@�U݁>���� <�:�?g��Ĵ�>�I���_������kMe���3p�gMfA��v!���}v)��sj���fC�˟m[���Nuے�	�7$�ʾ~/��:Y�/B�������(>W��9y|���q�?��%�r��3}rF�e���y�UU�-�7���:ɓ�?LO<�h��C�$n-"&��eTi�:��*����^�!;�d�a_�R�ˬ��O~�����<�a��J�N���ؙlgtξ�0(��ȴ9��q��ւ���ϑ��)]����t[��N� ���O������̧6��7�Yb��fM��K�?���mMgt8ks���]@7�\Em�����&�o�Io���F��v�����jӫ�j/9T#T�YxJR^0�jE_M�&���������R/ϴ%bmg_���jC[�~����t�{�S�X����t�Ud��̹�iZ^�1�$|�O=.=���q6z�R+�I.�-��e�&��O���C�OMr���a�W� yΛqE��������gZbg܌M�+XJt�����y�@ޓ�� �:,d^�~�vH���� �V�o�Qd��+�X��>��b|��>K�}��)�"��8�{�=�@���_��/�=mfsZ���>�'M�^>�E1P�+o��4[�-�lQ��{��O>j��#��RHfk�4e �:�`��H�f L���^���T#�}�lb��t��7���=���A�=R�>�G�Q0��y&�)��Z��ua��|�`�g���Y��Q����2Lƭe2�>���W8&���5��SfB��c����n�韡�Ͻ�@�%��E�p�<âa@�D��k3p�0m��e:q|���o������VM��֪_�;�Mk���b ֶ��a".H^��(t�������7޾&�O�Í ��&�K����"�ᗉD��8��3�RR$���g���}x�4RPȇ��ЃM�돭P��U2���g�^�F ���a��<��������_�����o
Yi�`U�	��-�`� �z	l��{cV��$���ܧ�����pe�׹�Ɓ��:K���(h>�lW��:3T���	*foy+S�x�_�3}�ۗ��1���{P�՞G1֧K�M�!�2=��tky7={�Cb�̲�R]���� )�_�&&Yq���gF����\��;\ 8�����i��qu�f�_&-���6=aޔ�U����^�W6{�f�
�(c]̞��d���$F����f�:4�U�?<w�����:��/���퇷�U�-8Q�}ݾn_������  ��]�x���������>U��`2�KV�J͊"���3�%�1�5���Ɍ����ڥ_|�~��Osõv��TE�	n>U��,��d�1[��K�L�w~�ҫn�N{�8��l�G��!���3����7l�K�.�l�a������i��B��\�e��q�ѐ���eJ��݁�s�4�u�����k���`E�������&Nl�����Pܠ�8ժ!���SXή�҇3j�R�$��qї W��w|���UJ�3��,̽��:A)$(�<CI��g7���#2�̝-���)2<M{
3�1�6���Yt`�3�(��T=���N 5��[ Fn��ܛ��h/Q+1i{�`z�:%:�ϱ9�o�H'M�I l�A�
��Ar_���� ��grO�:Z4��$��ȳ潜A�%��t��j��`����{>[vw�Yuν��6�nt�7�&@���I� 	R"%Q3dH�����~�؍�u�������i��̌EJ"EQ$E'� 	�h�ܽ�Tm��e�y��|�~�K6�;�LV�_f�ӕ{^��$����Y�1��x.��WݲhI�H�P� �~�T�À�|NC�A�4����~E\����M��i�k���f�MɅ�m��i�A�B��?	�Nh��"��]��W��4����q2���I�;+|��d�0;�h��F��G:�K����(ԷL���;o�ׂ��[�!���[l�U��ɖ�Юm��m|�7m��-�����ǵ����lh
�� ���PsF����~nl<�J�A[�G.1�<s���+��gcH��:�~��*3+�%[EoB �r�pL+�o�/�#`��Za�+����Y��k��s���� ��L�wE��(R���o�����̱>H�����I�O �)��u� .��J�R�S��&.-9Rf4[���XeoC�Uق�]�	�yG0��;��f��=K���GdQ��4�s��1JW�l�V���o�o�
褥Щ~��/��V�7�=�CE�=���H��?�7��)��]DG/��^~�]Z�e!�Q�����r�|�v��H(�,?K��s���<������%���wY�R T�P�u�d�>[LV�ΗLG�ԫ{��k�?��oU��:�|9`�K��q����ߠ����bN,%�k��t�^� �4+�$����ƫ���(42+�-��G�-W���e+���z�1���y�̱W�2�gO��~�}ÍG�Di��Av������ޤ=��O���ŏѯ��oR�gɔg>�c�����{{������\9�3������Gǯ?&�"�s�
83�@�@!�@�F!*w09Ykg�������2]-H�V}w1���o��~���+'$[p\.ř<�I* �w�`:�l��${�����L�O=�H�'��O��%(��ܘ��Jyo�q�{�.if���rc���mN�
f���h�<C~��W��E	+,7���\֞�<�k���Fy�;�we޴Xp`�����e~��i�`�E�J����i�������.p�,"���Ȋ�c+�r���~f��U�+W�k�����,*Ԫ𕭢�P��ȫb@d3���y�?,93���n6ғO>H��0(q�:t����w��nY���d� �n�Nd�ڜ���9{O_ѫI�E�Q��_x�����7�	�=�C�L�d��76��78��+��d�r��}둞|��W8퀋�KVp� j�~9�:�g5V�'C�"�J亲I��	Ж���`.忹q���Ƚ�O���i�+@{Yx�fR�ǁ�2��I�T�����o�w��sŔ{��x5�a�B_�٪zh����Pf�؋�3�Y"�89��W�A�#�����+�J����������W���V4,˥�5�ʾ�5�#�J�����{a#��\*7<����P��.UKRL��ʯ�՛��Rh�>�v[���`Ҹ�B�+Qh��H�>0lEZ���L_�wߔV8 �sE��K�h?A�A�(�2��YG����!�+��7M͕���t1�v��(��*�$�m��wU!t/z�B�����ُ?B��o�������q�J�|7�q���ghF��J�p%2���-J~�[��e�
[� {��\Or�$hd��״���[�]6��^h�*�z���@�`�оHG/�O/��Y�W8K��;è�'�ʑ��4��T�n�)���`������@�x�q)#ߛ�J�1!�_���oe7�?���SLG��=��,A���0��K�;�LO<~����"�׺r��)ҙ���<_ZѠ�,ws��	+A��+��׼�J�Ѓw��l��l� ��!M��2L�oil��h��>�_ꖲ��g��H\����=w_O������rgS*�4�	P�d�I�|���TY]����r��.Ϲ�p�P-?P�/�-����:�1�U�2�R����3��/��d4pM��9.�������O~���VN�by%��Dk�>.�{Y��g�NXr�����3�YX�G����cZ9�*L�\]��Ԇf�9�z� ���i=���G� ��H�G�D��^EM��?|?������o��3d�`�sBk�l6?nQ���r�|�ӱ+/��ｽ\'u����*�-�rc��1��D�^�s�r>1`}Zb�#\�a��Ԟe�����k`��}OD�����~/��d�[�0��ʻNE����w������h����j;�׃+�r�&f;GЏ��v��N���V���]eh��yg���Z�h#([��b}�+w�{gg�>�����@����2��&ɤ�3S�S~�ꙐZ!Ncْl��e:�ܷ�8��+?8|��_P�<Y�q�?�?�?�?�>?m @<u���;�}}�{Va�'��'��9�Yc�2[)3l�QA�"���S"x��i��p٠�f���P����-��td}F[� �sΥ����`��!X5@Mm��`\5�V"���ʹN�,� k9���^��ܷ� ՚]A"<N���}�^���3qz�Q�D����u��d�5``p���J�����=��k��*X�ϬϧjX��K�6qw�GՌ�M���f���俪��$�����fҠ�~hv���߽�T����M�5!ȕ�~6T:���%r=�1��u�X�5�v�88��5�3��M���+�ܕ�۵��WdL�3oZ0?�خ��om#�"�17�Ǽ+�F�Ab�+>hm �N6g81�JGv%��ϳ�Yz&�c%��)�7�	A�f�pR���Y�����A�Hy���#ﯜ�&�8�'o�g�R3$mN�f�k�^���>���$��x`��X�@"�Z���g�=aʯ�F��zH��!h�{?���8KsǦUȠ�Wpo��y� ���H+�<���*��f ����XC�z&�zL��"�җ}��5���	����+r�jx�tk��&��3��yx�(I�F@�Z���is��:PI_�?c؛�G��8u��y�߫Lh��K:��3��]��w��2V���y���ř! �MO0���uT!ڸYlerՉ�����>�{�1T�q��&K����eY���Vi��F��8�җ�^A�k�����z���]� �h=����Zł��y�ӆ��u���B	Ai��j�;�s=��H��=�0�/_��8լ���d}h*�;*�~dr��a���v�w��֪˹�+u=�o��0�f��ٖ�x	1��ݤO�1�����s�����!�>���)y�HvZr d�ƽ���y�w�����<vG��ƤY���"S�6�@>�}퀈*hUe��m�-�QYA�,S��6�G?H����e�N����2��?�&��A��C�r�Q�ȗd� p��g�ާ��>�6K0���.]8(���� �s���}��O���� Y ^��e��<ϭ/��I���/������ʸW�A����9G�d�r!o��sc�Z��{F��"]v�z��<W4g9!���f>��G4�����`eWk�R����3�]#���Z�������G��/�N��2�9�en;�΄�B�<$I#�7���o��y�#�Ǟy�.�h���"'A��@�V��O�Ǩ�m:��rmXOS���b{;"xg�t�˳�2� �񛮿���:���~_�F{��%S��8�Bgs9��d��)��L��A}�ł�}W_D�<}/�qG�&��gܪΦg/;/hA��J�rdI���[�|�ڑ��[���u9����Ӱ
�������%�lm�&��Qۊhy�Nh�����i�`^t�X�t������^Q�-���6;��G�-8i�b���!�Y�>�|��U:إ{�5_�v{W���vP3o�Ŷ���g����/���)�b��`"�j�L֬�.�\��gν�����{�,|��[m"pՑЛ9��ٞ'�=�`�e���0���{�W����~/A�뮹���:���~@L�iɥ��-�g�Zf��Ζ�m�u[�����Ey���]J=rIݎ,+{t@mɊ3��6�=W�7����<���N*��0�Od`3k}%g���s���O}�~����0et�"5WC��(��*��ۻ6�(|e�;�J1�:9{w�q}�����6ɺ�kp' D�ɫ|F��D#�U���m������IuR��Ҏȣ��~���ч�y����Hݠٓ���f�c�D�eJ��(qԸ��]��hϲ��3_�Y�5%2*O}?�UPb��Sp�c�m�Q2�#�{6�R�À-)@�C&���k�G?z����Y]�7p��у�󬲓��ϕ}YJp���_X��k/�G�@Æ&/�gpk���.Z�d>�,����JV��;g���0J��3IPY�Z�ee�en���?���~�_���� 2g�B��VB�y)�^��+k��J���gp����ct��^Ɏ�nT�x�����a��U`)�����u[�����}��<����������^�o}�%i{�̬�$:��D�,��|�e�v�o��]���Y�-k�3���>z�#����UX�'��i����'�CiiO��h��D�t�	���Ⱦ�ɂ�\iI��@�~�z��S��o��^�*���kW9�o��sY�
s���窯�y���)t�Ek��� 蔙�@;
����-�Z�&��S?xK�p#�(AC�!+�]�V��e��g?�A����s�IRQb�W�`���LҲnÕ����
f�@�y��{E��(��Eߔ��/���N@��b��-����i��(��t4ЮP���3�������Җ�<����o~�{��+��N���3������/X��*߹�Ԋ�,�� �yG��v���/�:ʛ�mP�-�	��U�x�� l��jvZu=�	4��_� [�U��T_^Y�%W�O�ֺ�&[�xB6�DmZ��N]����Щ|���
�|߾rVҖmQ���JA0�@C����7�ζ�p�a<�'7-S�g󗹾Q�7c}�iJT�Qhg��z�k˸�{����)ze_'�.��(����-�1�mA�ze݇j��gݿ,�̢g�ozׅq-�<��b�A�[��5q�s�s�s��~~� ���_}ŕk�����-3�w���W��O�����Ӳ-��^4��v�(K����Ns�¢�3����8DǏ��j�"+�a�E���Hh��@��9k�O��F�l� �K���Ll���OT�E0l�#�p���+���n,ja��1I�<V9+*�.M��G3A!����`B8z� 5��?�
@��"�-+�d�9��Y�f�#���iv����[��u�m9�i Ѓ=�����k"t�(2���p�@-�Z��`�iǻ�v�έ#9N�L�	^-Լ�&��A�\����*����l�a�Ó���]��5����@3A�q%��.8�Ŧ�j27߷k�����X#=��W�A�2���N���ڵ�R�p�Uݾ1�Z-OO�w�t=< ��JbI;mG�Aj��u���:�d]��5ch�ѯ��W�d��wco�s BB;�a{*g��V��T��A#��_� P���m=]��W�#��|M=a]����!Zzk��u(�?d��YזNC�n�� ��n)�z0s����W/@�y_�����Ÿ�nT����5���Q�,4��h�o|ڳŽ_[���u�:-�����΂:����	]u2�ОN�����l�Uq�m{�{����hh�je�S=��Ά���jh���F��дH���^ D偐���R���Fd/`�H����"�\�jo�uϒe������6>�����u�x;�lDx{����*G�Sŉ�ox0�o+) sLL@X�ҿ<��P���P��p�uT���2`��d}u��qw��V�s\�#[�ѼL�T>�aap�� l*-XcH��<s0Tޅqj��efgu���		��T���������~��9���{t���p�1Њ������I�+vxŹ<sa���9=��W�H�u��5KL�WS�|ү�#�g�M ±C3q��>���U4��3���~��q�:�x�l��/}�[DkV\VwE�!Ke�`e�~�݁�6��������}�$�n�&%��4��J���t�?��Ti+�-s�^���+��,��D���:Cޢ?tml��������<�jV�n��$#����%��m� ��>z���O>A{�D��dY�Y�uV�BK���6Y���>=;�DU�	�˙�V����u�7�K���#����ik+IM�娕��f�1m���Y/��ݼ����'�z�����X�JP����?ZU8��2@�.��BG���T����;�q@��%	�<.k��r���d�'�[��կ=g%ʃd~ru��r^;�l���gұ|��{���K�ُ}(�t����Pm� ���r�c��_�3�ub��J+���X�j�ߠc�T6~�Y��Ӛ��b
��������Y^��a.�����e��N���rN��|%=���y6Ke�]�Q��)����&#�`B��.@�39*_��r�I����P� �tX����o?V�]��������T�<�a�9)�����d���=k9���5egn5&["D����=���ij���lMȍɀ�=�|�����d8zU����wY�$К�Eٻ(��[cr�̏1vAh3���"=z�>��e߂ �,cX�/-���I���̪(S�&�h��*o���C��T��k�d�w�X�]0�_��O���~Wt���G90�ً���R��邴���˿2��n�6?��İn�n#X,���ʯ�y�"��7I*>@'�}�\�c:��RݍmN,��
͌
��Y�)������?�Qz�W��o�B9n�?Z�4��U��2@*K�.rt���ut��W>�]��^�蠬ʝD�����&g:҄g�d\��{ɢt�砓`w'D����PC�ӟz��]��~�4�洌+�1� �;�2(���
�1̴�M��)2�Q�X��~��k>�r�;�H�s� s
��iU�h�؉�)Mdf�O��s(:,����r<K���G���?��O�.����6W��p��1�XX��ʾ}�G��]\��(%��l�JV2Ј����v˦�C�9'*g��I�ԞT�L�]�<K���g����O*!r��bAˢ[~��G���E��7��1EWa
[�L�<�$�q��X�d�w�����<F����G=�w�`�d�j�*#V��F���ѫ�������X��� Xe_�Tk����B�WJ=�~�矦^��W�)��ȃeٳ��.���ߥ�� 1��m`>�7��ѣ���E����}��a�M�떲W�˦t§`&��\�$C<��%�e�=�u"�����v�-���?|�o<�d�,�t'�/<f�RD̍��=녽��8th}���=ܣ�� ��41���7*���h�;�sk�����
�U^�ܷ�wԀr4?��urщG��'����_��tB���荼�|�F���4U��1_)���{���"۹J��]ec��c��f����DT)��L�f�3?�6ub�4���+�I!Շ��gc��������}]f�3�&�A:x�6)(ȥ<�d�Ŷx���s�×I�8�*è<i�l�6p�3ܙ���ߵ�y;�֯#� ���|@�����>���Z9��������ʰA�V���^m��qz�X���j(T�m��ySB�c�g���Ҭ��c,�� �������6  ð��k6�9p��[�}v{��%h�WJ~�j��:;�/�0V�>�{�}�U�D�G:Ǩ��s�X��W_�>�r��t�b͘c�ړ���X�/7�����pS!Ӹ��2w8�T�'����!c���ZX�7�~�~�sV�SJ�(VF;uĊ��b�u� N�T���P��T��x�Ԯ�B�`hמh��`�
s�ʅ;3-��*l��$@.�S�g��=ށ9x�l��6��w��	O�5@��2ù���Jx�D҂v�V��S�m�s�|��XSj�f���m*b�ɀ�=c�#�E�gO��w���f߇&ӿ��;X_���'
h�������Ю���=�G���h�],��s5�<�+j�5W��?\3�v?���vL�	\q{�y������C7	���w�Ú�5��������)TpK;���l� a������q�88�۠4��s4���oֲY�ݕ9�~�I&x�m�k�N�fͦ�me��L��]p��Qlk�Q3�����4G�n�g�u�PP�L�,ӿ�]��8& B���w�a��,�1&�@�������x�fd'���v�g`H��+:d�B5�l~s��A����L%�sc�SK�BB͘��,�76��7z��at���I��<3Ʋ�$C%2?j��w#\�1Md��6��@��슞�^ǘm��u�;1�ЌWK�ւ־G8;��Җ����4��:��!�Nc�qo�A(R?8���-	�d��@4�v��^��������2yE��4ň�E�q��տE�]�A� Gdl���I�*�Q��"8=��V�J�]����ޝ�|�w�i��9u�-�W~��_����������%��1ȯ�����"Z��8���}��J�{Ky֒����`Oʀ4�t��	���R'����Ќч:zLϚ��Q�K���4(ݗ9����c���-�/����͎��n�,ӳ��.�,p��<���}����j�u+B����m����!����Ӯs�T�Tg��ez�4?����
q^�r�w��o.U V�=��$;�k��.�Ӓ��d�rP���r���1gwS�[o���z�ai��m�P�Y���d�hA�z��|��i�0௨"��T�#ȗ&���s�1\u����_|�~�w��N�{F�^�!
Є/� �f�q5:�H����{�n��*�eWAP&���!�Vv)�ֲea:eVF�q_����G2����z)!�y����cO=J�������֒R?������V+`��:�	.�r��c���s�Y�uk{��6�7�Jm�U���b<c�nJ�Nt�`'P��.!*k�{�G[7�T��������g�op0��3�b��j�U���,!H_hs�6/|�.���'n����V>(q,������	gd	�d�����������.c��ڴQ)Ʈ������ʎ�%����a���/|�+t.�Ø����=�Mo�)r���˾���z����B�<�.τ���r�.�x��u�F�=��dg�/�Vw�;�n�d���`g3�<I�T�����C�t�����|�<|.��lc�U���sp��Ǯ��>��c���|��]�Xee�^$�d��a+O~�C�Ɖ��#Gc��3f����qK�Bu��Ç"�������WJ������q0��Vv�U_�wZJ}1����7�t��U'@��E��q��U���=����F&�r�u������_e�h�%5�T8�ynOQ���K��?�>=��g���������Ң
I{���v��X6�_�[?t+]��K�l�%��B{��+�x���H�u��t�X�HR��t�5@Z�q�
�`�T� �(<�+��y�r8I����i߾5���|S�#��6�%��Q�r!�˙T�t�=7����\��<*�!UG�T���O�m�)-��
����u��	 S�@d�E*z�Ǣ;d��)�&:Ē��>��>J��_�^|� ���8(��=����=E_���+�*�J\Ѽ��/Qۊ�q�A� ;)WVo�M�� -����O�t�}��j4.�=�Zt�w��g�$�W�z�w_*2o�U_�|L�60/�M�rj���e}�9v%��'/�?W�Su��*ť���u�a����נ�7�/ƚ���q+f)�Ќ�br�ژ��,���s~�s����?���93����
�� ����rY��,Ӈ����2��T��y�xY��b��ٛ��:fc��LӶ�D�-
�A�{�V�uֽy�Xx�L����<��=�{��}��-트���i�nUƴ�08�{��K�������)��=�� ������̳�]^��3�)8��.���
�=X�4֫�rI�U{�v�����|�����
mf�Cy���J+2_[@fG_qH@E{�$�j����BU/c� �7�ۘn��N���O>�oغ��K�zS{��lG�kІ�K1�с�6v����`�Pf.z�q?��c���
�|y<K��ء��^D�,���!�� 1���>�O��6C�5U��ﵢd�vy���*>�C��vb�2���,��9]�ߏN��o��S���V�Ы��	A�A��f�AqPB��ʕ�K2��</�Z�^,��G>U������������?��i ���wh�6~�c�;}꟞=s��o�R�M}���8���D4P��ղ��;)����1s�!�o��xa蛑�:�t�[�˯���^�G���0�7j��;J�
Ռ(xF@=+�i�j¦ eW8��\���?�x�~�^Qm�����������򽾅����Z�W�2q�%C����mZ\ǔ��i`0�l�����&�6�d�n?��D4��X�ϸN�Ci��k�!�7�FF�#�48����	��6`g!�#FV���}Uyl2�͙36-v��uf���v~Gㆨ�����C;���B��j�Ub =ڹ��v��hd�[�*4�q@;n�P5�U߃�c\ P��Li	���D�˾�-mL�b�3�<9����E��V!ŧ=-PC�O^� k�y�c��z�4��_��Ax(��w8j�2��S��x�~��2cU��i��l��|+��°���b�6��	-TG�WIpikK@�����t���5�f���0�i���i�2�:�����e�C%s'��^���!ٙ���um��݂[�e�32?����J�(wl{�%ˠ�抝a1�s�4y�qD�1���{&c�FK�����x��f«�y�#<X�ͮmAu�7o�Ҵ:�L�!���Lu���E�UH�<Vm�o1��:�
f����Mv��Ң�F�~dTx�� �d��5�����)ߏ��l��Uh�&�ݑ����<�:�4��}=�&��ksKr�Z��¹��I���su�ա�@��C�r��v�@Au�d.������-��W��:�F�8+� ����s/9;y�N��h ��U�!�����	4��$�3�ڙ�R���EՐ]��}�&mw ӄr�%��c��F�s)8G�5��\�~������W��_�ŷ��ghkc[{���֠�=�]~�!z���������hi�|�{��ڍ.��Oemc�{��/5�T�W�Q\�@�314J��d�}V���;)���8�E�Ӓ��F���c����֛������G���|��<.��=���ti�'�)��� )��(�T��a�u���,�z�݁���ᴊՙ��+b��vRE�J�_��� �n����C����/�-�x��os��>�_����ft����L�\u�,�&�bg�2Uy�!�0\�}.s�:��B��O#�����oH
f���(����u�.9����_���?�*=���i�ܦ�hUy`vC�~}}F�_z��|�Aڿ^�f�m��A\rpQ-�+�@4����E�Fn`F�O�K�B��M��ѤwB�o�C:	;��GF�U:A��s�n��j����^}�$�>}Ni3qi�5�����������+�u<C�~�d���A��!�To hW�����6_�,0Q��(�����X0ل~0��(m�=W)��/�����'���5��7\��i9�D�Tt���'�#�]�+��,�a���\�O@��.0�`-��Y���x������Г:fd��f��D(3 �j���J��{z.�iV���]n�����r�^x�p��Z1�j7�)f=<x�n��rz��;�tw�/v�N�2��[;(�`Ȯ��)��SWm�U��_�<Un
_��j�%Tr@�+ H��|Ay�M����������������R�?8�:�%Wh�Ce~�̍t��7���F�)�2�Q3qe�U��i5 �Ɛz*@Xi�rK2_t.�%���"Ac�h����1Fח��˞ۉ�w/ѯ����o����+�wt���0J�g�A�<HV6����Rz���|���e�"�l�@)�+@߱,�qt���`����5Y�.�����6�����L�Ȟ�\��.�� -�\��?�������׿��[LU��+g��j�c�`��(��8m�2�nѯk��OxS6:۞��0���XuA���O�2��I�� A�+p��(Q�i+)s��>A���E�_I�'_���z��8ݺ��8A��G�\v�������+�tN���a�c�]�9�>o�@����1�w	�\�Ҧm�7T�.�����8�Ng��0]c%�>�G�GϿL��ߡw�=E;;e~�:�$��e���;v=���h�x^d^�V	!(��FՇ&Q!4�`������e�<�Hs��$D��Γ���&N�=9�,+���{o��7������+z��wigk[���=�U�`���}w�B��w���9Z[7�s�V�]u� �[�����Yax���`D��q�rU�@(/g���"U�̕`�$�07�s��_�}�;��_}��6OҰ3�ub�0m��V���B�OH@ }ٿ>jKHt��Y���v3M�#&�[�B�y~���Cfg��S�o�3f�Vp�*��χ��y��t�uG�E�?���t�l�W��KƼ�S�DO���k�{�������U��S8߽)ԟ�2��fsUL�W���,��u
�6�}�~X1s����/�3������'��o�������o���-��M�/7��]��y�Mt���	m�Y�5K<��::�9M�Sf��|��������?�~Ya���6���ɕ���{C�-ʴw?��.ml�N�1��G�1W:���c�<�]υ-z��t,���\B�{;
py~�|��!�Ϣ�K�uMB�U���ʦ+�G��rͨk�U~�@VyΙb�Z��wަSE.q*�7n��(������i�HSg\6��kT툄
����ċ��ƕ�<�39�����'�hc}>?9Ù�b�
!��r�s�s�s�3���+ '�wk'/�wѷ��;��?��l��9eP�V_�~8pS&+�����/�77����CehP��*JX12�.m�_�>]�Gw\x]��C[���	e$��k�.gФB4E�:G�}wd��� �Y��߿5.����kg�l�N�� ���M	E��lξ`�87���ȂB��5�%O�*� ��������ŝ�pd#�6-� �?�{�~���⚯͵� ��%�'�`o�6m!P[
�c�S<h�8�=����{W�9�	 ���&c���ѐ��9O�.�Wa�'���<���5� ��
q��s��D�m�@?��4�2�j����r=��c����j�h�hJG'���'P�%~O�������Ch72u��E���h�ǙŶX3 ���l�:=Gg��.�����F�^�Rk�c�5����;>���.��d�Y��� %;��!�ǞтZڬ�c|ϚRp�X��:����G@�����}�����o��G�bc�危o��)�>���"��=����ۍ؀D  )�h��d:��[{�X�u�*&WQ�]{G}׀c��.T�m7�s�́ un��6�����AIY��,f�l�9���(�*�^���/�_W�D-oW���W Ie>���d>$4vLչ#?U���u��:��֬��T�kx?�G�o2j�@]��
�tc�JG��\s���=Z��i���z)\���nG�9~��ە��&3�c����L��y�]B���a���0�VOh+S`ͽ-@ ���{�d
�0����]�r?Ĩ;:(�T}�r�ٍhb�6�?tM�O���!�*���'�5ˤ�Ky�g�K��q6��+�/}�Q	z�>}��~�m�8}Z2��^q1�-z7g!����`�@��z��5���U���
��:�:�q�R�X�K3GU�q˲3'�8"{�����F:p �����n��^}�������$S��t��K��;o�����Aʔ2�����'��(��ʜz��(C�,���[�EN; .����3�F��p���Q�ڒ�o��+_��,�ݤ����}�r��|�]z��hks�콀�>B�^u9-˸W;;�����M�Px�j�	-]��,%9��ʘ�V9�T�ڭO���a�[{�jF�q������Q�����رCz�y�}����<M/�����I�)sY+�uű+��cW��l�؋�4��v�u;ĥb�=���Ȁ5�S�-�07�+GTB@����ͩR�~ ��7����
-�a�U��.2}�#��b�t٣S��hg�#���'���^�5� 庂�;�Z~��:JgψT9�Ò�w��;����x	d��N�s������&�]Vg��ν��<���.?��]����o��z�3b{�f3��k��{�a�.k�M�B��<'�������^�.�d�`~0�-h���~T�BU�j�Lk@I�P_�P�yɉ��|җ��yx��h��]��<�A�N��e[_�C�y������`��x5?~�A}7������)�.dgȫ6�\�7t�
�"m{˃��*rv���b��,�Rٗ:i��K:x�/|�1����~�~����ko�39D��z�� mnn��xZ�L�i��V��+�>(���`�1`�A��=�!ǐ�#�_�X�~D�c=.��2s!��
��w�t��K���� �^�uz����I�#�x�&���$��KǼе@�Y�q�3*��yҊ����-��ش�0=��<5{�-�u�1�`>s����>]t�b�=����77O���3_u�1��W�I/��-�u��e�.;H7�u8z�p�Q�ƌi��b�5.���(���$֬:��hӁ�/w�ᕡ�v;e�P@xl�7/2�}�:ͦ��Z3���������:��g)�l��|�-�я_�j#}�NǮ��n��F�*�mll) ���&���y�{�k��@�
�1�֝l����Xn*u��'������d��{�M�"Dd�ؗ;R���q�x,��E���<U�3���ޡ�_y�N����_�utɥ���F�϶�8�$9�[m+��!���L�?�2������`	75|zn��� &ɂW��𼙾�/빧p�_��Se?Vt����}���֛'���]pp?�{�]tY�97Ϟ#��b�wk���u�`<�U��F*o����̮�`Ȑ ��cJ�1π�>�Գ`�i%������>�1~�M�^{���A�����D�����ܙs�o�~�����G�[��Ut�ٌ���(��Ǌ��!Y�[3����`�`��Mm���D)�� P��EIڭC�^��\�̷��rfv�i����n+sy�Μ-v��'��"��\?�Vx����}��+�"0/�$j���a��u�%%4�s���j��rL�n���[I�0�t��p��������X���msZ+��Z���/���>]�ʞE�N�;o�C'�NƟ�E�-�&�Q���UD�����_�%R�^�}?��[&�R�`�X�a�=����xEp\ϬU�4�ѽ7�����Lm������Q�3�m��|i�3}%��x��rVϔs��~E/�|��;;���������r��J�V�*ì�q�lQ�T6ynr'6 �^�|�lQ��_l�k_�9G��:E���C��{�0�/) _��r6��(' ����<ن��mD6^$R�lю��|֋Mp�7�O�:�/��{w}Ϟ-"�����������'|~�  V��э�Ν����#^�����y˗_�굧h��%��cc@��*SL�O(�O�h�夜�(���bŕU!6R��^��^�iY��E�z�hoaԗ_p!ݸ� �[[�YҞ1�[.`LA��z���J�36�	J^q�N����}���׷���sg�bܞMK�P0
@!)��)���t�f	IYN�`D�P�0l�,pP҅|㻦�W	����<}��{U��͜k�e�ke���]UF�%���5gP3֤0�E�_�_W�0�(~�PUn�`�f�xVe�"�cԞ}cn���fj7h(<P�B44a��腡�Ҁ.����0F4{)k��v����7XF�������>�_d��I�6X��L�x5W��Em���1c?�{3u�a��>�ڷ8#���{�'�Op@D�EsmK�`� k�����Sژ�>譖�u�`P��^Zd�T>Xnj�k��d�=��Ӕ��q��w�!�U3�ă��X�A�v��k�������D�#���k�C��f;d��  衙���Un<�D}�g�X@����w~7R>�}Ahw`���wT�3^�V�'H]��#F4P��5��8厷v0�d����]������ f7-]�'3�N��ȃ��Զz��� �={�����sf��E�q��'a��Eo�>L�	�O�m��Q�q�5��2~�kdt��;9@n��RM����6���i�qg`Թ����A Xi*I�ր)>�D-o�8sll~��Zk�lv��[�Z���g f0Ch�o�$8�U���zƾ��qNx��j�� �r���5 E��Q2���G�s�H�4>2��6�	��j��g�8P���s��/�y�F)�7�0W�F����=���R��ЍR&�����Uܝ�T�I3�y�,uW�^���������ѥG�u����\������	"����Γ� YGΰg�������QFƗ��Z{����a��}�����Ϊ��stF��hOX)Y�����>c�jE�a�.<|=��}D._��� �Xv.��P9!Yײ�R��h��9K�� ��xg��1HUG�hp��	��Dz.ͽ���$ȥ��ei)YKA��:n"[�=������s`	��r��1\R����~ g7B��3d_Tb�(h�5Y�\oY�v?������U����`g� .�}��A4IV  tNv��`2��[^������C7�x-?�=�)[I�N�j����&���A�eG��dur�/&=Seo!$@$;k*��'_�3l�V��nbZ�,�=�K��݆��U������q2�f���L[綅��qNݢ���u����;Ҽ���
��2�h|"����b�QQ����9��h%��e��#7I�]j�W�j���,��U�1,h����x��%9p�3��;�k�t:;~)�ak�]t�>��c�e�`�����S�W<?U���y@�R�G�iGV��fZ���9�>k&j����~�٘��߯��k�Q(|��fl��N&ބ�G�G�+/��D�*�9����r�V�[��$W��DW0��X%�#A�B���_JT3P.��<ɼ����-��&�^F�-Y�,d"=�H���w�Q}>j)�IU� �l�}/�y�-n�U�T�N��o��sX�ׅoh�s��A�H�7� C�/=��*���S��@w��H��!���'%�HE$��Q��V���NS��'E����~:|�6�2�A���6ϔu�3mj��·�:�C"��8�C-�jp���N�ܳf��}�Q�{���3]�2dm=�ʱѡ�frT.�a����u[�VX\8�w>~7�?�������x-�y���0�ZK�s����C9k���)�V��@¤}ܵ��tUv���l�l��\�j:p�1�x5
r�eo��e����?k�[-������t��뉮S�6g��>yBx���g6A�6dà�T������У������>pI��މ`��`��/陋�>g�����K���J���(v C�
��윥ͭ$g��+�����Z���o�=-�
h ����%������RÁ�~U�0����\u�OdvF�G��xރU�OZ9�̃���t� ��N�]��ADrf5�����i,�ϊLY_��λ�KE*_�r�rc[ΞP�X}F�OB���,��g�q���ժ�hv�JE�A fɫ�E����zzO�3�/���5\����5�S��9�i� @�J厝���}�?s��=2gy���������H���i���`�3����=��TiR}�`ZMIu9ҖP�ߖai(|3��F��+�TJR��/����u��	y��#ʿC��tV[;�g���KE�$�5�Z@W�+"Af�*�Wd Xk�a㚟"�R`��t�!���gOwJA��Yf|�)Y�^���@(��G��幝�?��������9���m;��p�ު�Ф�>l�0S��f��5`���)�����#�EK��)�GTAR՟e��$��S����k��'V����t>��P��'�>B4"�8���f��9�G�ݯ��Jts�0}>[t5��-��s���\GG�{蒵�t�l���5��S���p���ӂ��hS*k�r��Q0-��d��h`���Co/7��q�N�1m�է%v��2[��g�r��V��M�������}��l����膢'�psߡ^	}~��Ɠ咭��8�9�9�9�y��]�?9)b�Č� ���si��Gٕ�����S�qu~ۯ뷹fk� Z����$e�+IQ��mv��]�:w�Mz�7hOQn/Z�#�@=8_������#�<��I�x@�eq�@�ejU�p�(�'6NӉ�zg�C�`��)�"�O3 �Y��~T�X'����`�ٌ�a� +��\����	�K�\���h%��!�q�
��c��%�~5p��Up26��9�=x�k��L���]���<c5L�C��:��J�8�,�#Jg+ՠ�z5�����Mk/�`j��N�ZJʑ|T�v.ԻWR�6TU F�1���ᥩ�=]�mZ�{�+��~�}J*�Ÿ��
:3���L���k2��B��~C�����iV[��O�{�����`����5���Kb_c�,�6���4�{�y�U�3!ױs����K����c-��l�_�4�����pFf8���4||T:B 4{
�#c���c�N@~a�{�����CC���gs ?�e�|>/���+d��5�Z3�����j�@�:ǚY��'���`�ь|
����9۵t�g��S�PP�.C�G�/IV�p�)��Ι�=�)�5���w2�6����	>m������u`!����]PѮ1b���}p�+`���Q^/!o�'�ʻ�|�O�s���Y[���*H���#��Z�-	�N�*�v��D}�(�g����� ��\����R/�8}olm�`<²�4��tŋTKz�>���O��   G����R����EgV=oA������et�q�m���ʂJ\��T9���zv���ߡl ��x�Z�� }uH�`�����k�%.+_�� ��K������x5^�;8x	p�խВΡ���m��W0^}_Osu(�9i�ShĲo��58��.�
���:�%cOZiq�2�1&� �.̍���d�g+�im�P�S��({|6G�������%;l6�vP�����kp�e2'�`�����T^�<���ᝡ���܅o��Ft���8��>�iA�;m�Y4�lM��Lu�I)T�9��^�H�8�Ot��U2���U/�]7d�*�HC��x��yN�Ks��2j�ިR)M�Ѕ��������<a�����-�u�d��^H$�#���=�/._7�ڍf���{�|D�bU�4�3��o#W�Ӡ�Wz�26LR�7@�(�P��,��9/]��b4�z���h��ded����n��l��,�F=��'������j0\��s�=�!�^2\%�_�d���b7S0��N��[���^�V�҂�����Ԓ\�������Zɳ�U�*����V?�N�m��c}�GȾ0�f�RD��l��O�1��u}o<�lB6A����  z����!�B�������Q�.�5���z-��%+U��]+���5A��3��S
��^Z-�&KF�|�c�zT���(ۓ4p[��g%�/�3�.$�Wf2LF��jmFr=wdv�hA�`%�e�2 &Q�Z"���T��)Ƌ�J��r�Ƭg(�Я:�N�{Mե/�[-%Ӊ�_�����;�h� Ylt��@^��`���i�Pt��j��B�@F2�������()e��lэ�y��eM�Lb����# ԅ1�*������G�%�S� �A`.�����BߥF'�Nx��x��0��͇��MRT�܏" �)3�-�eMF3��>��+B�
������1O�*m�8�Ϡ"�=!��̟�tϐ�
�\[^m[�I��h��Y�bT5S^�4ݛ��v�6_�@W	�6I���<�8����9e&��I�>�+[�$@�1hE�eX�YA�1�%hͪ��"Gt�hp�r^φ�j�y=լ��@��"���.M�n]O9�%��t^�G�O�����T��̞3�����zpl9�?�'�AB���T /e/I�R�3��e|#�k��W?}�%y�kb[,t�N�N��Au8��/	u�(S 4���~�gK8?-M�4�l���~�ڏ���M�|�N���-�J�`�D��й��f$���2C0Y5�`��(f ,�#��h��J+ �X8J��l+[��|v����]uQI�IYO��I�7�̅ު:�`�c��t9�� �x�9����;���Z7�J���$e{k�0�d�B�+X��Aز�u��T�o�����,g��m��U�j�z6��������?�8�i#�������3C����h�����z��Y�Wh�P�F�5�����KX�7j�3Yq{�����e�-iE�eL�W�tj�Cg��{��};(�GZ�1�mg#�fe݇�t�|���3c���_(��'���=�J���nn��*������������?��� @���^�*���K������vT]�ГPX�;J���h8�ܔ܆ �*�;L�X�!�QUtDud�$�mf�E;ڜE:]�vj<G/�٠yQR�;�)�b�lA�"�1<c�!�V؏E eyk\��r���D�*J�Na�˙8�A��݉�Ov����o�B海���0Ǽ!s� (����re�d��t��x�u���ll�@@C���!Pe�Z���с
���]N�{!��O� ���xYX��Z�s����b��䀀L�
�@}�������~�휒�Ֆ ������`���Wm�{�����߼1E��>���'��:l��t\1EP�5�D��F9)%���z�ܠ��f�xx(���X�e��6�]�6سa(z���kK}l�5��kpv7�!Ц4�h�-GU�'��U�3覥G�WP�i[� �טӄ�Q=����3rmE*�`�m�^��d6�ɞ��f�{�+�Y-JMH���9;`k��V�/��A��ʱ�:�k��TaA�d�U�#��\����,gd��*���dN5�ʃ6�]��=��7-[�����2�lQǔ��~�����J�Ҍ_���g�g(W�0�� ��/�3�!�)���W���V��yni�.��n��ܐ6��kk,6�B=~n����2y�3�uI�\#��f���Ys�
���2�+ooiҜ2��I�������v��#��e��@.'��ڔ������xn�q�3Q��8C�[����}NN(J�'G�9�r2ø���P����1yw�Jt�ۗ�M�-{^4�o��}ڊGKR����WGBjD�Gː�� ���D�AU7���r={�zF��h-��K��U� �P*�"������Po�<L%�g�b�����8��Y��4A?����1a��k���j��F�;����%�2eg��10t��\��F�o���!�`m����γ�HF6hS�'�P�D�Ҧ	|z] ��D^'�f�S�=$��-X��xq���	T�N�*�X2@e�;�������9O���U�"��V�D�Ոu�cT�,� g�`��E���T��ٝ��7Ȥ[F���G�G-_ Tǫ�wג��6��7f��@���1 p�+-�e�}��e��fU���i���e~�fII�bDK�L�=7�k�~5*hժ�l��W8��G���I"̷K!�^=+s
ɲs�W�`�Vu3�@�3z&:�<���Q���UR���*)�]�Rth�Lq�m�NMߠ2������E��&�,�F��/cr�`���-]�}�� �]H \���6����z�Ь9hͿ�:�%���0{̲�c@��,1y��@+m�Z���i�5��ŚW`.�?�{\��y��=H�"����|k-����}Qϸ���qz�Q+��"�U[����*g��<�r�&�R�@��&��Wxa0�$}�!�&�|�:�����f3�*��n%���|��Zd�l�v���a��u��������K��a�Z��!�Nod� ~�,�*����l�	��d�J�3j�~G�1��>Am@��ٔR�`!]�t���I��b�x�k��cg�y}��O�ɶ�����h���ʂ&l� D[�_����-���&��Q+'C�	����n��f��*|����Px����D��/�x�����+�@+�%����\s}���	=R�R~n��l�V�A��J�N�Х�
�t�:��}��C=ō�ȓj�Jx�f���������� F�c�.�*Ph�F���.T��:�
��=�v����� ���s��4 Q���b���fD�蓂�/��uEˉjw����W��-/\v��#�߮C6�T:T���H�DU/0��\U��	`u�������5�h�x��`z� �_D�eϙ��_T�3��o��1:'�Q�����Y���f��.��{��
����{���5ݵ=)|���HU�k+е	+��U��G�w��-�w˵cjqy��5���ޛ-��j*�)���f'����@`o�߉ܠg�3�&�1lѼ�㽹�6�\I"��р���B8A�3���3�q8�3���Oe�C�I��3�G�X��q�h�4a]"��Ʋ1�(%�@��u�*zI7n��Zd���}Nm�����y��j���������������?��� �j�1��_�����o�����$�;�A�YQ#���jF�=@��P��t3G����8C�M�_�9Yy�,���!׷�9]t /Ό{.��ِ���e�.9k�}\2*�f/q�&.� ���P�>��e�K�y�	�vUR���he23��X*�j0�އ�)׿7����ￃ"2QF�+M�q�z����*ƭA�� ��m������0۽��E����r���i�nd#�N5(�Q�,�ێ=�r�`�����h�FS]z�=��ɞM��극����٣�`�U`:t�P�p���Vu���>bd�n{�5�
T�~_} V��To��a�@�4���1,P�eqg��q��Q.�'�Q��A���f��}0ڪU=�Ҟ�E	��n_�\icQ�͜�У�C�9�-(�+)��P��2@E�w ��g�Ih�L�P��'����� X+}���0z��y���v�Z�/u�w�����O�W�-TpT��3W�S��y��fCCc� � A����[�~�+�`p}?5�a,�|��{��9n��)�p�R�n|���g�#5`�����w5l,�RE{]�@-�����D�k���R���_ BI�K �߇��Sj�:����Nv6T�_�V�=7���T�Uu�ʅ����FM��(r0,�"hyWTD�yT�@5�:���ꟴ�u�8[~���3��:�4�qRyŗIq�h�wr�
��\��A����p1=�]m���2�g��47�P"˖E�3��� P:�������v j�Fќ�l0>��àC�4����ox���}&T^�
(�Ӓ�Z��.�?����Z��kQ�%|ל1�j����|�:
�q�\���4<���n�ɚ�s�IKe���9;�{��f)6g�-
4��IyKɜƅpVB)Kd���r����wp�	өՏ@��� ��aC��1���R� {(
�PA���`'!@�d��R�tF��M*F���C�{	�I/`�g(��v�<��X�"D�<Pf�$�^�	 ]s.������Q]/c�.W��K*H#!�Kn�9+�!�͵ �4����R��:��N��pz�.T�\�+R=c���&ɥ�N�\����(ٚ7�gZʅ�3zu4g��d ��
�����z�����#U*�w��p�Pu&��^v��%]'�*#�S�'�!VY
P$2��L�BC\R�n��a�΂,C�Zrl��C�'���.�*%&j;GAT�0	:�y��d�f��f�!��I�_zV��Z	&ٹ��7��kr3Z��2�^ᖽ	���`rRdc�LNF�W����Wz�܇�]������x�V*�yq�1�F4���� �<3-���C4^hA��͠�L�T���4�$��
x
����ݭmA깓/.4^*;[�_ZB� ֑�j	ZZ�x�w�D
	5���>���,�Ҡ3����� �j'���F�j��F.ϱ�i��� ��)He����Z���� `�� ��^��2�$�J`)ZP�.v�j~:TwD{# ��:c�y�$	\�)�N�:i:h��l��W��kL.�<n�!I��U�@��:ڞ�R����|��.M濑�#�,�p��IZ����-hC�@�����N��y&z��1" �J�`*����zB�Yڔ ��=gsЭ�*��[��<9��T��ߒ�r������@���e���!�8�>95�u��jk1����~*�e����VI���?ic�L��d��(�U+_*W���T����M���ث������7� %,��`+�i�9�(U�B��`;c�t�@�t�I�g��4I��M�o�Y��7=䖓��g|L���FB� v`��DC?���V��}������P�D�$KP
jsD�Q},��	<�;%�%�C����Ġ���
�>��WJ�����U���j�ڵB�u20,묒=!�+�?�&� �W�~v���=3��f���:����PETۊi� +`j����g���4o� E6	Ң�ϣ�j��=�����-�!wU�^��Shv����S�WۆyF�kB���`��9;d��Y�H-7�=��� �9;0�s�Y���<ʯ����4���'t����?X`��u:�D���
�Em�:"0,��M��l �:Z	����?��߿��[�x����˅���?�?�?�??��Ӯ ����i���[������M纝�9�^*:u��o:���D���N�����5i�U���2�e� ��Au��b����Sc@����;r�(���q�,
|W��m�&M ���	�#��m����#&k�M�IC��C�{���16$3��
W|����F���^w#��E=�@,#��+��ϑŅ��a���<���z�g���~�h�&��7�4���$:�d������]����"�ͤpZC��왥���� n���^(?�$�@������� .�mC� �����8��PB߾�"����k�o;n�f4����N6�f4�w�/�rc�N����ag�ȒT��HTI�8�da(4���j�`���ʩ�^�G��z)ِ��VsgB��u�sH�j�z��J6Wɮ��kَ%h�!p>[��8�U�4��0xa�!�P��p:Z�P��M�zF���䥷����Eg_A7�<&���G�c]��4|����E�I��f�,�ϒ�����9�H'oRC0�_0Z�=�%0�&|��O�~A3M�Ɏh慒�X;]�P���Y��p0�ct����x�+H2���sc{ !���p��N����S�伥�sBSνzXW�-�F��51u�c�l�Z��.�<.s�|�9�*$����gZ^_i%���~cc�$��}�	Zޮ�[[wd%uƁ��T~	>�9���TL�1
mw����]Fƒ��lY�R
6��4������o�:�T�y��0�E*@w�G�٤\y�U>PR6'���y��%N�46���^Ø��1�B���$Ъ� �|�����G���0��P�@�~5�+�F�:�OLM;�Nr��o�i�l��[��<�
J*[�E���Q'΢�1ݠ� �h��,�<D�����12�H+q؊tq�\�k�@�mV#[���%�r���b��W��),�`\J��y�~�{���4�f���@�e ��6��.�<g{�9�% �k�[�^� �@�s��25�	�[��#�!P�j!���k��4���F�u��͔����es�+������QʜK5�3��2 �OpBnրyWY��=ñY���?wP�K����,�U��T�~�?��� a�	�����m�z_t�٬ײ����e�У��R�f �Y����#X�M*w��(A�
����ܫª���Z��We� �{8�	�@r;�����8S�ҩh�mu�|�8`6ڜ���?�޶ǒ�:;���VUwOwO�P��B�(�Ԓ"EK�]�^��À�������a��aY������!Ɇ��H�H�p���pfz^����8�yNd6����R�]�%{���V�̈��9���Սl��늚���X�vJ��.q�H������= 0�;�B(=��~�6��^3 }���+((�D'z�7Į�M�$}c�>��ZA��>��g.d��lZ�W�$kA�t ��fv�;c���w������p����ș��m�X��A}N���̀���~v��Cj���ϗ+�'k[�`�{�� b�0
A���s�u��Տp���^��nyl��;�W(a![���3�m+�+��F��u��q̼]哇U���#���u�z9 ��̝7�IZ����,�{��	crr�=����&L�������ػCS�=&r��m7X��Dlε��*�j�tP8Y}� ��h���>�X��)`޼���������vJEI�Ā��Ξ7���4c���4�e�#� ���}��\��L�A�����IYGy��()΢Q�&2s\"(�'�K���峪�Uz���քӞrܙ��9�����&�j��H+P��S���mP���bM��J�o %����.�CVt�� K*.q?��~?�g,0���ύ�D�N1��St��*ѭ����k8+�M���^��� .Wc��
�y#���Ч��*�Ы���$~n�x���70���t���U	Ġ������T����%�7��ʅ�"maf�� ��q���~^�%�y�p�+����.�yR��dԑ'��� FcA�A�ˁ�Զ�#����Ў��<\u��xN�4�b@"�b��KطJЄ�%�`��x���v�[�L{��r��d�~&=6����G�K���r�*���d��~ob��}���9��ĳ���E�Mp�3
ǨT�q�-�n���Ged��)���ƾk�C�D��v�����R�s�^��F�j�뾿�lC�߀�0��	�j��c#�́������}�b����x��V	p�s���ƶ�k�;��s�k�5��y�����,f7%dx!��@eRi�<�a�&-y�K��R���J���{a��dωd�2hT�=��wc%p���5�Rָ<W�^��HP��5G^PV-�˞�ެ�]+{���,;6�d�����ׯ���ߟz��?}����[�n��u�yݼ~��' x�t��?z��{��߻��{u��:簤��E&��ݕ>�z-�l�N����h(EH�H臲:�P�4>5�D��P� ��Ν~&��,����~�3`�H�1e�Нu/d��;zL�QpC�s3�Z��S���=Gn
N/��}����^�7n���p �n�}F�!�j�>�H6��lh�7�
�z�������?��F�e���#=:�#�N�����|�-}���.y�U�c	��ۿ�V�m;xl�����з%���^��#�B�Ʊ��_
.�^�]����� Ix����X���q~q�O	/�/����վY���0���"m����ٟ�g5�5u:���)�0w�)�^��u]��_���
�f����0"� Szbw��k/��J]�d����M�A�A��g���]��碾q*/{�y�]���3��������F|���z!G������z��|�3��u-H჊8�kO�l��.����[��z�W��܁����k��P��n�ڵ�=��EG�k� o�.c[}���^��ގ^q���  �����3�/\��V��w�I�|�X���{�9�~�hc�����+$�sYG�lee;���� ���NHXr]��8�:�U�t9���.�N��� k����l��' drG����"2 �n��>�{��ou�}O�T&�Y����g��L?[\낶�i��k� ����u�>#���)m�'���k ^�Z�.qM�8�͒e���We��u��@���S_���
��e|U�Uk��{�	1���������M|�h�]'�n�W �ˈ�������
�����z�R�+�~.����r����v�,�#E/��7���n�#��dW!���D�=�Z�)�ߟ������Q&��k�G�%@#��|WR$��Gy�� ��S����d��z����eLz�	�7�J�j3^Նi�M;���,����qU���H�1���#�q_ȟ&+�LZ!k��q4?����[�u�Mv]��މ�N�Tϝ�����x��W��`+3;S�!v1J֮�D6=I�X��2F�j]�u�~>�^n��ɒ�����$���"�v�s�N��J��9z
��)��A+R��R'�����e�8����59�%i�	�,#��;\*�®�4��#p�z��N���j��Y�$3��� (&�A:`»iQt�}]����Aa�X"��}[�d ��nx��]x����XC�-�|L�c<� �>hk��8���x��N4�L�&0�9h����&�p|<DbQ�`e/��G�L��w�d��1ۺ�(�㌺�b	���vDGT����E�R͡Y�K���޺�wZ�|�(v0qkE��`���/l���?C֤���^�������$�q�ϩZ!o�h��u�G���;�Pt�YKv���Q�+s�/q2�
���d�b1�XH���� k�%-z���"
PT��EE��>;<E��9�|�uU�N�h"�υ���� ��fA=��%��,��{����� ��%m�Zbl�"x�8���Տ�~]�P���w��:��y�S2�fő���h�m�/��f����>JP׏��ܠ���b&�8*���b�,��Gs��ܿ���QA4�����ף�nK1��Fk~�ʱ4���3���H��ҝ!��8�#\%Eʘ�M��>�r~~K�VcG �a^�ڞo�t��q/��ꦡ;On�p_q
IB�V	�2 �~��C�U
FV��wqߌ>+c�3���;Y�����*��;��Cf��v9b�A;�1&���%�iH�O�W|�M��W6�<�})�hi��E�(G�ET�%�����W_A���{��͎2��Dي�	{d���3���|pLi��r�S(������S�ȿ�lB	*���2W��=W���	�ǘՠ_��C�qgv��O���Љ�r<��`�.rP����s#� sv���q��R��˔Ԗ7���_;}2�G-�6AuW~�8����%�<F�5��������D���Sn��+��޴�\!F�$ߪ��3z�� V�����bv�JMmm"�A��u��B���|��5|ѯKZ���ct�'��3:cͧaD׽B��7�}�B�8=.�r_u0�^�q����&=�Y2�u�9�UX�����\�x7Z�ޮ[��f1�γY�NV��c(�e����]�?ɀTc��ǁ���Wz�Q�c�,d��}�܍q� R���u0���9>	Q�]�Z�� ��I�ɠ	vΆ�lcv[UCd�J�]���z����lR����Wd)�������:�yu�9�v��{���Q�Ry?��ExdD���j����g���bYG53/Yּ���o�9�]~2�/�a>��C��?��z��*�<�tvo*T�$o`t?��|����='!��~Uw�ؘ�m<��G�������/>u��y{ץ`"����u�y����8 `�����g����+���R���9.�ؑ�"�lJ�P Mv��u��?Az��n`a�aA);�͠(%��ь5Gf�A�o��Ka&	�YJG���+���s$�ϼ��=��������s������l�j�Y�#]ʹ��5���ؑ���w'��~���P�S6l~��%��u�"t�Zt\�x�ͽ�^���0��U���]�e-�].O�'�B�w�)���;Ko���s�Yd�E��;ܑ��P˺����!��va [�=�\��-p+ ���eA�މɮ�F����Я���4��<|a�;�V8fr���$��oՀ3�	�P$b^ј]vE����䅏@G�y��Tv�ǽ����T�}&�����NfOLv9���ғ(tԻ��vݲ���j��JA�B$����u����I`˂:�`�"�����tu�yPu-<� !\]�2�
�w4�� .�3����F�UA������s��#�7a�Z�tl��ǜ��2�$(Fnw�)��P��\���g�zR�T��u���_0���l;ǲ�
�U~�"��p�\�h�ȒxLn�z�� ΐ�e=�^*.|~��Ă��+�抳����y�<�Ё?0[^ȍ��(�W�e�	�@���U2�-���'@����Y3����`���׊vɒ���kz��%���=i&�ҟ��`p���B�)8��\6^F�}ٽh쀷M�(n!���M [Eք��+t���:���yGaOa�*l�Dfr����͹3*e-r��{����jN�ц����Ā �q��]�����~�	ڃ���K��aO�ۋN��A~kw��_[��AVog��IN���� �u�z@��c�rf��h����kZ��g~.~�rv�_�l�/ߏۋ��`�=�Mڮ	�v]��{K��[&���	��v7x"��}��������T�P�,Ie��u��u��vl=w�f�Hq-����R��.�<峬�Q�k�PwZ�VA���:D��[6	 �`�zH��� Kx2aiI#��_0��,g�nu]e�Mz��h	s�#�8j��B^�ya���Ve���r��@7s�ǡ�|ql��� �B����[�6f���~�&5Omo�룥�k�(@U�3	j������.]5�F7L�R�^�[�o\�(,?�n3-a��}&[��o7�j��x�I�d:n�b�!����U����Тd]P,^ڂ��lt�yӯ����&E'���	n/�:�3�U������y���9�6@�ʌ�g�x�lr�X�m*C���V�Be�Ҿ����eͮw�Ĺ�ќ�l����+Lj1G�0I�.�tԳ=�g����/{w���H�䲮o xl�3����ln�&�9wx��۞�H�>SC-�U$Mcr���y����ԧ��Mc{�C���8�l�9@7W-�X"�B߽ˎ��~�sV�gt[{r}�zC�ʧ���n`�����]��uI�����Q|J%�+akd�d/�8S�֙�X@����k	mc����{���� �f�L�;�[�Xח�����a��ZѠ��M�B�;u����)K:���39Z�6r|����̨/��#�C\V���Dvh�T��q�E�\0q^XP��Sw�t��� p͚�YȌ��q��Y6�\	�'������p=Z���}%���L'Oa:�z�4>H,N��I�nۜW���'GC0�v�돲ޟ�e����M�iaV����	<q��$���`#`r�8���u�M-!C�3��^2%�}HC�a6Ƃ�U�Cq�w�{$n�]�j�2b%�o�v��lTL�r91~S�u���B�Y����,�{�S��r:�L��i19�z�
b�B���@V-\o�yAⶄ,@" ZJY�ZU��G�Y��r~Χ��=y&���`OR֎e6V#@�n{�C�� �9/�j՟���t��A�q3G��֐I������Q1t
�R��`/ � {ц-��+z=ͥ*���Ԩ_]5�:���,`�s0t�=��D����P9�QL)��eW��"D�����x�_�jM���	8<Ƚ�5/F��
�ř��'�����Rr��-jKY�P�Mo^�4ݢ��^AT�0O�>�.X/eW�[� ��9+�}�ϝ�-��E��3�~�A yG�#�P�ޜbk�zY��8�u_�@՘W),v�g�A��3@S�WӰ�ވ�d&���@�$���k��8��s�ϧgy��^�HV&��]A{Y�7�"H�ǉ,���� Q��K�G�"��G]� ���69?6;�)7�8��`�~�ch�s�s���T����@<�s��sn{�>nB����|�����J��j؏d�O�yH���da��~u�g`��������g w��7��>��x��@�Bm�'�]�j���d�����<�ϕ�&)�*�[{&���7�����'�W�k�K�C��`/����o1w����>��v�h�@9�W�������6��_&��*��ꮷ%t���l��������I���Kr�����>��O�س<�A;Zv�!O�{r���k�n��~�TD;5�n��u�yݼ^|�� ����g�i��W>}��;�]'mVk�m�9-��L�VR���/��#�Z<`x1
�ΰ&��ԎX,r�u�K�9"�����L�]�;��s(n�A�4����k!2�ðw=��a������|:O�zѹq���[_���	�-R��>͉�z�|����=�c���:���K���Sś޵���Wq��3�Pkw ��������g������d���,���C6ଘ#Z2�Y�:���]��;�
i� wk��i��1���5�x��;ٹ��Nt�D�N��c���i�f�C��A���>�Ƀ���SE��#!����{ݍ����lL�ɶ|���w<�bź��E|O�&G���tw�c�l[��� �хEs�|���Q�(.�Y�Ύ����^��g�:r���,h�!/=|���tf/��bz=Bk1�#�=v1������{���g�nΔ�Lt����/����, y����ez{�>o�(r争���s�`���Z�c����7$��i\���S�=6��h�05�k���:A��]ǡ� ��g%B kN�����I/�K�=_�����g(=7�ҏ(7���s��.�ς�m�3����^�>]�2س�K��\v��Z�\�	(�~�d��B�:-*����\�72�1�%�� ��k�h��Ͳ�Ԡ�2)�֬ �J[���Z:PJ(7B����ZhT=a�=cA�ֆDd��l:&=���\���f#�Rх�i�]ʙ��2��a<��;���C�EcFM��t�3�.�Z�f�����r���#����VsU6.?+O�S��L�,�U\}P8�v�e_�%X8�Z�S+v]؞�IA��������O�����\�'�#/ �o�����lK�SYgR��n	�V��"� &8F��d���҄?ͧc��������I�	шJ�ۆB_f���Q���{9��-:�Y��np0]k]���{����Ʂt�q��ĸ�K i�g;�����g.V�0@���n'�����"�{�TNܢ��_H��8��^è���F�S�zK��C��t!WϟYWϠ]��0�I����(nG\���r�[�uj:=?��I��t����=֨r��=9^-�(gag]�օj����J�M_c��yث�s9˭�-9���}�Q<�i��^�f����D��"�KxL��V�]�� �.��E��9s��pm�g�$�n[��@D�v�c��)�E�^K:;��ɴ��Y�!Lc����]b���L�(苵��%���i����0�v�{}�lݑ�%I/��r��5����5]vU���}ZA9�c���j{�خI�+��|8��PC�-NF{6����d�+uw/P� ������ACn~%m=�5��� ���v�٬�v�/n]�8^��~/�xe]ۉ���%�Nw
��v�~ȂP{���O���=����:HO_WA�s����׽�����{��f�^���"�&�d�QVs�� �a�{-�-_�f3���Qh�"��Pe+h�﯅��1:��ҏ�"U;���Mvn�}Ԃ��U������ ?��M��:uۓ3GSu�
�_[I����F�%�Ǎ��i��vn�7�9����\���3�8Tk��8<�tT�����2��Q.�6��^�c��,ǂ�SP������_ɨP/K��#��}�s+tc-�M�z,%�+ �R�_I��In��$���A@��"@?6��b@��x��G����O��P��8��\K���!�$�H�g�������E�J���ø�#�7�1�@p���������8�����Q��})�N)�́X�v�M�G2*X��&�-������gM�_���ل��ȋن��:c�Z<>^�΅�5�3���^$<���(�2G@#ζ�@ͭ��|�#��	�Z�k�11�{� �r�K��5/V��a���붷O�_5�y!�vh�|f��@���88�`��2�ݾ��]��*�P6�XaƊ��A����iw��1���'�V�;(+0.��"U�����T?�����yӻ�vQ6���2�0�ט`/՞�?��^��N˚�p�V�"��c*P��q��ܴ�;k:m{/�٫;�m��/��V�U7+n�"V�,�-�L�j�({ݣs9<bז�`�uwY�k.T�-񦘅q�-]&�c�K����me��u��M��d�7��cm���E�)��
P������L�;��8���gJ���]��Y�����\!^�Ƕ�Z�PFsBd��@��Y/O�0v��[�hG�{ Ր��`|���캓�/�������~�c�M.
�+3�|���g@RT��f�c3���k�?ٳL�hlOʜ��6���3����+U�3����B�xDQZ�M�I�

G�`�G�*��r�dn������b�\̯k/:��	�g��,�#˜��u�VS42_7ql�uX�fc��d@T�p]/�����xhI��c�� >�ʪwK���������q�P8v��_ӕ����';o�Y�v�Vl�Q@e�Q�4���^�����.�qHs;k���&$�[u� osS�ػ�|�3$�%!�l�ٲ��!)�����5Y�'/��X���0w쌗�0���A \��u@$0�C���N��9g?)�9��W3&'1pe����x����Ѯ�c��l`�f�<3@����t��}�<SSTi�����K�w>�̝W��)��-)=�RuS��yݼn^?�� �?���������^}��o\�!?��\G�������e�fv�:�"���#�Z7�����Ĥ��� �-Q�Z&�Uُ%%�Σ�uU(_5�KX���C6�c 7��� fY,�����≤@g��t�Q�:2�btz�U#}��#/2n�9�sG*�@3�@��u��g�;��M�w{�XdM�o�S�l�ݭ\OX���q^��*>/7���I���L�Ɵ��l�7d��z��g�4�;H���Z�'	��+�G�F����pe�������>ȟ���Ł��k7�Pּxދ���ͽ� 4���]��V��o�g�m�v}�ݛ^	t:b/�3DX�&2/��*:���9L=�&���y�[^�V[��֕�Y�N�z�H��_������!�!ևB���u���f{t]�Ousߥ��1�(���(\K�N ���{/V9Pc����[qts]�\2��l��o��re�j��L/g���}=�л��fd�d֮�~��z�����;hA�L�@R�'����:�����ρ�r�l�7�F�ӗ՞��\�}��v/���,x�M�EP���^�}���,9���?��3=1�5^���u���`M(�1z|�(����_,�e�_�d��A6� �Q�a�9	�M��OR����-5�Vv�v�T�38�oP�h$n���]ޕ���9��f�,g��~�ud��ܕ}� .�#��S�2Z�$n��2n/;�JNB
��\�������|_>��/�������3�>�|H�v6�-u>)Sg��}T,��
�ݍ��CE%��X1QI⦐����3"�B�ȳ���R8P2�,��^ (��~+8��J��v��EB��/&�z���@�G=h���1)i�ô���SY4�8Ztq��A�H���RY�K7ڶi�SC�2��/�����;w��w�sۣ��l��<���w?���p8��c������5��ٖ����6C�|Հ����(���
��% OR�'�����E�-�����G�b�~(�mw�ğ&�N�mg�R�����u�u\Q6��Ќ�SOF�0�U	,}|f�ٱDY�#�E�0����U���ޏ��;1a>�ʥv��Y�������χH���y��;������:hw8ړ[����uz7$@���oE��	�tB�w j�nJ��ߖ;�Q���L)k
�PHF�)u���6$���Q�������\���R��Y��S��:��W��#=��D���k읬�r�&t��iǚZ�Y��d0��q�~v�V[�)v���"{q6�X�=Y��Q�\�Ͽ����i�ZU�V�Ȑ� ��	�@>��b=�n��5LABb^��T搬�{�:"��E�Δ
�� 'QdIh�h���&��IP�����E��o�s��2cr��u��P�*�s��ậ���S�w�w���/_�l�y�U����ھ�i��Lru���|����9�ٱR����+�^��(���?ɭ��4��MGVe���� ̓��4v%l����mc�P�x n��ɩ��y���]�}��|�g����˱f�iU~��Kr������O��pe�^���P`���³�d�p9˟~�����k(	���8�kv^бp$��J�|��]v���Wvp�x��hX k��&�w�t���!Lr�?oz^gU|�Em�AD���$Y�1�zZ̑y��y�?�_�T�g��<�Εb��ӌgӂXct�ƄF�97ni��pT��0�I���A�F�΢��ǧ�-o[óIN��R�L�z�2��A��@���1��џ���~�����ki�40Gpn-��S�_��� j%�g�v�G�%u �2�~q����d'����z��镥�g��T�1s��0r��?eE�A�q;S���]������Δ��;�3e��kSȔ��a'g��C����#&��<�a Ĩ�QB�6����vp�e�����$��������I>������\�*����J��Wf��z�-ٵ߻
O�Dx=7}�l�)�y=���?� <1ݪ� ֕l �lgW}����OИ�m�� r����#Y�Tzp*�`����=G^^���m��l��-A��w�f_G��e���hC�NE>����G_����u͟l2Dn���MԂ��r�K�LT"k<-�v���2U9���;+�oh�	|�n����:|'�GW�>�O���K����£Z!4�>�f��p����H}󻋼�����i��-�d�����(�BhN=�����8���
2��J�
��eO_��@�J�?)���ꭗ�Oe7�|��B���`�L���9��Nj����˽�|�ߑӓ����Ig����t�m�0O�����sM}@�g�t��?��\�k����cbV!6�H}��Tt�����ü�?� �C۝ؼ`�#�2g�z���7������8��Ŝ1��%H_:�]����#si�f�g#����z����0��10����+?+�[��r�_��ߗ���/4�.��g�Ϟ��|��K�������xy�l�s�j��}�O��b͂�x��2b�"l������x��CZ��M٨�: ���.U��7�(��F��_����~q���Iһ�����$<�qk��d�f�#(���;j����/�1���~�O�z���4�χqx�>�:��^���T4AR�К�Q����ʉ&r�,���AA
 �`����AO�X�l>/�"m��W�����op}y��j!�D��=�F��Y|N�a�5ev���7������p2��m'i���WcM�憎{����e�=�3��_S��J	8�Π��7�ņ�X"��3}P� Ў��|�e�Sw����o�ӷ�����n�D0���u�yݼ���� ���g��������o�g��w����y�~Uʘ��d�s
�t���E}��-��S+vw���$D�uL�2�ѯM����:���M�-�7l������3լ�U,^P��j�`K�G����5�D���_@�fIgț���Zh�^� ����0�~�	���HATv@X�h��l;�bS/D���u_�~9����"��I����(4��=+,v���r��D��[�����w-�xd���YPN!+�����B�"X �"���V\
k �I����tzs�kdW�H/�ּY�6��!;��bI�=���_�+t�ә�0gp��:��q`_�LN���=��Š:��|�`N�]=��&^�-�w�!_3Q�H,Ya������.@M��<�n_��H��Gw��'���[EBgH�)|}�:�V*`a���+���b�m���p�kݣ ��2Y���z@�l�[pN���}/*f���ؿx=�VzT�-�2eRsOxBQH�,U-1�ڎQ���l*�(u6�ԓ/�\�J}�5��-0�0"��-<:����L�ЛH�f&���L�r����&��� _�"�6��������%�+S�s�������
�D�������!Be�A)�jK��y�|@�4�����gvF�&^H5��$�Q�FR�:Z<��(SV#ѺKe��^��3��,3]�Y4�} V3��/9����l�@��Q2��=�ू�:V�"P�Z	u�W*k¬�r��Y	EeN�ס�h�h�3�h��1�p�z^�G0����DP��3�ΎLC�-x�fsm�C�9$5x��)j�r���3��Y�cg�Z�s*�O�a�g��8�Gpf���x)�&�"��>�
eO�[�{�����VDm�vkE�I�}MDW�kz!l�o8�(>&+�7Q �gQ
����N~�>���3)A]�Rx{?���7��������t������|�޿��YZ�G�ۗ= ʸ��p�o���+���������|�*?���}�����k��E⃿�BnF��9��eX�rq}u}���׿��۟{�����=y���K�e�M������{��h���g��[o|[=z$��|,}��$�l�s����p�ǇY�{������.��@��)���q���(�,}n����3�Ej�l��U��\ �o��i"�����O/�I�dq�#��(�Z��Y��Y��>�1P��_�����u�?�'�\��ҋϦ�L�ϲZQ�H[+� ����z�cb�'Q�;h��
��"3�w��k���g:�M�J/�s�<iֳb��P6��-�3�}�)#��=�BP0vd4��F#?�5A_���fL>�6E����Ϩ����>����x��2���ψW��� �0H��W{�qM=`ۮ.�~���pu�wW�M�/g���
:E.����<|g�-3�p�p��$�^���l�AjYp$Ȝk�ϥ]os�0N�%�JVLJGI���iIj�B*8��wy^��Q86#��y����v���{d�4e񪃏�{���((��+ �L-�c.�S�Rz�>���?��|���jehz��pmk~�օL� �O�H�C���`�Pm��[���q���yW0�k)חbq��#�t.'ȓu@Vne���5���Z(؋�iA���$(ri;��9f�t�}�Y�0n�y�r���Q�j�{�w����=�_�8z��C�&uݢ�34P6����
W(���;�e��M�<�����i�������ȆcqJ��V	*}a,b��>n���:`�m�v��q��`;)�� Z-���滏�s���yF�$��Ϟݏ� �@��g=w�N�-2f�θ�����Փct\��
PZ����}�ʊ�,詟z�>K^�{t�ş+P�cW�O��L�/n��D��+_�B}啻r~6J�
2�����Ç��o]���>�3�f��O2��ʊ8�f���]�n;���v���	�����,,^F� � W۟�؇���v��k�-7��e�g���ۏ���RE�� �^̆!^��U>}��7k�q�|b�g��jc;����F��G��Y��	��Β1��,�M�e*�{)37e�a�w�J�[A���ya�L9 �K����{� /�0�^H��v�yl �X���5����g~��=w�����i�P�c��arց F��޻��c�A.��^v��C��85>��7F���ۑ��.��@W�i�&�kEΙW���"'T�:<�3��PSֺl��L�d�{n>��IBhk�4 G�M,<\~6q�������>����P{����cxq������#�_����5U.��,w�b�+/�tWvgdj����|j��,����gM�g��D}3?���[�N]�Lp]������m�:�cg�[4w1xz�� (;��'�5F�X��������}�4��~�5y�ޅ|�Χ���Lvʀ��I�l��t��-�{P���/�^���<|��+1M�;i>L!<�1�B���-
�p�+��+_�8y���n>=��wx�׉�c����y��B��7��q�M��Cߋ���~�:���K��:�������ij��L̏�כ����u��� ��9����|���^�1|9%�9)ǬQ���I:1�1mN��NL,��c��u��#�)HZ���:���^Q<��6��(r��ҍ"$�͡����X����:�?=T�'�@ݔ��gQ��n���?蒓�N�^��& ��V�Q�C8��<�G��
qb�85W��'�������,Á�Z9��.h
�u6��u5�8��m�Q����u}��H&
�KR�ZzI���ł+��vG�7bb��Id����烃k���&J�\5s�X��X` L�i�RLZQ�͑	�:`'�� /	юj�@ c�i��DG�梪/�.Lf�f&u���3�@X��)�5	;���~�z�TrHD'c����]�	l=5��[tc���Mb��1Y�TV����`ge��pTW(9�g���L�՝�o4@����,e	�;�3;�ed��D��^�i&���B�8(f�0cAR!��⾹E3�E=#3Y}�&��f�Dg�m0+�zR9K�9���(C�����&ԯ��IE��Ncf2��E�%g�9/jG�6,��\L���|r��^t���P-�Z��
�#Vd6t���]�����}hw���'龻�}�63�£�+Қ�ĩ�u�r<Q;c�P�%�T��4��gR
;6M'�<�=��h���;��<�\�d[g-&����p��k|_)3@ ���i޼���n�R���y�@eXS����za�:9)�cOl�Q�=5t|��(��u�� ں��ԅ�Z�?��4��n�Q���%γw��>��Z�� �g3Ҷ���}#l`��H�� ���́zp1��v�`A����&SK;W�&8�[������~�=�&�ΐt�������RW (�Q"�+����=��;V6�ۊ݇�0)a��5�� ϨNU �]V@�%1鱰�3оCN-��n] bDvu(�a7�z���o���p�?���B�n?}$�]����# �y�� ��8_^^���P?=��m����C��Xⴜl�e�"���ܞ.�l7�h��|W�v����<n-:�(��o���]�L�i��mW�nQ{6�JT��)҇��A-0jN�X7��<�1^,�.���@�0%O�~AC4�]�=�8=e�%c���w�jw�d����F�N����s�舂��@�bE�
�N]�Ż�Y趎��w �w3)�-A�ص5��8��5a�Ѷx�р��f��
 �Iut냸ϻ2C%���BMO�

Z����I\�fV
���?P[mzt	�nf,m6;{��\*h�mk"�4��{q��/�I��T@L�s���$&a�Q��P�a`;M��]�>�5yV�bI����O��<[!��l��}0[� &��#w����ŋ�
\+����uz��g=Ď1`y�G���ɾ޵�X wmt �!�U��8g��,Ψ���;:b1w��x�+u�,b��k�׶wd�ʌsxՁP���m�f�י��H
�٫ɥ�U���
S�Tg���ا�"�bt��i靻�q靭z��h�Q��������a�̲��{��x�Z.���T�����+��L����#0����d�H���
g�����6��b�JFA�ڼ��{d[+�)��\�!Xa>P7BN�{�E:h�wa���ԥ,�h���Ϝ�X�BG[�什�K�b��F$�+�����FV��O�(Z��}�]����y4�+�]c��^k`z=v=�~�2�h�*�lU�w�!�Ꞻ�/?'(J�>F��ӂL�@� O�-�5��X��jo���������{V�YS���X�FgzD��&8"t���!���A:�3�T{���İV޿��kיۗv�G�����Or�:�ŭ��>Mr�;���v:Z"�Ծ�����hkH�LN)G6���3��y~F���Zn�q���u�^[�[�b�nj�6`�B,ٹl���96�Ξ����T��ΈX<�� �!.<��2\)ˁő�c��]�
r{/�W#�.�?2PRYe��K����
R��/���e��@>�u�	�L�q4�~�v�cN�`�$k���%2�9��M쾥�5���L`�
K��#�2���[��-�u���Nʾ��!��rͥXC��3/d�?�30gfGt�t�4G��4q̌��Y?I�?�#A��g�y�b�=����W+��3��1�~�u#���@����а�^�����r�]���]�]��S� �W�S;gXK�3vI�	��B�j>�V�q)A����L���Cב&����g�ٓ��5K�g�g��lo�xl��S!���u��N��Un�M�t������:����d�#G!��u���@��B;
`��s�?�|�=�>a��=��ޜ���˽���g���m?�Ph~שj<��NeXvqz~�voݚ��Y�þ6���E���&#�(������c~����'�U�;��ǟ�؟nh�o^7��׏��I3 �k�{w).ώ��'g���:.��\[�S�o8|��g�Nh]�o#�p��5�QTfb<xqO��B�M��l��sG�{ǋ����fv��f� �*0��@�����$N�@�U�.�AO��7�+Ꟊ�^�������B3(�&b���dOA�Ĝ��;8{%8M�� %��@1��Z�1�/z���v�ً}=�*���v)��j�y�4�-5��m�Z�5y�&�"�����0�-2��: vm�N�����Rt��"pfm�Wq]�liA�����5C�+l��o*,j�L&|΃�RFG6
r' 9�����Ѳ�g��
nR���+U>�60˲�=�q9��mEt<b��Q�;zj��@80����.���s`�Zΐ��Lt4R�Q�u��Һ�#M��Q���(�U���j��^��`�n֝�B��[��&t�$���E�T�r`\�24ZǺ�[�����i��06<F@�𨉢��s�l�ͱ������I8�L�>D��,���F'[d�3b�ý2� ^u��Ir���gݰ�
��e@n���*�!��;F8Ŋݩ<�r�4!,�,�d��95R�.��v	���@�:��P(W�dg0#���x�ER���Q�iN�K3��q�`��g�Y��M�eCj��m'偉K:[�v����ق����;#�,�O��+��kSg�i��ǿ�1H���M鴭�~3��Ar���^찄u	��-�]g�l��(���!� �DPj*B|�]Z�Y	L �5₮�����"��?>|��im>3?Y�2�	�0��
*O�q����:;��o+����&�T����BE�#;�:_�81ٶ@&inu&�^W��T	l�L�z2��C�\z�T��94�����2��fB��HkD�$�.�Ǐ��::�Zu��o��D���g$��L��'�i�D��l�3�b��]Agm�<K�E$�`ݔ���֬�������C��_\��_<n?|@��J�o���uL���rW,�N�������;j>�f�j��
��ν�䟁m�i�laD�
tU���̎��u��"�5�o�v�q��(� ��$>Sגɤ֤��� iv6�3���,Hh2V��6[���"k7e����n����W�dO����ex�R��չ�����b���f�ђ��Y��:�Y�h�=� �9�d���i����h�W�Ϥ�D�۫6z�����A"0�I�r��]�	-��	l�OsE��Ρ�@��l�vy�R�R�0t�n�l���O�I||	
>z�A���+�#�>���K�2�m�?�H�!�AQ�c������&_�e9C~H�Ө�V�e3�9�'r.-�` \-����#K�gP�gRe'�>����?�w`����L9|>QTc�Im+d:�Z�$��������@������ȸC����`����)k@�����i�c�����a�k�O�mv�{`w���|o�K"�z�5��?1�d�׃њ����*2tR{��;8{
�9�&�����R#+��m�\�������e^������)��[k�!�S[�K�����1�˾l;ы���SF}̘�-C��EE]�{��Ci�탘߀L���0W0p_'�Q�la�����t�1�%��CLf�p�;�Y��?��v�P�c��L�8� Dl2�vE;�@��-q�@UB�Š���H�-=�����R�$�7HЏ�H"�E��C����I�=���O���KALkT�R�Y���m�t�	��fF3�EB?ӫ�[;T���[YA�j�1�.q��嶘VX?:�8h������јϵ��u��K��Y� -��~p��I�a0k:���2���ϖ�N�wԋ�W2�K�2�X�b��YW�:��¸��1�m#�	M� �����%��h��h�c�@@�V�U:2���ٸ��/�YL��ם ��������` #��ɝ�6#����[�7�wѤw�Ez��?)�ӑ:��v�T��fj�̐�8�r:��x�m��S�WTϝ��_���ʵ�TH�t��4Lg3�%���z�ȰcR^��\{��F�0>\e{h[����|䘡q�̞]@O�B�ɦ?mߠ���]_]�	6�Bv�v$_���p̙�:�t19SG0V��VκGQ@��w���7�A�y6�˒�Gl�?V�>;��q�Q�;C��}锩K����ٳg��� V2�,���f��?HD��ߺv��G��8X"�?#$�����ӽXi��l��0�s��t�i&؍���yC�^Z����j�?�,}�b�4'9 ���f�81=��	9��֮��eHHf1K�ɕ2%�&���|��`a4�����q�D;D�%Tf\'��=���,	���8Ю��1 �zZ�T�� ���L���"�'d'rfwN���|>%�<��������'�y�;���)�߼n^7����� �J���j}z>���^�e9��8�h�R�+.����/��Q��[p�8A]������I&+�Y�d���|$i�ɭ;�� F���݊�Zi�1�͜v�4C�U����򋖴$Iv$5UL�	9ߋ�8�#i�P_,1�f �<[�xAՇ��b�s����hW������%	4�fPP��+�P��hC�i	��c���$�5�'�uf��e X�#Rv萩�|��$K�-	�xQ�d�Ĵ'��Y��`~;��:��pn��m�4.썕5�($�g�a�B�*O�٬ue� LP&\�بd�PI�(��Z�vXY9�\�|%��*0a]%t7�v��4�v\��d��K���&�!���G��Y�o)��ƀ� �����;�k]z[ڠqS\;瑘�Fqe���v8�M��yl��U�`E�Ly�B���-�֢[���F��\Fv����F�`��f�:Q�1b ���%��h_�ö}�0ȍ�s��'�L6+@$��|��	������}�ߧ'��'I ��ǲ$PdR�s����ʞ���L��N���|�N�Z>_e�h'���-҆�G~D�j4�� ��oӡ�tb5�y$�hB��V�L`�[�<#�;tz�E ��@��XA�C5R�7W	�Bt��ghv�Q�n�/f�S
R@?��N�����E��Q4��x��!E�#�e����Q�����(�Ij���]���m�5���/�?�N���@6�B[���PX>���v*�:�@f+B�lB���"�\�א$¨��ٗ
�iL?�	���v
:0`��%�t��co �0έ�M�.͑�)��<S��Ť���O��T&N�S�2;��S%�'J�Oh���[Kb6y�5�Vg�Y����v�
T�MZ���E]A�N���qCF@��k��BX���jk�����b�]|m��&X�w����k=�N�g��g�=�i�\u>�%�Ά��r�?�'c��:�#�BJQ�2�Dpν���P�[�i�8�w��ڠEd�co)����t���(yb�O��O'��>B�}Xx�d��=���a/>� hLfr���S�L-J셧S�M,Zk��Q'��'����P}��I��6p�j�4��0��W����ږK������z8�sc�5t�zQ��9��������-u���F���,a1�.�'o���
������� �eHV�e!H��M�{�V ��޻>Gf� IJ��)�XǸXѩ�O��aH ���,�A�ޟC�1Z�Af��d�Ɯ��`w��t��)�n�uU�]$�H��͙��
�X���ϵ�^C��µ���^ _Y�Jm�����X���ܮt�=��O��Uc�MV�;#�����P�8XG�l�E��P�!�d�B�n7���@qߑ ^�w,*��_A&�!# !3��z���=�����~��;ә%�s_���#�x�7��3U����;z�'�'����>��v0�@�S-��u�G;���>C�gn��^�����\�8�]��p�"!���O�F��XI��3��~�lebT+Υq��6�/�������k��60��J����c��ʭ����O�Z��eg�nt�SESG��0��_�t'��NgȠE+{K�8�J&�5b9�M�}����w7���^� 8�3��,�N�j�T�(�7z^�`A�`R��ZǷ���
�vP�!a���`1蚴6C8)�vӚ�ϩ�/֍��@�늂�Zp����(C�� �%K�ۃ�L0ew[��:{�n���:��x7q��+�${
�?w�\A  󍁷��G�y��;(�}/�^�j	Ʊ�ӧO�O�����Q1�b�SHY��e�Z�ˣͺ�.[��>�ڹk~�]O�?9�!��w���.p-��CQ0v_E�6�G����Dm�&�0P�&�C��{�#.ϼ��s�c�3��Q�Nh�{�,ע#u��פ���ۋ��� �a s�23����j1�Hϟ���k�@8-Oi93�f��Ϭk	\4�Ͼ�"��2����v����-ޣk�~�1�t�$��`ϫ�hޅo����V7���>&l�Kw��u������,�2=jg��u����A��T�Z���\Q2��������b�|�_d`	�犄���S�=�X� �i���[m����s����*��oߒ{w�I�i�~������,��� (~��K�l�=������
��G�����շd_�������H �G��i_������W��T&��t�cO�y8�Î���[
&p@�U�n{<�>��kq���F�.AÀ�3����x4S�[ AFc���)E4K���`8glP�n#*�q֞k69,������BB���x@wY[ ��@��ޘ�; �׾�<^ݻ��U�٪^��#a�m~��2n^7�����o��; ���'�������ౖXG�$�K�^*C�wJ��1��s8�
�e�W�K�eSi�f1d�擖%�)���v1%�
�@ߧ]�^���y.���x-��i>�Yr�@�Â���zS���!i���������iRES�iW����C���aA	�����A��yT����<�D��N��/�����4g��i�S��u��B�g�c>��,Q��?��&��]�.�٤i(N�:�ӵ��͙�2hZ2�3%�C���_��%)o�������,^��)e0+�5�1���q9����̬���ڽ��=�Z�uՄ����v@׿�)F���������mNg����l]�ʝn(��\ZPe7��i9��w�{�� �fsTty����)�A�K8�S���p�ɲ�b��?Zn52�����Ӻ��k�5T0����Uo̺n�z�<#�&�:��"ѧ:�)�e�f7�8�C8�k�58ě���S�ǝ���v'�kB�6��;�ϭ%���2j�Q�_Nr��*֢���&Wq�Sl��df>�J��A��h�amn$���z�:�L�A<�C�^ \O�WU߫t��2�a4�����Χ&��G�����=Sٍ��
�I[�S{߬gF�I�����k;����uGy��?��b]���f���E-����ZMl�]�-vYNaI�1��PGX���t�n[�v�RNMj�p������E�Ew�0�L��1��|��`E��dP(d��G�ب��v�؞}��d2m��gF�*w5�&1mM��>��C[��G�����i�`���ĥ=��=��JKZ}���|ܵ�lj�h�njK��>�f�3��v�T��t{��E�϶��΍9�ZGi϶o��h"�zi�0�C[���{�s�2�� ����� W�#��h������Np��:Sj{��f�BM�e��Y���Y�j*��j$-$MO6]�֪�g��\c�Pٷ�v�`��&�jL��O����ڍS��x��,�l���� �<dC�  ��IDATZy�]$�Zi5W�ْ�9\@o�����4AT���Ο�b�	��ϛ�<d���Im�t��u����q��U�E�8+��"��þ���4���t���9�2jw=hC�4e����>�Ҋ�����>=�-�,�-��·f���4;��bTkVe�h:bl��|�Йm7�Ͷ�o#-�����L��&�\�'�9�VTd��oe��[�FS�Ci�0�̆z+��xh:�IM[��jb<�y�M_��,ÔU�
�������4a����Ÿ�˩i�fS���-v��Ƕ�ozE��>�ʁ�Of�ڷ��7�6Wi�RSuM��%j[רs���2�rViz뤆%��N2,��^��1J�c~�\G�=�)/���t�jk��F.��,קC�Ʊ�a���VZ�y�P��,�� �ЁrU��������h
��Kێ�g���k���r[�/�����T�J���3U��t��Wm�I�󱝺Q��˳���D�������{]]��1/�:e����
��leb��u"����Q��T֢`!��h��ˠb];���&9??���ؾ�t�����v�a�@pY�p��<�Ȣ���M�jRВ�@�� aע]�\��J�ʐT�+��ɤ�6�����n@/�iq@Y����V{�ݙ%!����Hr���녴\z�+�:��h�]����xuue�ʿU�X��`_B1�Î�މ)�'b�$^������Q�O���o{����������]��n)�`���<��:}.ݻc{��q�]t��bSD�A�V]�#�n)38 �@/m��z�ہ)�= �%m��#2v Ǟ��u�y�abR����]�xN�\&K��+R/��h�uu�D�S�Vvk�ׁ�2�V�nB%�
z}�V�� j7�Ȣ�'�G�tC1�����$2@y�E�9�>=�����V��V��B�x�l^����,>Z|�8���	+۝���9��⌲+� �`�=���3�og�8��˵$�1/(R��j2x�rd	w��MC��hr�nv0j� �SN���&!�G؟����9\_{��Ё6N��  MR/9`J9�d�B9
Z���XX�=_����IB�4�M����9f�H��]Q�
��� ]q�kW! �����7��y��@V���[���2�K��VК��s��4���)�`f�w��$��l��[tj'��Y���@��3TX��- ����q�	�#z	�1D�VS&K<[^TEgu�z��$�������Z���s|}Q��(���&��Fa�W�_�d�ܾ|����ϲ�?�,nIףV<�;�o=�����"��/�Uʏ��e0��^�4��>��;��W	�2�@����%i�k;C�K��!&_�[|�[�z�P���R��~i��:��}�B@��b�H i��������I�6�������Ɗ"b@r��1 �<��,!�|*,�	�10Ee�!ǀB�z^���g�s��E��0t��@�0P.��$;@�ݷBp����3l{מS��9�A�@~{y��A��K	"�0�c�K (�θ`�U9
ъ�]����o��@:�-����|$H�Ѯ��rf.1����:����ʀ ����nsf�:Ƌ�62�����&q�3i |�ty]�:�ul�څ������]��'���/��|=�/w��޽_�<y*�?��=��(-�";�h�~��i	�]?u�d?}�"��fGٻ��:t7ѵ��@�4���[w���{�_z'ڵ�c�G�j�b�����J�?�����9���dn���`�@,�C�������A�$�"}ԅ�p��'}/��3����=UV�~�3�CE�����g�ɦ2��D�HϢ����Å=\C�����}0ց���{h`���AIsu����o^7��������� `N����o�nݓ)���;E������?Y~���_�8�����ҟ���9<��-����?	�x���o����K�ʓ�7�������b����y��_~#��Ǉ~?ͩ��>��~�t�;��Z�Sz��ß��??{<<�����+r��A����r����t<�}خy����������yx��J��}P^�{/߿soy���,x�����~�������5��I�w_.?��?���],���o~A���<	W�W�ᣇÇO�崄v�կ��]OˆӸ��Kz�����'������O�:'���j���N~���|��Y��>�%�����?z7�)��4�����k����~�sK=.��>�G}�ԃ���i|��7⡜³ó�3���|n�ү~i�hku����i��)~�ݷ�7��Fzzx�����b����N��/��r��E���G��O>��sz㽷ғ�I;�8�}��ʯ��Z}�����ޕ�O���{w�w�{'|��C+�{y���u/�����g�kw�{=��}���������Yl�e�8�]?��/�;��xu��3�	����?�Z:�S���qzv��k���o��o/����'�=*�..������7�<]���O���������?�������｣ ���M���'����0�=����k�?�����M���{���g1}띿�����-~(QK�g�Y�G_���b7����9��T��z�v��+���ܹx���P~�׾�oO���k���.�u�<� *�B�/ߺW����/|%߹s{y��{��t��
�/~#-sI��c�����K�����~�ӟ��>�h�����yy�]>J�3Bm��;������^������ ߹};>{�4��w���\�+-p7Y�P�������/��R�w�xC;��)����}+=z�dZ�j���?��˗����V:;}���������i���V�}��pyx��JQ1���~�~�׾�%����o��]�s��F�R.�vwꭶ����_ɷ���;o~Sn��R[����v^��K]�.�ɽ�{e��_�����+�~���<�W��wߌ��N�%�����s?��yW��</���/�7�|3}��o����>�~T FS`���W˗Y���������_����NzK�?_�O�|��Y<���s��|��/��+���rz��iz�߉����p�_��3ڲ�:��Í���t#9� �@�$���HKk4����k�ϟY��Y�F�ؖƶ�%Ғ�%R$E��(�`@$��_�|��g�ۻ����="�D��z����;�Tծ]u���o�bXG�ʯ��d���������`��x�9�zΊʄ��F�w���wa%?��`��Yy��i1?=m������U�WF�tM#�C[9ݚΏ<����{��|qyQl���Kg^��i�J3i�V`��V	_u��kr���ګes�auG}iW/[EVX�	�jv���R�V>��+�K��o��#�[����K"2�t8�_}�j�P�7����g�5�߱F�XmyQ�.o:������4��.K�Kƅ��֫rN{I�J��K�b��=�ګ���/�ˋ4�ϼ��ػw�:u�� ��9r�rǰ��;�R�wP�7e��3g��ʂ!����+#���Bd����G	(;{�L�we���u�x��k�N�c�Ffچ#��*��?�?pD.h!��R9%m[�
�峯XI�K?X���B9�N印�9p�pl�|���۵�U�VVw.�	�PbӍ�����bign~����ߴ�⵺qϺ<ZC��GōWݘ�]ܛ��4��%��S�Z�;����%w�B{d�w�pw��~��F���r\���]���Y's3��Ťb�wʓ��{V���~?[;�ܳ�d]Z�`��>0�n$b*Riu���o�V�V�"β�v�������땋����;.R�3|�+�����ړצr��VW/��z�\�ڰ����V^�V���l{NL�f�V��N;�%����`�;m���S����̭2-���\~��	��+K���/<cz5�>�y޾нhffa�y ��l��ިH�t4�����ϝv��޳�'�����ȍFR/��hev)AT��Ucz��}����m��S�[��Y���厸��{��N'�nm�;;�byy�<s����W�[�3-�{2����w��Z#K��$���ٹiW�֫�^w.���^�w���.��|�¾D����E��wV���{+�:��ИwʓW]�{�ϻ�nq~��(��o�Li/ ��]u�г��ܟ5`�R����� %�Qf���U�*{�P�BǦ�>� �Qe����KU΅�f�lI��� �{�G�J
hy� �����٦T0�@��n��D����m'�T �� ���B�P�0��r��[�U��
N��Ύ3+0��E���G)�W՗��@HAဂ�� 38I�rV�K�NR
Q��){��Z�B�
%�G�_ ]�gC�:#둤L����E�����\-��)C/��C��D�R�`-����o�L
j5�O�I��*�TV$�R�T�eJ�H�<ɪ�k^�3 )��h�@ ��KΘ*U0X Ls����~�ʪ�����V�Y���0`�]�s&:8�yf;	���Ef����i�
�`QR��
@#h����T��Y���m�n��U��qi9S�%J&\��������Miה��`��0�@2�S�. �k�c.r%���E�����A+�K;`"��q�pVR�azU��1G���E��7T���,�LW��LA �/�D�d����>�ɯ(��9�O���8�X�Y�y�� yA}�m(�����P_\yK�G{~<��2��j��Q*�\1�H5M���J2�A+Y�&0wDp�v<�	XV�,=&2q��E2�Gy���3�#�$}�Ę���2r5%��y�@2��W(���B��4��P �P���A)&g��KJ�*Q!��:�h"�VK���(T9 ��{�(I�!w�ǓP�*��+c0��EU�J)/h�ݛ@���tͅ�n��>���v��u]%�m(��.ُ�(u+����*���sjՈ��R7Kx��ϸ�f��r11.��5��W��V��W�"T�Th"�N�����x�{:ٽ\kZ!K��B�ʲ�l{&AA},���J�Y�)I�s��ő����@g�G�X�)�/�@�1J�4P8�X���&e�|��U!� 9���l݂3��*������a�\��L.u@**H�iRypCh�D��?W~�\�R1�?�E:Oȵh��d��R0�&W �����Kx��"��s[5�+tjr��ؕ�$]��ʊ���]0 �۪�+�J���HRL���&��T�5��h��~��2�pQ(�7W�  ���B����e�����-����1)�ȤW��1HY×������"��ȽP�3�%�ǩP��G�l�"���u�j�D�v{b{gΦ:S�{a�����3:W��!w�K
�Mg�؇��-e��r�8Rc�sS���7_���8G�g8g3HmV�_�J/Er.@����U���d���gg�,��ho��S��`��XD��1XN�E��HB����Į��cB�� ���3���B�;����,"�Td*�!�!I�~%e_RWj#x�p=Ζ'E�0��`��2��l!"MUF��q���eW�-�Ǆ6V�3��M�"%j��������������(]�H��"s�� 0u������ ��C,����0�8ck�4ʑZ�7T�A��R�b(�C�ZS�w>$�n`����+,1i�6i�6i?�'E @�z�h����C[S�Sgk�Fq��A��c��o�k�rC�i��F�,���/�՗����j�?u����-o�{r{yf�i[�	��k�,���e�[��l/�gB��KU��ݏv-�\���er7y:s�+�oN�����ѹ^pǱ���o�{}*�vL�Fz�<+�v�����s�Z˫?����Ź���ټbye�3��<��E�n?���ϽV��oL�v��0�E�/��G������ӓ/��(���%�{�ҩڷ��V��<[kYS��w=��~�F\�p5d�2��������H��V��6�N����u��ޒ[����̑�|���kO��~��lm��w��dizA�S�8�DqjH]�g�����P����9[8�w����}���}ˌ�� �c�c������_�C���s�S��:�?�D�	:�CG�mF�ԝ�Ɉ"��S/O����3g�,+�O>�+�ls��Yv�X��Z��Ҋ��������τ��߀���x�w�����q�ˆ�Z9�/T�rd�|�y*<��Y��̤���/Ůi��%���9�r�y�[��/}'܎����[֌��>p�{wB?HΖ�Z�sq���C�в�ƙs��FO������=���$�gO�td��������6g�^}��Ln=qKt�57��`��I�۹Q�yi?x���?�7�<v���^u���ʬ�;�=�L��Wa�������{��+~�e��s��S���a;�-LwF��R�VQfYat�+q2�_�_�F�����|(=�tl�
��cXYy�(F��Q�_}�Ͻ���/���,?r�}ה�oS�7��Co{�������o��78����uKW���<x�8Mj�|�,1Ϭ�q�?���L���z�n�Goz8;�t`$�iq�Ny�5�^�s.n\�>��?�7g�N{�]�"��=.��G�a%�(��N�̺��;�O��퉶zV`�׹b����w���&7�K�����7�Իp�����a��R2]�ηZq�$��ߍ����~����~�/<����%>�د��N<ݮ�j:�,ׁ�^>����/x�����WΚ��$O����3�$��8t�5,���)�w��a>t���Ƶs'ҟ�#=�tFeff0��Չ=,������S���N�b����ۇw�xKd�V��"h8�h�ۯ�}���/��L5��Ԃoe�c�/�}����!�qJk�����8��놞�yi��_�������ǆ�����\�m�Fj�p�E����Ϝ�T m�[�wu|����sӝ�,�D�U�^:�������o�BN������T��[���Fl�r��(�8��5M��}���/�:�ϮYǗ�*{��F���
�e�=v�Y������|�3�]��w��S������F�뒿6��?|����`�~}��_����X�����eW:4��'I�B��i��������DY������ߜ�>z�����ii�F��&]�Yȱ�������v�D~�n�۲��X���Hv����c�a7)ܺmF���g����o~�-j�5=�T[F���</��&xV�fx��'C�����g_�����7Ә6͑��?/������O�^�:��?r������XK�#��2l;v�B��k0ǰ_������7^�vzYׯ\�=��G��e�6b�a=|�H	��{�y�3�Y;4B'^O�'�~���$�4��-錮ɤ�|��ӯѽ�_s�9(.�R������ʱJ)�k�w�]ο����s���9/��9��i������x2=�N`�I?+]Wnȣ���+�X�ݯۗ���Q���'��4��&���&���w�r���/{��5��}W��\��|��Q#p��PQ&X���n���;�N��D��}��;��o0����2�����U��Κ���n?�IW�K>���q���*��Ľ�H�j��q��������l��Wߛ-O��<A��t��C�=�K�_�^:�}wzy�WEvߕ�;�N$� ͏�m�ȝ+����ꟻw�s��[��]/Z�MQ�8qO:7=�J���ү��k���F{ލ����ox�]���'�w����j�C˱�<Ms�w���mϿ�B��׿�z}���L{�w���w��f;[�k�������_z�ƅ�SSf��Ym�����'���-l8r(ӲL���p�^�����_��R���{�)�3�e����� �7i?b3t���A�CF��k;@�1u`N��щ���V�@_�eF`�Jm��>�$�/�!.�E��2�m��
�UA{
Х����ߡ�]�<����� Bnf�3f� �W�c��@��jwrn,��
�1Uf�
p����)�D�_��F_6"����D@�}�u�)K�2��Tl���<�����W2�ҥb`D�"9й���YO*㺒XUY��A�<�
H0UC�����,S������*����^ ����W@��s�K(�t�� '
��Z� p<����d�_��9�������0%�!wL��
(�H۵H�Զ��l;--.˪�ީi`��6М���N�� W�8*�dP���*H^=#��d�8KP���#i�6�.J!4��$�n
�:ۅ[�ҽ�u������6�5p&�ep�3~�0�z�^���v�\�?�gR݀��.d��\�����|�H�b F�X�C��H!T)LN���
Q;:�� #A�`4t0�,�Bb,>+��QC�m��|ףq�<`��Bd6��t��{�7�(�)�� �\{��MrΣ���<' ����������P�T��kOK�����C3��?��3�����B��o��QVk��KU��	Ld�ـ y f�{X� "`��7�+e
�k����)(c��7☕DE��r��V�:e��V�R���x���� j��~��Ŵ��0Xv�z6��O��O��%R�6} ��C��ʇbo!BG�Tݩ\sv�R�* 6�ɫK�Jn�D_�!�@��|�.�N���Ee�HU�7��i �R[)X	�V�-�x\�@W�����Y�\�5���ªl 8*MU���@�T������y-�/�H���,���1Y�	(��'�c%�Uy}�8�K�"���E��;J��z2��~E,?�v9F��D�{`mʓ/�X�9 �T	�CI^Tj�2�M.J�ؚ���5�_�"��d�A9]��T�Ae�c/�WC��JJ�@��JI�sH�	| H�XS��Ӫ!�ta�#+��j �R���R�
�ƵT�Q͛�aG�Uf����5?�APΥ'It9�Dذ�,���j7�_b
��YW�#��]|�_����k[�R����ɟ�����P�べ�$���m�Ey���]e�S��./Y��0� �ZcR���n�sۘ���Q��;�����U��� �+R�X)@���y�H��F����R����"fA̔����!�`Htm�4_$Yr�>�>��T�J�G�]�0B}�U��#juy~�JŁ��\&�dUB:�6x�+^��n����b���������uW��n4�ꥋ�����|�ؠn�"��4��3�iQ�O/��Ez�@#�����a�����PW�?l4�C�%�wԈ�aC� �*�cq�Q�mf�X�����t(ϙ1HB�ޤF��j��3TBF��ԟ�]���VjB�.M�2���!DE�(C%E��I��t�&U
�Ƥ���T��3�R�N���sg�4�������C>7���򩰳��6l�d��EI$�E�:k+��!�{��vK�ꒊĨ➅i@����1i�6i�6i?��'E (�KQqձ���O���У����ܺ�����L���ƫ�l�V��w�{��ػ><���_���5��!���s��:�r�ɜ(2M�IS?)������?����8�t���ݻ�Rhzߓ��9y(�r7�m�w��h�<zl��g��p��7u�XXLg��^���\`]ypM,�r�ü������ɗ�8o���|�����.��-�۴���50,/�����"��y��̱c'��+��}���<�\J�<
�/2�Z���SO}c�]���w�}���O���*�5���Ǝ�ZfV����V/]����Z~��W��>��K�z���s�^��]��{&V�?��c�s�g:O?��/�<]�]4m{}`Y����fb�^2�n<|�;f�z橖�^�I�w�_������8����������yO��wf,���(]{�ɞ]��Y��5僇'��~[+��/�Yo,ܗ�YFp���m�(R<��Gv�u���z�ҫ/O���,�;u��7]�{�5�,7�g�
��0#�q�N\W{���VS���~.
M���|�A=c�L�^��;q}������o7�����'?�]���7]#�i��Э��?�ޏ�ϭ��φ�v��f��m�p�����3�76X��������k_i\^�l-�,���~���χY[��քhy�4�8��C�k�ɗ��(,3�ۚ+n��m;�i�;5�Z�M9���=�k|�>�z��϶����6����ؑvM��!,hX�(�w\u��˯~7p����Ղ�z(�+�:��R�D5�����ӿ�� |�C�5��͠'_��b�(�-�v݆˱��ǎk��?�����0?��o��8�ΰ3��5�hx5��'ݦ_��V�����fq����n��p���|)0�ּ��j��냭������*�<Zܳ�1�M͊Y�6kkk��{��ħ��~��[i4p������kn��wR'*<��s`%��?y��j���n��Mﺃ����a3ܒ�:��Ϡ�!;e�5�{���﩯�C�,��)N�l5\����(iʷ�u9W�c�a�}Ͻ������Zk�m����a��u��+�(VX�c��s���'~����Æ|m��;��2|�o��Ӎ��t|�]�=X�":^�����g*��-���:�c�^Kk��i�n��O�~�~��9�#zr�fn�55��p�4�-�����N�{=�M����W�ֿ����-W���gH���9����������L|��&��5���y�שwz��h�J-���z�C�<x㽵�zj��nz������.���YQ�lۊs�}�]����~=X;Σ�xO�p�;ǡ񇩆u�U��x�����������z�C��i��;�_�J�,-?��m��3~h��?����%��#ǱFw�K����4�w?�h}eq���/</��Ͻ�x���Zi�]/��+�V�������x�����{�΍G��o��H���ȱ�}���A#v��Q�V�׾���V9U~�cI��ߗ��n%��j4������z�p M+��~������ ��^$[>�κc6�5片��}��	��Ͽ��|X��o��P}���Y��G��{�Gk����7רYO���I�pw,�ʹ��ru�1]˵o:t�����}���M�������$��+,q�hmz��'�������|)��;��3�i7#��N����{�'.�3���O������i�s��7/�o;~M�o��0����۶[���a����w�EY:O���y��>����l'��5[�+���к��۽����Ԍ�^��c<t��IM�5�if*���R�猹� �����ϼ����ۯ��l�͡�$���s�Q�jvm�v?���g>���������;l��H�c�bJ?k�k�ǻ��ۂ�~���-W�P[؛��[r]�˱�(����s���õ�N�C뮷ݗ-6fa��h
"�q�����?�Ώz[�Qx����_��Ϲ7�v�qh��붲�r(��GOxS��Zs.l��E��g��o�/Y���]B��y��Ia����������η����x�{�g����e8gJ+�t�0���FA��n�����ɰ^��������l��kF�6�0���P:����\����+�FEښ�k��^p�(��� ~j��<p�TzQ�#��f�";�`�N��F�r�Ve�����A� x-�����8�h6D�֠�%��0(��C ��Bs8X�xA4�G�^�O�Pw{��qS�\�D�f�2(�F4=��"�$�q]�R�w��a��l.�.98H�*��/�P-�F�A��f�)�r0��TMVH(�����X\ ��s�z#kn�?N(#ˋ|�V�* ��6g�!`��3�
up��ȅ
��y�j��Z@ͭ��`��9����8c~��&�ۭ��L�м�e?�9�vt��S���Q`xm}���^��Gg�f ��!� ��WSަ�F��B����1q�j2��k�"�#ٻm�C5�U��'�m�H)a@߫�(����)S^�bN��qʪ�(��FC�9Q�)��Ae��3 =��\�)-�L���������N����i�,^�m&mL�� �
 �^���(G�t�� Պ�ʚ� 4�1 �/������7�Mѓ�����F{r>(��N�l;2(G�L��/�6����2�����` �ѕ�ilt�ɵ���gK�!Hx�V����3��E��ئ�O�k��q
�G���!=�h� �P���[��"O$iy���xv�
6T��}.��C�#&+�Qmy#�j��3Q抟!�B@N�q�9��zMLMu�8�j��h$������z�\�³��="h��?�����8%���`�({�S�^��bUj@@��B��B_��Ji0 ����0�LT�Q�M��-_��CVmg�-�
/p��Dh)JZ� ������$��"��s&_�$U�o <��F�xr�A�k�0�H�5��W��;�KS�j����Nx�ʓ���{�cd��E|Üؖ�HS�*}`U~S�_��RLa����"�� �hOH}ʊ�� �=3g+��T�E=~��\1������Z��7��!C�"�}W���8�o��А�2�7`���ׄ�7U�~<e�{�&%�Ϫ]������/����� �hdY�oR�v�.X�ݬ���Ҳ�R�U�VKa͹��劄e�9�R�9�j0XWuy^) ?���~���B�}��(���n#V�}F��S���5�;�t��"!�	�oc��49�X�cђ���
�,.�RI��e���܆0�ג�T�I����i�[SS���}:W`<@���@�a���q]���G��C"K�<����}�\����5�JQ���[^��\�>�J[����{e�
l���s��Ǫe����3l��9��F�H �N��A�@�"Q�����K��TA�{;��A\�Ø����>1��+]���sU��B����P��ЪK�2"E1�OM�-�댭KD�.�/�����_�jM�>�d�:�O4�-�aZ���z��ଉ}�p$}��N���T@��?Ⱦ�>��l��k��L�tfy���4��\)m�����4��<��A�T�Q`wo�7��t����HT�"�a^I���s�O*=A}����pFK2*��<R
8�U�#$+��"e�i��/����7�F�G�� �v�rAE�uJMV%2��-<�?J�G���D�@l��B�T^E�x[��;rR+��ϗ��@�U��}��s�x6Y@LFJϹ��aE�l\��I��}�T��H���
�Y2i�6i�6i?���N ������Խ���O�w�˖]>�w>9l��[r� 7�y�[O^�H�0DK��Qx���s��ֹ�xT�vfw���'�$�O�ӺܰvvvF��)������>�tx�����z�s/��;3��M�n7�b������p�W^y����y\�k�x�cI�w�N}9��mwl�q����n�I����u�0�SU��g�ۉ4��]3j��>|E!1�<�m�A��֓_��L�E-y��gϞ�|�M����-:}y�K�u��Wb7:�y|+�����Z���,��qW��D�O�"^ȜQ�t������G��0:3\n4}���e�W���ֻ]�ʃ�Vvk��Pt��XMS������W$�����rT��:�ɗ	y��H���}�.Ҿ�O���Q���]}��e�v �r�"u�R>�)ؑ鄣���Ρ�ck�N�0�ח�z�d#5t�h�n5�n��>:��U���#PgH��{(���~�%n6�f:��C��]�x�:�t  ^�Q����˯c���d'v�w�����6�u$_b��$1a�ݴ;:���׼����̙���s�d��Y�C��]�V�[ȷ������1�;[�����I{uG5�6x��n_u�foyfư���٨�#e+�l0^�������+�W:����% ����Ws ������z���x}ݹb�pi���/��:!��ޙ�eI��~�C��`o�۳#'M#y�H~f&���U�v{)��h���w���
��s|��ҟ�벭�4���{G7��^ʥv�5����)fgi,�M90��hT����ٓ{�Țy�l�VAH�B��'>6x����cW^��=/�I$����vU>k3�I>��ڿ���7�xc	��|�L1���c�&�x�ѹs��#W����j�خR7k�-�3��O�c'6bc~y_f%���tA�T��4�q�6�^�z�>��Tz�ųq��ʮ�77�;�y�h~z����XYXIA搟�g�sE�&�����G��w:�x�I{yy��q�|!��*�լz�7:q��NӞw���\��뒹Z�Ms ���n%���it��i[�W��L�8l`��Xyҿ}�>�ȟ[{��]������uW�����^�k\q����ܸ0���gl'[���Ã���XW\1���,jD���O�읝,���u�K����G��r��Z3�m�MѴ�o��]u� ݊����gkqq��"��c�����v�=z�{�������N����4��>?����8��c�Z=�o6����� ޤ�_�g��ΰH֓���2��e.��� I(��{��dm-����S�}�2f3�Ը3j��y��E���o�9�6��{���Kc*�u&��=����]:�=�v�w��Ç�d*�:�C�}��vJ���e'>45��~l�:r�H�E��hd�Yu	�4��[�5O���mu�\�)�}�rLy��S�Tv��eKڪ���&j��_+bŐ�����y\�Ͳ5�j�S�q�u��H�?'��ƃ^<���R�iH?�&�$U��{��u���ݟ,�����
��V��x]����������څ+҅w���F�C�
������>suu5�����n�?`E*ߵ�&�������%�-�����}׵w��Ya��H�����Z�{��G���\�ߵ,ϭ��i�}3;5j�kk�f��~|����W�_I�ОI���[���e�@��g�&��qzn�����/[�n�/,4�em8��������UQ��|TYeXl8E�Z%��!R �䠺VP�t*k���"���W�_��EW�l�E@���[6e� ;`7����9[	�x�h���8��]��猺���g��^V�oY�z�\WZ�ϋ\�ܨ�
(�>�)�YXaH��a~��b� �_�vK�A�~��` �k\�4���� )��΢oُ�����ݝ��{��n_DQB�}�W���Z�r t�X�QVJ!D��f��$�-��j��ِ�� d�@�@��L���9љ���99�]	X�f0���$
��Wz���E�K����;�]���I��ld�ebG��MsU�y0,)x����l-YZ\�{W���G�;-�kTc���oٔil��hX���g"�8,L��3�LV[K[3i�)�ؤ�pN��T�0��8�%�zCU¡�2�93��-WY�do�UI���o���l�Rm�zf5� #����r�0W5EP!@�����?��T�Y���F���������#tr��k4�4�0'<߈�#H�`Kkc�0��5/B�
�a���5�*8Q�N�����䘢ڽȄ�tZ�.���:�u��=��V��>�S����k!]  tMj|�Rlmo��|�<��xDrl � s�$�&䀈P�A��plY��.�䢲�*%�6D����>�Rk�h��Yo����� �S�7�U�Aİ�ЕRFnJ�&��a� ��נ�3e�ze�B)�3gu���^Uj0z�x��WP74�K8i�T�GI�cO ���&�9 Xu��%�Ɏs6$��K/L�E���'�J�������(m ���F>��V��(��Py��jT>B�,\M|��9J�D��c����<'~�J� kl� MA�cy������d�Rb�HA�|r�YոW$허n �y�?���!�}X
� W��5U���u��K�P���.��\�ڳU�G�3hҗ|�f�F>@�[Ŕ��D��0��
����1 �8��P*e�!�n�7/K;���F	B�"��ҿ���@����(�&�
m$��*'B��
�S���4�ar�<'�D��B��q��N��7aP'���B�0��u��g ��lW:#��v�D��ȏZ���#����"�)�Ңg�J�n`(b�.	 �lr.#T�27ʶw)8I/#�d{�E}k5ZtùLg�c��o����:\1o�1�2�����7������F{�NwH6�,�Mc�2��7�/3I�0*Uy�Rj&8�Oh����-��^��)Ր�� �i �:$��rΘ<��`T�>�`�w���l���l�y���0&p�+�v��F�*�J`�^Z�P�A Ù�u��>^�=\�*�S�,��n�����M��Ǻ�}��Pr�!Rȋ��@z���/�ĕR)[`�p���n�ϙtƣ��^��&z;}��rO��B�e����c����u�'2g���`k�BT�O(-�/*�Ϛ|N)��h� Ӵ�eaʂe��5ܷ��A� x�G����G���7#�0J� W�Q0��8�
r����� �o�I�� ��.��)�A(��&�y�;��$�u)
Ae��C�ޡp��0G+��2c 6�H��D�a�֕I�J:@�I���(1]V����8���H%����{��̃{����5���;LK����련�-���gSv6�zOb���7�I��I��I�h?)�L�L��>�i4�
>���ن�Mv���6q X���������v��l�v����[�_h�7��[7�pÛ�i���&�7�8�����##������u�n]���ɓ�7���G��V�u�V����QZ�G�6z�������v��������k��O�y��{+������~�����n�}��mo���p������ڏ�c��&��ڷ����̏�?�x���L��o�Z��b���gy��l�yJ�S_��~��]���/��]�}|�����4�L]��T�G�<d�9�eP6$�B-K�����s�hjn(�Kd��W��"P�d�(��^��!��0a��+m�9kz)���_~���L�~����"����MQ�}�g#,������Td�P��i$*�K�>���
�T���
�!\��gDH@d����v��נƒ����un%׾UA}y_ ���]����#v��O;]����o���@ z�mmQ �e��7PU��9V���
W`�P����"��	�[X\$�qaqI��͉6�t=�6��RA����{eT��E��� �Ϧg:b)Z"E��k������G�sCH���:�Ȝ\���@:��6Y-ǁq�U��d��]��\k�Dc��Mؖ�Y�!����a
�*�t�� V�Y26��* K�Jɒ�md�!3��c��i���`�~�J�_�C�"`_1���U�P�Ό�����-��z�u�*� �*eU3I�Tٛ���eF��~@���:�F�cܿ�d�|V�HHN���:�^_��"�mnn�mi�������r�M��)P�~i��ʨ&	]C�s����j���.b��@��Y�p��C�}��`��R�`��/ϧ�8�W�&����0�2���xNʹ�����X���Jd���˫��c�܍���E`�^S<�
�"#�u���b�k R���"�ӵ-E�i�={�������}��2�4SF��æUP�8���������RL�Sbay� �.�/�^�&�n(����&,��ප[��8{R�)8K �9�Wٟg8���F1�����=X V�Nw�T��\K^մ��8$�A�)Hn���2��>Y����R��)��?�gR&����f��[e�C�ee�8��J.q`)���89����&*���(��6UF�GY�>��#�?dÓt��C�k�*�"��6�� ��L�Ȕ2��LN.����qX�z8QF�cD�`���6�47���1C�lԱ4>��1i�	�S�����*CZ�D�x��\W�ϩvKLMM�1��s�£��]*�TA�5+�Pf�cUdA�?��I�	���,�^Б�����X_됝n�1��E�1�n�r�.�Y(��
G-�Ƶ&k�)Y�wx}�_ Zm�z@)	�!��T�#mT��-�}�\��)>6��Z�I�Jd5�SmZ&��`�.y�H�#Hk�bcsS�+�n���`UO�}└ �"����{le��:�'�� k���y�'U ��]��r0>����[�@��t��6dW7�u���,�& 0��P?,���qM`1�P ��g�ŹH�,̈�r��]�$�6�;=i���zkZ^[�͍u�P�|��2e��J�cg�K�(nTunҍ�p�$���!����L��,p}y�?>��`@�r |?�k �S*�`+�]�1JǠ�MmD䂖\o ���~�l���%?c�֞�Ģ-���l�J�p6�f�0������%��h�ϩĽ5��3��l�r���I��4��w�Lݦ9�} �� ����&�ٖV	�F�`�5�Us33t&[�,��斈��%�.ȹ�R�ʾC��W^��<�Xm�"$〈�a��*����D4�d$�}*]Ce)�ʯ�\s 3LI��5Y���j���sE�w��b{��vQ��"������ �T��gI�L�1����=�����8*H9&N���2"2���SfLf�2��.��U����`b�
��J.�u���ZIa�$���	d}"�"���0IgQ�q8W�.N#�����h�3<7�Co(|(��������3�Dȳ�| ��� �RIL^`��~`(�"ۨ�}R�p�*�aB��I��I�Yh?�R�_wg������C��-޿���ǵo���-�ǵ����MڤMڤM�O_��{%����߫3K��C��~'�g�������U�t�U�3��:ץư�
����v$iw�bY�- �-\���H�S1T�)v�JJ�/s��k
#X��WL�\G y�l-�$���\4��X��⨚�J��@X���,�_p$L��*�	 j��, o! +�7=�� M��>]O��a�,U�����Y��O��M`���.�J17;G�Ph�6(��uרoB�����KUƎ��U���*C�PZ~(��n5U�gB�T0�a�:^��\!����lY��;�W��"b�fi���8������� ej ��P|YZZ�ll���k*��k�"�YI) qew,��K�A���]Y�%�)7�E ���p 2��ך�	]W�m��eC!.�7�q����+���C ��Aj ��f ��m
 c Pg��E��y�2�Zji�r�6��_*�n�P-C�����8��%��f�|�@��2g#����#eh�J���`v�TMyz'E ��2�E�����+�pI8k�	苔;2{�(f"�r���"��0��C��X����UKfK�,�� B���P���}@V���,�&1e�P#p��d9�[()2��.5�� �j�<����x`%��ZXs
&C�d���D��*@^ͥ��L>�P%,���E�R ���ۻo��g�o�_�I>�sH���Լmҳ�K�SV��L ���v�M����7Έ��ui���&�������I�Ң��0jP}ya(y�rh*5�o�]��zNZ_ h�o �SZoZ������٤h�@!*�,̜�~�)?��&�W���):��9�8�.�ɾȵ��2��L�I@��?t�f�"���TB������R#��b��K\ߡ�� I!{�S�Ծ�M�e��p�Z��7�Ӹ�C>��� ���'5�` � " ��^w@���F�^$�TJ@T �Z9D(�Q(��ƮL]�#����"�°B�&�^�64=3C� ���J��	��Q�)�J�K>ж=�{��w�Ƨ�3C�#�
��������C��FW���N�2�Ib=c&��:��v���6�_5�*�������;'�=H({�J`�Sis<_�d�D��P��(�1>� e>�8��@���ۑ��eq��*ك>��4�y,C.@ 0���{"�TR�<w��:�����:"�(���An��lQ~���;�#��6��)4W�n@DK��%�@�~�8�I#Ls���y�M1ՙ3ӳ���&�s��H����U1%�䍾\�\�I�c0K��\Ư$e�C�Lt(�:|:�q.��P�~F��{�3st.CF���g���t��ew��OD�C$7�oԹ�@�2,�3�D8]�ؠ�Q��66��O$dR[v�%<L>���T���/*�`@7b�B+�p&���ÿi�o���Ԥ���R���ǧ9�M:�@-}�*��)e�~��'�kT����7Q*�f�#���'����|~�{��3�D.�(�lgϜ"�$��T
4��C�c����B�E�3չ�H;D�9����Lr�)7@%,�u��������ܟ3iŧ�+����8��	5�ޠO*WP=pHyS�Oy@��H�J�)����t�i�Є�r�w���ʈ(&�'�V� ����KX���HI.�W�"��A�a%!⑥0�܊kFQ(zވ��=)\I%�H�#���)eEd�� ��T�[����������MڤM��L�I) ������OڤMڤMڤMڤ���[9���L�6?;��Mפ�Q;C$H� `W�X�S՗-9C1W! �)1�3��B�
@pB�?5E�P���t X�L6D�,`4U�9�p��H��x � ��T@<�S�ht)�u�T�� ���<���g$A��=Ů��1+�K��H�A-�v[�Lψ�13� H�갆�Xe�K(s����e�'���IL��{"+��͹v6�~gfG���-g!+	�[�<���U�cQ��:�p�p-g�:9���S٩ n��ΊPr�TB�݌E,���ֲ%(S*/��;�XŸ��q���\K�ʸvF~օ���؆�A�5FI�$��(��v;��&5lgj��A[�+�$�$J���dvhE��|%�o)�d
n#3��<��E�YQ��T٘��e�dϮB��6cܚ�6����%�aE�uc�3��:��9�8H�����ȉ� * r���Y�ju9���T��C@+2Ϩ�<�r��Q"2d��'1�����,u� 5���G�}�IA�L�K{�#���V*��`���<���<�[SW������4�� �<��C��YW��m�ȸ&���i�y�$���g�ɻA�_g
��b��zV��ئh6�T�����`�Ξ9+.]\��|��_C�D��&&��Z2d(*�|����xE 6g�R��Η��#G�?PY�k�O�Y� 7T3��7\K�J`�vz��F�9^�`e����F�A,x���X��\o��m�<�����I速SK�U��
�#0$gE�Tzl�"�`}����S]c�8v���U��tW�T�F�A|T�W �]�}�� �C��"B�!���ɷ�����	`������D��R��%^�
|��C��Oj�_� ()e���� �)�@ p�+5
��b�0T�j�� �R�񚨂�Ɗ-���J����̸>Օ��ڨ�ö �RՆN�
L��U(��Rۥ����&�J�ðY��?�7����L�*�o+����1�~�}D&��룻���u(�Jq�P�*�	TXj�4GiD���� /�k�JB�Ʈ�&��KEf�d?"��kh�S�Trз���,���g�
0����N�%��Q��H�k~��W�.\����s��;�&=�A����'߈�'��O7��+��c��uM^,D�k��s�K�fW&6�G����s�}{	d��G&�%m��S��:I�hO&���5�{��$DL�|[�ͦuJe<&��������� ����S�C�;�����Ҫ�>M
�ݮ��EcY|��щ�e	����9��(GQ��́����ʆ�"$འ=kϊg�M�L�Ag1R�p:�PY�3��r�����|�o�����`����?�)^����̥�!��Q$�R���l�$V��t&rYU�F�Y\:�%�%.���y:�"��Rd��9��C�0�D&�܁�:�R(s����Ӟ��L��_~��/8��<ʽA�m�S+��o�2Km�B�⌱�
�:�j��zy6�و�
Hq+�˥�h����I��3vF%8��A���3�w�ȼW���D��H�7�ڪ��~"-ƴ�^�Xy�6Y-�`B�i����u�J!h���DgȜ	��m��w.%��i��Me�(Ã���9m��)J���� �	�X�߆��B�"D�r�(+��I�� jl�!��B��<��
��X����D�y]��dZ�,忋R;�I��I��I��o?1��MڤMڤMڤMڤMڤ��m�儚��F�L�t0M��1vP(�N�Lò
�1��Z�;s3Ӕ��"YҀ� �((��@�L&(r�VE�d�61�  ��\{S
ȣ�%�몬4<�����HDqDD  y�Y�Z�I��]�jtr������@�*cӥ )�����$}������h A�Q�@��W:���組�Ƨ�� ��!��-Q�T�$+�hQ��3☂w�~���)qǵXs�|��Z֜�ɬ
R2����
�����E���DR5%���[�wd��V�tR��L�.�U��P�<��Ⱦ�U֜��� � K�R &=�Њ��6g[
�T6�`���9���u���ԵT�g���-����2i�u�Êp�Y���X��Z��b�E�&�'>t�8k���2d!�
p����r�\�$������]Vպ�,)[
���� ~6[u1;3˵�Ȉ`/װ-T�e����h�IF��3��6-�Qzu� �҂�W ǶRQ��@�@v$��Rj$�Q"�aDc��䠃�B�p�HGeYI���*m\� +�@��e������5�L�����M��	���Au�-&����RĢ�ޠ�<)he�i���%�K&HDQJ�r�d�P&|�q��Lɴ�h�O�B�s�(���gs�?�MA�����"ɖ0^i��|J�k��I&Or~ u9�m?9�+�J"Ma�m���q0c �0?Dܑ����eF���i�?O�&�i�O1�x�p��75Ceȣ�����+�A�j�iޑa�������d(z�Bժ��ڦ���1n�+�R� ��%�~Ԭ)i{�))h��[��Uh82�K�U8�dΊ#�'"xO�q)�/��x �!�cOp9; #��T2�.T &e�(kB�%���ZƤ���';1����R&,�.A� ��I�����B�M�l��i�)C��{��|9A���&����cR�!��/#k�c�Ka��7ۼc��Л�,�%^@4���E�K�ؖʘu�����#����I�'�h��υ=+����2��WE��$�
.q��	 ��@��|=�)�|s�vJ>�d��|�	'4T��VB�l�8��P�?kԛ��2��h�H�Q��a�Y��7�^���]����HG?�J���C:8�� �6������z�����<|�dD�G�	��Z��s3��E�*O��Dk%K��Mq��q�����kʨ�J�HM /��Dg�T)
�=̘ࡉ�Ee��X��Q�3���	���7Ԣ��?rR'ʨ|��+�"�|6�jP `T~������t�s9k�H\J�}aaNt{Ȩ�	�I
���F �;P�J��@��+p�3�Y�b,��A{�4�٬��p�h�ި�s�LMJSr�Ln�7j��$&߁������`��.��+ңIZ"��q����vK���*��s��ߙk�b��%��̊��E,5��y3����n��"܈jO4�>���Vd 9$*�s�{0l&�b����r9'Q1���>0 �	]R��7�aI�`��5'E�ϗ�7�I���YA�W.���Ύ��n�U��_��:�V��M�4���}�"�J�����@}�W�_���?�J2�JijT��U9� u2��qq~��A� �h(}�e���c�������J~��0��TD	�E\�ƪ�"kX�m�y�O^5gƃVe��I��I����6! LڤMڤMڤMڤMڤ�j��/� ����9�*��Tr�e��`����
����2�X^ԡZ��"X��Qv�!�*|-�Qm�\|�YR��^�3PH4<G���i��)�l*/���� ��p(v�;"��0H"!���n@D!�>VҟB��gG������l�.g�2x`R��~������ǆ6��ll�G0@�i��PS���m��L�C���/v�;$q�L�u�G#�\��D�`	
�S���EY��#�5q�����,����/�m�@��뾲*��R��(�H"ΘS"��(�Ww:6K����}��A; ����b����&�ls,�mm�`F27r9�FEDaৠ��Jdc" ��9H�Z�@$-���&g
�=�[۸�y�lO ��V�8؛�.��VI�\~^`�J�ݥ��Ib_Ρ�/�#i� ���F�2S�eS)�
��O�KRXJ� X�T:�
#����2)�e������2x�u�D���Y�|"�N���P&��AK��20������4�G;�.e�SfaT;�n%���Y�B%!���Y-u����R(r��^{�]����سk��{e4O�R�Lw���u��;�f,vթ$�!����W �m9f����0�H~[$���PVXX\�n�2��r0@+��q�_��3��,��.�`<$Ǘ��H"���k�o (�%l�\����C.*�R&]SҸ� �-��=�$�҇a�Y�G�<vT�ϒ���D�A]��m/��-�j��}�.sP(�=Vs`� �x�P ���Wd�)I�sQ"M�m��T
�g@*=g��-�� x�rn�>��K5�!n��;lm0����o;;�Dj Hn�1٠RuƱ�l%`R�ئ����Bo! �0�R�e�2�	�LD�?@T��-'���ܠ��A@R5�KZ%�~��-��,�+�s�7 `x�y�!��1	@���9�����RL"��j���e�� �a@{ �(�za)�TՕ.M&paR�aV���c4Tg��$��,ٍF�� �͂$�Q7~(��vw[���Q�Y�'��D�bR�Q�/W�	�25��T�BVj��D2�LhMN��!���V'"ҜiUg
}���`�,r>K�2jr��@�eW"��J����I߳-�+=�/A��҈�-ylZdG��T�ړǍ�R4�|��H���綧;�(�@-�0�[�"Jc��X.\�rJL�
HQcRI���"�%|��7�XD�P��mD�09K�Q���ر�b0���ؗ~g�^��� dE���TAǻ�e�/
���H�Hy j���x��9)~G�*�`�={��}1��[�T'�J��hFIuB��� �HsY�$H��%��P����O��W�D\� ��I�D�O̒�kh�&u����"�Ec�
��X�DBm�������L��q��	�uE"�[�LMj��'�D�����< �������lۨ[���T�e[pn�j��̜�t�"�T�]ՙP�4AX��f�gmA�
~�F��r��d�þ0/#9w�9"?�=f8P�-���X�E�Vq���<�k��1=��0�L?��`�X��+(s��J;Н�/s���^]�<c�rXj��.�
��y�%�h>��a�Jux��Hp�m/@���<@L#�T�����# ��
jD,,�̈�ox>�R�1A��ߓ:�Ҍ��J��,�=4T	4��τZ�r*����a+rҫ�����6i�6i?SmB ��I��I��I��I��I��.^�X�?-̢�Hg���9c�P kYV��b<e�%s���L�P�z��}��dpA?�`怟� �
��Be%!K�Ų�$c	J�LKe�BRY����,P |��P�!�pv7�	@�"�n
�q��_�V7�gRf>�׹����<�$u]�ʔC�p��g2�o:�Mg#R�o+�{�ܦ!*	zCe���
c���33���B@��Ԇ����nO4M�I� ��?��)C$STu��0��e�Y�`����<�g�P��L�L0�,I̵{��@ ��@g���E4�*�Hwx!e~n���_]]%��_�� 7�kU�`9�#�,5���L�E���}q=��&↜7����j(��Z)UD[���&��9���ȼ&�p�!KR�o0	[��{5��c�D\[Y���5�s��AN�଼�DsU0Ye_�3T}`�kh���7� p��xL�Ϊ���R��r9���Q4b �.)p�6k1�Ae|���b4���`IǠk�6�Ekc��	`@l ����fK�$ٕ���K�ǖ{e-Y��@A�|�)�R��
�O�>8hz���\c��6�9�^3���Ȯ̈pwSիW5�,���$3��V��غ2��Q7�2������xF�c Sg��(Y�:�TΩ� �qHҐ��(�Y�P�gZc���fB�)�T���Q>
^�$�Z^�?������ֲpJ෌��m��S��Rh�Tm�����:݉%P�X��@L I/^�_|��,AĈ?�u�?����������/c\�TOVkj�Ͷ
��w���k[�-ǀ��"�m��o���#I (+�l**�a��8u2�ۻ�?��+ɩ�?TGz|�L���
�<��2��˦=mͅ� 7��C��HM��@^�����5ܧ�5|�Ğ8�(����2�\�����r$#�� ]�wW�n�qtδ�M8 ��V'�3����-,��5���x�JkQ�5�9��+�2��ʩ�����h�r�7����_P}<�'��x�C�*�Z�9�Aw9Dm�`���H�Z����ׯÓ����9�C�$�4�K�c,�Ǚj��Z��,U�'��0F�̒,��->����gO.��{^ܾ�}0��=��1�׭��v�C𜭼E@����ü|jݣ�܊�NIV���m�tG��G��Tggxe���B'��g�V:w��dE�
��$�k��gO��_}��}����9	��񵁁V*	��o�Y�?$VG^�%$���Q�����x�f(�{ ���>=:@0;~Z�l�>��cޢ�HO�,�Qp���B��Tﯞ?���!p�|\���]\�xx�C�\�Eǜ�����'�t��}]��H6�OO�����"js� a�ܟ��O��C�_�c���UP���g 8<�{����7��+��\�1F	���%I� �N�R���D)�y���+�Wӭ�no�-�A�܉}�?�'�i�$F�y�#�E�v�?�g�wq�}8ؾ!��!�ᜠ�3�B0�8âTb%�ߋ�����;��oM�X&���:�A#�$HL���@뇦./�� ^
���D�+�S��|�e��v������}�{xb{�9L�t�ƈ��^a�t�Y ��������!�|UM��!���y� �
�z� 5sY�ڏ����}���r4����)�%����&R�'���VrEgq���C�`�mX6�H%nXB#���/�}B�b�&�����<���Y���|n.i����:��Y�cW�}|��L��І6���L�@ �І6��mhC��~Bm�ߧI� poӦi���@��^��ޤ��L� �� ��w(�s�/7ǟHB�SN�܄6�upQ7?� p�P��78_k���.3�
��B54��i�yd�m�g�6��+0Б���AwYl�J�l�qAH������%%^�:�� *Ra�)IB��{\
�Wf^�Ƽ<ą�1��9���g2��W_��7W����T��l��&��ק�E�l߃]�	��m7/Iuы�c��~�����վM��V,$fg/�����Uݽ/�c�`/;){���   ��qA0�e|�wo߱_$D�������Odq+ey�Z�S�������:��q��WM��5��H�R� wj���� ����n�`�2]����5���܈)�  ����@����ٮ2F;"C�Ҷ^�qK����@��;�ߑ��p[���5��i�R��=�Tʅ�b/t��V֪�����^�+ד�.�U�jݫ�S�𽾒*��ba��Z�pL�\C�~[h$�YB'�U�z�,EA� 8���/�qፋr���� G�I�سZ��~�����}x����r�'Y�G��i۳�3��<�q �8�" T۰n�j�����K��������Y|_�����@5 � -x��4�M3��j�✠$Pi� ޠ���,񑗽<�7_����Ϻqf����������|>g,���#Fw!�R��)���r���q�5x����D0XƟ̔�R�7�IF��J��,EQ+Fj�2��Т�X�n4�+��� ��e��4�5���/�=/.��ݭ�±� >3�k�F�F����fs��y ���) �P��#��$�s��
Z�T��l5V��~��qUz&xn��}���cx�3q�9J�pq^�x��9`��5�Y�����C�3�\c�c\�%���9A�#�S�7`�t ����!-� �56�<J0/b,�����z�Ŕ���Z�\�$K�}/$��?#^�Ͽ���}|�{��q����^z��T�)m���-}j�<׆㸧����?i�@�c�IN������k9)i	�N��� ���xZ�rE�Y�"�Y̝ϞТ���"�:b�H%���9����;K0+�Yf'�& [�_<��� u�1W T�$j�W�s�z�^_�g�9g�ׯ�?~
u>bN�>R[r�g1/�Y0�����}�/����q��ĺ�u՝��&���d<�U�Q^��	�����3aAh؁Hck��d�����}�e"
a�F�)��XF"I,�K� 0��_��7�%�`�c�� T��:a��I]�1aK�\8苗��=���$��泑�T��t"��E�ԱO=>>rθ'�,V�;�%����xQ)1�Kmg�m|��Vk�˘q&��/�$��:W�����.�sʱj�c��noo���г�oΠ��Qy=1�1��[�� y��5Դ����3unN$i�r{	�V���5VJ��$:=Ɨ.$�8�9I�S�τ}�K��@S��Nb��F��.<9��!���"L�=.�00�E�.�������� �5���r\� a����0F��Y1�+
�uX�������-�3�+��wx�����1�(�J�� �mhC�Ϩ��mhC�І6���'��4� ��Ǣp����u����v�| �vWD��R��&LF
��I����+@4�=�`S�c*�T�V�n���_�������1R�?6 ف̚Г �mb2H�/��	������9�,(�R���ZMX�Ǡt��W��KF���es. ��7���:���Ւ��&q���񞸠|��Yi{��<�-e�]����2jzEuk�:ޞ�R
}@ �p\��Rl�����-��Yb��T�6G�@/+W��x�*0؎��4pU+@^�!�h�rwċu.���$
��`T� {]w.�s��@9�*-2)�41��k8�U"5�gbC��uv��˺
SkF���sT�ژ:Ȟ��p�����Ç�tp��/����ShL�>�礍Ή�I�H��fm�/ ����B�u%(X�>7׌ĝ Z�磜�	�FB���j�k?���`����t��� ��"��� ?4f��ߝ� RI��Iu��Z���� �^��<�̐H5���ԇL�f\��{�d�����H8�s��v��ť8��|��m���9(ą=�l9��  ��X,©)��mzW�ĉE���!�N���p4��3�K�U-�a-��� n*�C��Z�@Dp� K�PLF| �O ���E�PN�8?#�����)K��Y�A�z�I�}�l��rTc��&5���|�5�i e�!�;����T��y�oM�?������d�xI��$U5��*�+��!�  l�I��0�� X��?��m�7�p��$�'[��BZ7��Ϗ��8�R4X{��]ɞty�k��3 �q�nr�M�:<0�:y�fY�Z	��o���|+P $�O�J��5 W�`��D�n-��p���"%�����O�.�3&�2����Q/=�-�'��1�u��j�<�,�E:�:�'r<�,`�*�^�^����͕��Q~TimOP�6�*�0��	�N��D,�s�o0��r��d�>�����5��J ��2�k��lo.,7y�w+bA@���8w�����:Ywq)����^[>3B���HX_O�.³��������*��$�����=Fc�Ǡ�GA���Yuu~�w~�<MIv ��Ķ�*���������7���+���T���9v�<�t{���^��I{AF�	��8�`}��9a_�=�j���b��7o8O �}_Ř O����s��S��XS��A�&�J��A��n2:1a/�!�!r̹CD(�3lp"G�\I�<��	H�*�!w&���H��JҠ��'W�W�lUVg:=�1����J z�E���^O$��#�<7��I_~�r���^c����A���W����[O6S!���n1n%��/m�v�|��PbĉM���8A'���I���=VO��kg�a��Y�c�?�g�q�g��J�Ϫ(Iω��Y�lgd�	����Ew���؄�	p��BۥЦ+������ǒ8"��g��s�Vq�B��K9�_7��J�-j�<�d�tВ(f��L�	��X��|�y�Y��$J����r�2��@�k<WT{ƞ�N�rp=��s9����І6�����@ �І6��mhC��~B-�ʴm���M-�}WU�@�ʚ�_���0�A;���n"2sUc�w6�l��Pr&���/�����O$n/�X`j��Г�~�E~nʠ4����~�vQ�*��u�vpk_�
�m�q�{d����~8p�
u�c�Ђ5�J���q9�C�^����>��.PٮP���\����E..��l�Y�v`5��ԹL��N�"[H�����	  :�??O
�uf�=/qY��x|.�Bh
:I��>S�+4�uGY��R��K]��w�iE7#��	 �s����L��� ��.�@P�d�D���űR>{�@�կ�.���"�05|ӪNm]�]|Rm��Ĺ��K�ީ�3�k�5�>ש �	 �l��}M5l�uMqh
�,��RI�����"q̸��)_����.d��6��Q>��/@e\z�b�XQ��+ �����n�����5Ǎ��i�h���Q��>��n�� EG�HD0��&g���Y�Z�{���iZ�g� z�� �#�$���!L�t<"�ٮ	�a�8)�� �6�  \��
]14�e2~��	��ƸM�g�ں5ſ���n���Qٓ�X�]�_p-U,[ �Ş1�ޔ��o�sQ�NP�{�C����<<�|��b��@'�T���!$z(I�7�#˙�c�6W �4L>�@�����&�	�
��|�f�15��@u)��X�0�}q�x&E�ٳ�V?���o߆��;���h�]���˄6�P?r�(ڠ2�" �;��O�W���o���
&`MT��`�ܑ ��x6F�Y�%�8���%���r<r�TO�����u5�As}hE�B�suD�ޙ� �7�L��w�����7./+�z�I�Ӫ��b�����8?=??ȓ���2���8�>lП?
|�9�5p=A����;ە����3�r���g� /��#��O��â���1�Vu�i4n��u�]A5��J���.$8�u���s���~N ��i�����]̣P����?'�,j������	��d��ߵ)��*t��p{�$٘�xj���`k{����Q���6��� ���>��W_�u�C�Q9s�|��F �a��8����×߼	�ł�G��b�G�Z���AOXa���*�z�Z�E�@�)���x���:a6���3�e�H<p��su:�.	��2�ѿ����}�:|��$T�y�--�qA�*�|�!������{4H��Q 2!�lc玎'���$ɬt[�����јۍb���;��FgW�2�1a���~vrƵ���j�.���?��_p_���7<��$�R\��x���=l��Ӂλ)�8�:�ӡuw��1��Z�����
 m����ut��<�R$Ff���)�9�(*M����ϼ��Z�8�������\$�Fn	��K���?��.4�Ӻ&aB}B�H��=�4op@����bo0� t������#���h{cjg��8c�8�U!�]���$&��eE���DD*�(ʸ_��8j�`�^�t����D�A����~�y<9;	��g��#�����I룟c�Mш%��B����mhC���ն� 0��mhC�І6�����v��R�ēw�e��*H5��ܴ��/65�h Sd��#��k�w�M��P�Ჹ��Ƽ��Ey"�L)cS�Ii�`+�O*����4\��2;a�\�S�:�--�k������k�����f݅;��P��L� i�6��- ���' q^.&T�9�S���������Է�
��u���Ы��������Z�!å�>�)ɉ�z%��նvy.�(���hB\\���i*`�6K��T���aGGYhV���9�7(�,C�[C�U6aUo����T��vl���$*��J��y^�"`0m��u��>���!��t�\��OU[555n��������*� ��tk�c�J�Zq�����ۊ�� ����l6�=AI CP��fuO��j�f����7�a�J`��E�8M����ň,�� U1.�i���i ��ON��?|�d2"� +�,��\�+DX�|�<�Z���������PM'�  r��2��MRƁϳ/O�uO����N089�w1��X��i�N���ň#<N�����S��Ֆ����s) :V�o(-q4=��}>_�ˇ��������E8O-���:���!�}����g���ʓ&x��h�� �nG�< �+9�xɉz_��/r�8���_��U��y��ڗ$`a������{��/��pHAy�6@!�צ�@�ǀ�����yՁ�e\����N ���0)��j��$B"���~f�>�s\�R#��,�O�s��b��BD�MIr������[E���9N��CX/7���}X,��#w�ȍ!�{TRC_��Y%1l\���\��{F����Ϭ^��3-թp�O�v�}-�70�*5	Έ��5�gnI�&>>6r�IX.�]��ݫ�*�U'R��Oǟ�#F�� µ���cw�p��/h˲R�#g�@�Kv��f��!��Q���E��/R�j�:�G(�������O�C*��@X�}��7 �7�{^�Ŝ��a�g��Py AUV{����D)�A�	�������ȁ#)k�T
	Q�l�9�(c�'��������|���x��d��F9�js�m�3�q��(͑o�7�lD�.�f�L�M����Db�f����xje��;��e��L�ë����t�q�aݟƼ�+��8W��6�NN�|V"����o�^�a�dG�� D�q`��/��Tn�@�ڹso�]cR����?�����Gqxe�7������*���s��kp�=6�����J.C"���3�i�دۛ�K	�,�ɉd+�nQ)�H\y���Ǐ�;�W Tu��zĳ��&����" ;RY��2�[��p���.�� �l~吢�}��#�Ӱ���%���$1�7���0���������q<��� rg�Vtk�LĖ��<�d,!.u6>��b9�@�[���������7���g�6����LG 3�s����&$y���9ϳV�(��4�4�9�G��pr~��qR H/M#�.�IV-BLS��D�=g�.�J�\��g�����(��P�u�Ag�`k�	�{��~GI�qGV��T�3�>���#+�UBuogY�����$R`��xhS�;)'�{���>P��3��G1��5O�����D�1�I��lUc��(W1�T��Y��n���́�I��j�w; �M.mhC��~m  mhC�І6��mh?��Hs��9Y�7mga/U�淦.o��Uuua+@�J�ɘ�g1r����^���K*Ƌ�2K�L6�|�Wj���D�������nhM�]SS�-�PCeVI@���!��1����sYZU�(�S򥦼��-\�Sq?��,.������)�F!a�	� 7{gn,K �Q�5�߾W7�@���s�v���~�f���m�e��Z�E�[m�ЁU�[�J��t��K���^W��j(���%)���� BWǘ��$ d����X\����Rc5T��YE�#�\�>��RmXBge1��k��S���B'��껢���ëH)ZhS������4ɭ�8�����	/�1��Wԃ�l���ј`)��߾}Ke��}Y����xM��� ��TV� i���!�]j3曔�д�7���Mj��6=��!5�13����K��1/��q�]i�ⲕ�8g�0?:9&qf��|F�����ϵ�a ` `��1(�``k�Z\�Lr��ŷ³�T,��y�iU��GR^h�nn��`��ĈFM8;=�^~����w��oU_��DT���fzK�
.�1� �,/!�Gj�}k�M�L�t%=h�g�����8� R� p_��|v+��r�0䮳���5�뚟��/ބ7o���-  �(�?���� �a��X�Zs��?����
Q� #V��*��$���W �`�H���u��C���$��cs$�:�K�'�J��`�XkK<�B �7�&qͮ�uءθ�px��)�%���V�>~� c��R=Z���6�W����ru�;�柺����;kb��aYޣ�[	���n��z�T�̋�(/0j��t6(��u3�W��E��U$�<����S>X����Km��g<�,1����R}۷�$�x���{�����s{貖��-b䗣�1�F�I�[���AAnZ�����PIfc+7C+�k9N1��g�Ս��L�����p<�m�^n�@%�j皐Xۼ�\\�:��D�^���E)������9�Yɔ�ׂ�R ���h�G}�Ol\��bl+��4T�<�.y?���g�R����@d9�ȱ��!��} c�0�1�@m<5�J{��4�]K3�e�9U�8g�d��/���ǰ+w|��_|E�W���א�vke����wO-��xv<���|�%�Gf.��Z���}�$�D:�Z�͎x�L͹b:>�3�b�#J6b��9��r8�b9�V{����O��g�I܄��-�~vda�{K�T���� a�0w'M�m��b3�2���Ϋ"N���cEP6e)p��rrι|�򫰯�0nS�+��d<��ec�0�)�V?���!�_\�=��'�o#�⺎�Ób�����u��6� �&���I ����q⢕4
�g@X��mT�g"�Vv�G?0ǾǨLV�gg�ͷ߆Y��I̧T��z�e�r����4�Ϻ�_�ʜ�df'�*[�sf�X�<M�|Kc񜘫V��qm��A�x�;�������r�@�������",�K:4�8��판IW�'�=gjg�D���w�J���rt��/����w�װ�"��%h�<�K8<L��}�,'\�{'��i��g%\|-�����mhC���� 0��mhC�І6������_�KN���*Z�=�㗀���QX3�SK)��"({ 2R����2^(�r*3�5�QM��T���J�=�vu���2�]���� �`�0��]}U�;`Q����j��7 �
cu����vit�x�Yê;�B�����O\�N��σ��NP�@���F�F����]�#� u x�v��KJ�]������6�>?�u��n>]�ޚۃ����%X�g&8���:��w������UAbL�����.r1��u����wf��^��s`;`�C�,�{���܀ks�p�o��o�_N�R�.�y�oe��gu��;g:Q��<�L��&;1�֌��^F!�;.�Q��kQ����2,��ج3��5��q�
���֓�-���.��/�`��,�u��ÔB1��ђ㽯U+� P�Bϖ�<�E�
w���+Z��-/����.J�R
�Tc����m��f���tI��P�:����D$���Y��(�F>HB�}�~���A6�x.�x+>.�N5�C�������x	�| �T��D� 	1�h5b 4Z���Q��@Ū��:�H� �kR�@+  hu�[��^�L%o� �ԀJ��))���-:��ɓ����"��ޒ8�A)��J4 ����@�֬�Vx���N�j{�����ﾦX�!��ܹ��N2�b�}0��zE�A�kb'�`=`��O� ���O�]�>r~ �\�nHl�q99>�Cr(��^~��m{�w��6!�sp��U�x�Zf���t&�'8�2���T�T����L� ��nc.�ƈ/F�C��	c�+����_�l�H�R񋼉��q�ej|n��>�|N��u'07�3 @~�2�1�9�w�uXĹ�=�{��[��(��xj����L�>�נH3˛���?}�7�Y�!W�Ƕ:�;�MD�Q0t�O0e�Kt��Ī�S[�����HP��%-�������*sp�
��]�0����n~/�R&b��1%����14�T�H�jg��ǮĆ�%3�4����IڟtV�:�
�MyVHYA� i%��,	���_He���sv�������Ua�\�}� �"�Q��վ�5U[\9H*���jv3���^���s��)>�.#p$
� �&�a���s�}y��c�ӫ����W����ߑ,uRDk�4�M��F�~b��r���5�B| ������☪���בh#�yC�9J��k/	_�������,�2�)��ٷ7��W|�ͺ�C�X��O�E�K<��w��}��7$����s?����!\��+Jgg'ܛ˴�}H��vP��6��_U�}�N,F~j��k����81�k�rTERL ������q���\<p���]��q���<_-7|��c~&~'@�ͦv.�3t�qH��H��%%�$4��j�7�
�����l�$\'�����y��!'3�9s7�e�5�kH�{X*�'~����.�۩�d��q���{���e�쯪�s�����(D���K��{X�f4U��h*<���w�pNr�:�iC�0�6��mh?�6 �6��mhC�І6��Xk۔��_V��uգ]h5���^(������t�u
�Z
[\F�/�������¼
U�����H�����y  XQ�����.� �n6$
�2$�v�~x��y���l۫�q��d�]*'T������SBqV��ԥ[�f�_҅>�}�S���g��3����&�{�9K+�nM����"���tEW��Ԁ*�����쮹v��΍��6�����U�jo�=g���=j�m�KSat9�ZMݼ���P�B��T�>]?��W�^Q�S�`@ tQ�x$�!�&ρB�� `չW��� G=�^=0e�^�� Ǽ�Á.���ą)@���F����puy���	B T�PN��@s�t�0����D�� �6�b� .	��9;X�^�}uź[�?<�Yי�Q�gY�8��	�^x2�F�A� ��v@D����a-��9:d�K��cβ��fc�9��U��o"Zs�9k0_4"��-�֦�#�CQ%u�y|.�� ��7`5ݘ�8�m�x�8��:�!����ɰ��^[������;���������`<�k�"�jkk6�̄��%>J��/�M��#xO6R��Dp2I2F  �Km�!�)��� g�x#3r*RQ�(�>�g�0d�|�5���/� �S����C.p ��H>��o��s�'�\��D�V9 Ԏc���1����R{HFe;�. n	A�9IE�9H>�e՝�u �2�5���fͱ�!�,W�����հG�į�#N8�f����X���@u'�`���KU5��~�G\7Y�XQ�欄[�|d�LD�9	^��v$Ye,k���r�c�pw���c���*c
�Q�_���bEk~�%���M��:$�9@u�Ӄ�'�c����:�>��k`����9���J��v=w*�mH�$ ���9' ��noi�/Uv����9>�C���1��>S	'�9��s1���=tnI��>$ġv}U�$������b�Z��T�H�MP�%�0���iK�i{�a�m&��w�T.2X�p�9:>������Φ�p z��c��y�rr��yq~0���*�\[�ۀ�TzF�)�"�R�+���g����~�'؍c�k~�9F
�B<�����y���W$�O��IZz�%lO�\�
n|>��ap��h��׃�,c���-����D�د�~�8��]������+�"��u��̸7����)	q�II7�~�3��9^r�%xk�����Q37�>x�����=r_�w��~���)�{����e�}�'�Z��H��� C>|��7����������������%'����9˪\_݄��}�b?�����0>\���_�*��E��*\�q a
��eݩ�v��|�;ț��.rR�;����-ʸ���O�A��s�D?�_�Jt;�|���	����
[�
�&�4��^�;�blI�Ğj$ܤI�2DNRQ>����ʴW��$��Sɡ1' �J�[k.q�@��-�g�ي������Y�;HȍX�X��k�+�}���	:>	�?���Nǌ�5H���F�TI�H*0W&��`N@��`D�����$q1��ғchC�І�����mhC�І6���'�����,ϲ6����,a�Ҙ�\��f�i!zAuj��N�Ki[����W��Bɯh���2��.S����סj���
e�/.����9�;.�*S�WsP���k�4@�ה�9�����.�5 ~�'���E!�r�1j������T?��n�����v�xV�	�Y�\__�g�H]��и`��ul�Pp�p)ZK�Wv��] ���v��G6%���/����xe�ek*`��.{2�����r/p�N���"���-��Yk�lh���AQHK�`PR�i�:&
��$�kNN&8�����Н��&��1����L�n�^P��d��vJ�Յ<��R��(�:�`V��}-� �Vq��?����������}\;���c2t��Fwk�y'l��Z'���̣��0bp�j�	^�����z��j��wo��;�t(}�����I����sSG���Lk*�ߨtAU�vIޫX]	z8Gn,�~�6��gjSW�M�N�p��H ��!�	m��M�ʒ`3K/ ���\ ��������~���tyE��8oШV{A�@l��e-p�1�9έ��4Μ�`�S[|�:��j���X#g�����}��,�:8H����,��XR�����J�GX�g�Ư����y��yC������tk�>�t��ٿ���%sU��� n�G�AQIZ����I��� ��H�9�QB�����q�ØS!�>��pa�v XbL�D��u�����Xg i�����͑�೾9����^��c�OF�5�mj�ݣ��(g~Ol##%�Y�W��?������9��1���{T��bbJ�ӱ�	?w��^o��l.��+��gˣ� 9q4��J���">�˸�8��(n��5���*>�aؑ��U(����o:}��:�`��-�����8߲�vb�>�����q������Jn�|��M_v��1O�\N�����;��WB�P�,E���f:��UK��>er�@I��sNfgfy�v�e@���f?ONg*�`.'�W88�b,���˝�n�3��l����y��qE����F�<�=GSNI���Z~��z�;G ���)؊�<�+~��p}wG��
nnn�z��2������R[�e���"Ϧ1�&������,����31��{!�T��\<��L663�Q�A:�`�R�ۋ[�)�%=&s���}R��\�X[&��T��]<S=��������s����n2���&�A�F	�	�� `�� =��7�|�rɳ��k���gOgs���ZNG~�JzW��C�U���Vb�Όʹ�S�����y`W��w�t���B����5���fI{��O�����|3��,�}����+�J !�����xcggϓ�X�x\�*�I����9͟���JV�${n�SL���&��*ŀ�C�GY�4���V����cW�cX���p³2��G����p����,���s=�tH<�:gz���Z =�·1�(>['��F"k�,��.~��ߕsr`�����iGxv��7<'��#��tzıq�{&��y�{q}�b���@h�%�=�#I+�w'&J��-y'��ݎ`�ӻ���X4�N����	`hC��~m  mhC�І6��mh?�6��h�<s��.�X����������M!�t����f����biJ�֬NS��s ��;�Ta�
�wԎ�� �a�U�v�K�U��e6.�@ � ,J �#R'�X���탬�K)���L^���8��j]��tu(-�Y��
ٶ�ţ+�d���@3���q�K>N���Es��>����
@놎Ga�a�X�ӓ� m̆6��ݎ�!.����&�ϲ:�*� ��/���c�KS(��,b�5�s�;a����)�YG�iz�v�d��1�<��2Ȧ�؍Tw����Q_���\�T��5�ֺ>P�6n6��~�k����k�ԕSAm��`c� Xl�:�L%2��/ S}T�h� B[<߄���pw�<yF�	��$o$R >�>,��Z����6�����Jx�}v���K� `�3� ��z�~��2�W���t!E-�q_	��J | �l7!1M����((1�L��	!��Ɍ�sP�a���>t������� �I�8�큂ƕfF2�z5�<��N��+���7����$�����m�3�b9$M���Aj��g��:�� ���� 8�n7��c���x||d*�J������ݢ�5� (PgS�צ� 8����V��>k�� ��2�hc��}=T���@�t6T�צh��c!5� �����$q�V����%Q@���	��� ^���K�&�59㰱fz�|��G�FtM�:�N��d��($d�V�E6�@i|rr�����	��T�~V�%��A�8ΏC�)�<YQ-!�MR�~/���u5�U=�)��
���s5m�+����>Trz9��pAE��Z�|.�Y�j�s�t$��.B� ��ac6�w���m㼤y�3C�a����w���y������{ڏ���?��9wq�kR��P=n%d\�{x[�4p����N]���6���Ś�T�NO��n�X�����1��{O� v�zUn%	A^�����/�bO�W ���+뫛$������఍��	@u�#Z��$%����6>��p1���Y����њ?��x,RL��<o�Ĳ��D�����{HI�Ri#�p~Q��|�j��}1�sIñM�b�/OIrl������8�K�=�XJ�k�;s�����F����4)_���]����s�(�]ل������3�}�	[O|��ȇ���?�D��޾}�����ŋpz6c�uX�OXk|�����'Z�/c�����ps}^�x�����x�&�<܆9l��f}���d���>2=[�1���M�e<Z�p������71v�iko��7�Ԅ|[u�왧�c'*Q2�I���m6�U���8P�X
��7o~��# a\���8\7(Ya?�U��HݢyV��q����y�/�yAx����W�L��Vܓ��g�iZ�$��ȗ_�O����!����-��������[:5���O�Oq޾��ux��7���1i��l�+	D�������t�8<��?��I�,I�-�����Cp~�Wt�iN%*P��_�D��Yg�I<�� y
g�Zw��~����?|���[:#`d�o�<���������1I*,��O�ܖ|<'�$��M��	r���|q/>���Q1����#G��	��Jh��o}����?>Q��Y���M
+3�o���nO2�8\��Uv.їP&�����rmNL�u�Ĉ:�9���2��mhC�9�� 0��mhC�І6���DZ�4� �I�f�O�:�V�= \���+ӂ�;	آY�A�*��(Nk\��f�-��*� {̪�C�]BUZ��ǥ< \���{�v��)m�Ё< n�>�eS�T;���-3��&!�@��l�Ë/�/�pY������x>����H d%�l�q�uS�FJWS�p) (��ܸH5@�@�����	�t���E$�} ���s������B�$����)��>�kI�l�4���n�Ju�
K` �^��=�:� q�:M�>*m�'���O����,�����s�-� �b��>@3]^B5�9��d��i]��Ūb�a]V�˛u��T��":3 ���5g�x����G^lڳ��a<8��]	0�u�)��8ϸ܅�k�Zu*@*�G����,fE�1�D��"1Le�)�N��/�ȭ�O�� +�?b)��-�Y�OO����<��TԶ�bR�W��;�8�Z�:^���k^��[�LU9�����	�;�%�CxA}SP�����;��M��<6�:1{сw�&R@㇠<>���v��E��R" d h�ǁ�h\�?{�<4{��>��ÃԜ���q�uxB��#��V��}89>�*�׉�F9�J��� 8��#�q����)5T�&��)���p��!����!F<�K�ْ�Y�o��2���,���_݆��1����p�?��z}ÚÚ��x�؄u�;J�#���oo���0.&$�����cA6�Zǵ�7/w��ߕ�}��n-f���jb=��rt��c�#�_�G!?*���={J�Lm��tz��=	X{xN(��RG�t�O �È����:ی9g_��t�u����8�5<�`�zv�I��kN�|�
m�����9	6qm�"��X����.�z�{��S���~�bȝ �S�n�^�� '� bd�b�|�d��uKq'��T��S�c�<����'{����YL���x �ǸNo�oH*�f�����Rsl��dY�H�k�2�K����4���zKr�2�MRẈt���p�0�p��ۀ��h�L�����V�;��v?Os�$�%:7l6[Z׷mb�R�C|~~A���<ȒD;�cW�� � ��P����c�3�k���(��8��<�dF�qb��H�Ls.����Bp}{�1����E0@\�5���<������ Q"_���ò(����O$��o������.��/^����"�$��r�u�o��oH2���?�W����|Eu<�m�؆�(@�U��8�e�'&��l�9�1"��pN��F�8���zC ~M������+3��O��$�t�g��as�YܣI6�ߛƹ�����y����Dy�60����$� O���|����D�N"b�> ��֎��_�| "@����0y9!)�;@q쵭�u�殄��G	��":96���gϸq�e��"���"�%t ���o�+����_|�c˵Ϻ���$,X��>'�ѡ��e����rTA��3�^�����eN�c�VZqA����,���F�"�gY��j�,����3G��X�cL�]r~>]^3�Á#M�����u��Y%3{K�m0RoO���y�D �� �g�����&�+Z��A�Pv��j�:DR�[q�W��M[\8���r ���i��R�\�!EVt�ƒJUe�����NXFGgO�W��=����̀�mhC�ϱ��mhC�І6���'�� hS\�5I�tŐ������;8�*k��ㅭYn�R޻�� G�Z�/���R`*-�ld-j P�A�R�ά�P��q)��e���E,�9M���,
 H��ڝ��T���v��X/LL�" ]���Oَg�K��w*���r߃|7ie�ܶk)�M�V\^�R��{X|CUP�� 9-��f:.e1&�4���R��W���R��r�=�X> ���@�?3�@C�"@4� wf늦��U�dz�Q6
U��ˋ�Կ�lv�"�TJ�U ��vE�_ f4�{^j��)�;�g��&.A��z|\RQ���h��1�v�]<ۥr�;̶��:к��p#�1s�%���P[�x�n�cEj�c��b_�k�����-j# ���-ͥ�nmLQ��=��%�dགྷ��u��J	��>�P�6T�Bi���6<���q��Ǻ��  i�	Uj-��O]ɞJm�} J~��Z�Ki9>
Ÿ�T�� ����c���	K���W	��T�^� 1 ղNWb�׻��f��p���}�A�']#���.�� @���d�B/ ".W\#[M���gϨą;�6w�h�C~��zJ�r�����L P8;���R����&�Ռ�EK޺6�r����ԉ2����a)�Y!+����% ^�����w|�
@.�`�~��9Ei��r�ʁ��� j1fq��`��^��2Ǒ.7�Y,��vǭ�PR!w�P��mH��`�l�9�&ƮV�<����gg\s �X.dvľaT�s �H�_�1\q�Yj#��.7bls�{dRde-�E�߹���V�q��U�S5iN	�YaNYX�k�]��>B���� �*T�bX����k ���bg�w�����q�\�a����n�p4;	Y)�w_
�b��΁�a��>���:��*�C2���;�h�P�g���rk�����	��q��b^�1aY�L�g����曒�뱾�Hh���X�}��X��z��#Ȏj^ �=B�;*���R����#NY��@*}c�V	���{����w�9D%a�1Ǭ��>6S�"q��ʐ��IB ���ιakd8���2�Ţs)�p,⾷VN�!x����v�^��H`*�B�r�_�6j�!�W�g�����}�����œp}w�|�W|�M�ۯ��E�������������.o8�Pտ}���,K@�8��ob�����ɛS�A\]]s�C�?�����&��b�^�8� k�16P6�.�|�.:R�&���tN!"��l�t$���A�/�����$�
����H>�k� xee�z�7�q6��u�9��?�S�x�qE�a�c�,�ށ=n��2�ԋ���z��fu)�H*��h�6�����[15��ag���{�=�'��VVf��V�o�>���2V�Α�f᫯�ƪ#y���^?���ND�IV���<��\�ӓS~�c�_H (�\��$0�Aa#�9)��Af䷤[�:'F�H���,�5��������	g�I���dG�>�a�r������#O������۱����+��@}OBo�Y�)=Xaş�y��S����{́���b�ϚnV�x"�z�0 ���@���2�YR
1[�,���-�`pdpR�k;��7
r'&���$Ϣl��,�3���)9}9�����T���&2�֥�� mhC��~nm  mhC�І6��mh?�&��IpU��r��~w������YW�ׯ�N��[\����k�� c�bn������]w0uJi ��T[��{Mͪ*A�����-.�����զo�4R@��ϗҪ��7R������0 h�]~N�1/�ȏ[Y���pI�<>O��� �p�3����5/da]�瑂(t�{Y��Gf1^�*c0&�rG�sZ2��6渨�v���va���*�e�� ��(�pO�́G'G�� ���TkϞ�|����?/+#�Te�B�ߊ���b>�)�js�!ğ��pG;�VJ> ӛ=L�9ەhC��CE�]S2&%H&T���uc�:��|��ψ���-�B�P��%���V�k�#V��@u^E�_�⿸Ȧb�T�K��EL�ʝ!�H�;E�wm�8�NH�-?�%
�l#Y�SR����|�1[�&l��̎��Pc�pwǿ�+��r �@����h�>yU##�Mu�	l�p� x�e)�~�J��+;֭��R��bĄ��)��Gj��3���z��W�W�(��r+��rG�2%��2�����W���N��qş�5��F��s��YX��d9�*��"��e<��=��+�A@7�~0���\H0����=p�%����� �1�<p}uNO�4�;�������7�$; >���G�mwP&?.I���2����U��Q����8|�]�ym��B��9붖3E2�X�n"uA��Z��N1�<	�v�{�!Ix���ph X���,�`��9���o���
0"�%m%��m=6{�.Y<]&�z��"���])��M��,�`�.7����y������X�MWuG6�`��؆��=�_v�I ��5l�I���	,����^�����a$���'��[�tA..�1�U�r%s=^�	L���ǽn�VMg W�nHZ�s�����;���*�pzvA�j����d~��@=�j��Hu�J�X���?�5�sDpBm��װ�b��ʊ���o�o�_�9��)�1\_݄��Y�j<�u�v��Z'�����LK:7����Iָ �. vؠ��[�.���YH
�z�s�<�$�	K���&�8���ۘĂ?��*�I�����߆��{��ӏt�i
6�7חv!�
��q�ݓ$tc��7���?|�Ioȋ���sL�����,�3g���� ����}��s���?���B�>z��������#n"���2�>�7|.�[ꌱ�<��� fd.�M�?��������p�I������7W�1��NH
XZy�=�o�	�A��-��/W���ć`��3�rZ�ƾ|G�^�2�ޣ6�wI7�pN���93�@�up�eXl�$ܷ�ip�����~��1��G��h��
�Ϻ�*�<��#�����׹�u�Ƥ�3�L�}�I�^n�#X��189��!\����t��ӟ�D���lU�8Q��]�rA�|b�UaƼD�Ϟ{�{�Ă̈�XOI�a�4ri�$�~�jh�B�@�(7��N��~��?�=0��7��8�_0�p`�yԭ��؏,�#	Ξ �L�&$P`O�+���td���j:�m��I�j������ׇ�O����6ѹ���gIwhC�І�����mhC�І6���'Ҿ��v�^�:.������0s`��V�9x�V����u���R"�*�d/�1�7^OW �����> 	46�*��,�`թ5q!_4z(��p ���.����#ֽ��5w�Hm��RQצ���\��ƳV��,d�XǞϴ�?;����=/�X�s�#`�ua�� *^��ԬP�� ��X���Љ)��Ƙl��Z�;(�	��ϥ��E�Ғ�B_O=x��T
���L* ��a����{~a�����t��0�RչꉵK�$��6�P��})�5�L@�+u ;����*QtI���2S��D?���e��uu	\w1�vX���kT+Y���M�t�:఍�M�lc��ဪ�,5W����m-�/.�Y�{TH��Py�yur]��� �Җ��c0� T)�]��&�[M�3R��'�_��F�Ae�� ����ڄǇ9���Ɓ
A�nK<�T������Y1��L�� ��s�ؠZ����K����:1�}�|�pr� Ȧ�w���p�D�D�c��ܽ­f�?��a�L����!�x��Z� �dS�5	 Pr�Y� ՞
Ȇ �v�!�&E��*Nk�>�	�XI �,)�P+�Cd8�<�>���.ޝ���ܶ�|"�+��g��~����l6�ky����h�>}�y�<|�eJP���>���Q9�X�R7��*��˫p{{D|!�����z����u1^����jG�5��)��Ԗ�����ZK�Q%���
$	�i�|��>������)�X�m��M8:9Q��l�w����s�E�A�`��5+�0�ߓ�0�	I���2�Kb���U�?�f#u�F�8�ݞ���Ё�i+7��,B�c��s6� b�fr�2�s8��"ώ�&a�- ^� ��
p|�Y��[�3q�u��ޏ�_vD��E������\��?ʙ��cr��xO*��'+[r�}O�M�C�u�O�T6kĐ3	��1A��l$ ���\"�B��t6�c��+��mQeT�x��'7|>H"�5:��5�u�_��My��J>�� Vh͵H���qyvI\U8 c4� J���g��$��H; dd)�Cd�=Aє�p�������*��A�x��`ة����S�ι9��"�In��g{��R�9��:���������➀3j���?�W����$�H�CR�',Qf�����ﰍs2����q.Qg�1����m��bs�N��:��?\".��7ks������B��%�|���0he,BkdQl�)�g�# ���r�/�/�{cgS�G����q����D"b��ݜt����} �>|O�|�ql��`��hmD$���`��k������N�3	�4V�#a.L�����t�����\F*E<��-�,9���C
��v��ҝ�\m�� q.����ɚ���p�8�o(����,pOw���z����A�ȉ�?Ƞ�7=�Ⱦ��Y�	8+%��/��E�-����\#��(�[�w����&\�=��w�އ�'��Ҟk�Ci�g�L8��Me�R*k����N��d�C��t�H�k�q�1��IN$�\���'�pӕ�I�~r��,�U��I����HX�xN�՚�p<�3~��{K��$��ڠ��U҂羚�ke$b��L���	S{�[�*��'����R#A��z�[���:ӊ�mhC�ϣ��mhC�І6���'�T 뤎���TU.Yr�Nw�z��W���v����TԶ��[X�vw�)LJgR,�15U��)�L)V�Ez����,��M�ef��:�����~�K?\4KU��]֓�2 �]��{�`
B���� ��"�;��)�aO*[{\R�� ,.U���1�j9xa�`[���r��:cŋ�V��ur@N�k�ga�^�����`9.qq��4w�|Gc��������̖���Ř+��a���s"�� �Y�WVUjZ�f�1�<z?C�ǪЯ�PVQ�n*��J$�B���w//p����2S�$�C�H9%��^��z"�-���|�Z�O?��'OyI{d�3.��< ���B �n��T{<�]�Rf���V��eg�J���c���R�HɿTVw`+As��t�� ��3�8� � �A���J�=��]=I�^�W�Ħy����
��Q�gZ5��E|ca̦3ߙ]4Ӳ>�@��rN5,-������rTh�4���^X������s��Eg���d��D�F��[�+�s�?%A�:T[�� �Ȭ�UG.�g���Hwڨ�)��s��5�p)��.�j��].�̛M���z胔j�]�<F�n�T��Q�/|D���j�g���b.?|��T���Q��wߓ�5���߇:.�*~���۰���q���t���*�p��(˱�[�֘�Kw���?ʈ��:t�GI+����}�} �#��9��Z���OTI����prrN��� (!A4�x�{�.��)�\
�8��7)R�'�܆�3I���r��,�83�T^���fr��q�����C*�{U.
�������*[�zk��R�4��4ۦ�E�5��%���N�����RWz�43{��s��<Ip��˂tē�����o���%:R���l�A(����M�� �S
	#;'b�ݳ�����_��1�,{Pr?C�e$@�b��V��5�^�-�D&+��u=�!��y�Z����d3��	��$�����<b}�� �u���W���.棣�Q��v��o�k������eGN��^�g��7�-������]�ֱ���d"u�ui�X�q2�� g�p��i��۷������:<��%9PZ��G*��������$����>� Vk��?Йc�͛o��?2W�c���o��gG�Yמ�����"����H%��}c�Z�l,Y:�%O��:��Y�T��a����Y�	|���q�~rD��P.?^q�c��6�J���3�����)�����l&RA��G�nc�)`�Q9�:֔*Q��/ۃE�5��Fa๫�	���*~�$�<�2N�7�I�}$�˫K���@0�Z��7<pϊ����9�~�����Oq����t���C�K�!����cӂ����\ѓ�h�+��՚�M�# ����8��~�0I钵g���g����qq��&q� ��9\|Y����+q~Y����'�yqΠ�_�t��(5`�����L�y�Q�y�I���YY	�l:f~C�.��T�d-������|�j8�"�(�=�9R)�T�0<k��pf�[J��.Z:z`�@�E�� 7��Zj���;���H�jl�S�"��'��3g���dhC�І�����mhC�І6���'̻֬��qɕ��w�c��ҋ�}VϺ��mt����xD;M(T��Nvf�]�C#i�L�T���ó�Xw��  8�^���S(`�Ֆ�<'`����s�jO�$L�}�L����Fn{���c��4K\y�v��PF={����e_
{i��@���S^�mx!���`j�^_^�F��ȼ�A�j���R*\��Pk�ۻ{��?������[�2�������	�T�}�/8��0E}�������0��5�`����n�	��ߨc�IR4B�Dc��5����% XLgG�5�8?'\<�<�Y���F��jr�>/@�W�RiYć�]�{�/���x[J}��C-�X#�� �V~��n�ɴ�k��[Rw��Hﾮ:�c���� Ȓ� ��h��8����, RS�C��4��X�� �V���
)��[�<�������V�v�����B��ʥw�۰�<b�ת]���.����1����m\��e�ג����8��S��~�,�r���W�_D�:i��Ǻ��&�v|zJ�m�TJ� �c?1�&qݮW+{.��8x�|L�2��;>Si�	��l[�/���O���9����V�ꂔ�i�hM)頷���ZWa��䋶0;���H(����Ix��?}z�� $`��:y�߅��}��J#�XϺ�[~���9���b��IQ_����	  NR�ʘ��������O���Rs��R}��r"ǳ�������.M�	�"�^]^�]���P|��s�ݡf��T�F�9G| ��3�9\��js��{*�5���nu����T� =H��$,�'@+K9����4����r�L��Uep��S�V-�ox�	�h�qJSG��2:�4�^ŹiT�Oɿ�����E�������d�\pxO�s��Z�G)�-��zֹ>��-?�jrX_Ӫ��=3p�6V�e{n��%��$�y��M����<�M��|���}���`A���;�Xo;g���<���� �h<�<RA��l�����,���G+�����5�Ȇ�1��/�ŜW��|I`}@N�XH���u�>���R�"ة�|m.0��a�<�mg����N�% ���׿�����ݻ᫯���������?�}p� %�:�1���G���W�(�9)���2~���M��Q�s��E6&yb������̥����?���_S�Q\ϫx>\m ����I���ʀj�j�/S��L�ޤ����8��P-y)���A�D~ Q���c�<99�b������������S�\���G�L�s����H�%��vF�a��8f8?|��c|wOr����+X%�35g��W�00��s��}�x�I���F�����c�q'p��:�t�����3��xP��8���ރ�����~��r뉯���q������?��8����rO1��P��_C��l�ھ��k�a%M���<S�:&�g��8Wj|�LR�"�Z������?��όM���'�������y����섳����<�ݧ'3!��T��my�������>�O�L��ʤ�1:�������cm���=��S�����ZFO8���[W�w���8�=�-�������C��&G����u�?�g3#ze|����ÜsK��yC.Zo�C#��s[�7i� �����-dhC�І�����mhC�І6���'ր���iۤi��S!5����~�W��_v��v*z|��f_�����p:;�%X����Wl����8�f��v ~fo���L��Pi��¬KQ?j-�� ��N�"����)��Giv�E=0���vci��VY�&5#.!*ߠJ�e>75�~���z&�"̡Z�e?�!(Q�8����	�qS��2.�g!��`o����έ�^F�S\����l�׫�.��KT��1�1��۾����nNN�i��F=�ׯ_s����6��:�z�j߁U���j�Z}HS:��И�;'�������-�p������7���sG��v��,�?B~�0��n�����oC����כp�cG��N5eJUT�(Ϻ����9�X|�-VR|��ښ�-ֆ��$I�e7�^p��*q�`*����9j8	� �� ��t@:�ax����X�îw2:�sr��#�%� �n��4,�	4��F`�A�^7�i��Q�o�/K]���059�WW����[���k9�����YZ	0�R�.�EgmJ7����ެW��J[YU{>�C�����R����~0���'À׀���nj���H��<Þj������"�����A�kWefL+b�7�c����R��Wn�P���B`��r�-�{��>��{�~d�ؖ6�;HF T�j���k͓�)B��هUB�1r���^?H,��~�a���Ϟ�}q�d
આ��HS��!��� �l����n�h�
�S��0�)���n��4Sr��wi�ysw�� ��)�;� �1���¾�����[��:&hv���N'5���U#�o�Lݲ$��
Hn
����1w5�t簕�Ú�v�^��w� @,Ԣ�y,`���iT���8h��ۑ��:s��c�hW�j��Ѭ��ك�o�PA�L��-j��t�@<72N�/��7�Z��UV��$x� @���.��I��4ޡ-��X_�	�w�p�*d���Y!�qW�-�x�˖�z
V
�}_��}���8LT�I�a��Q����G�狠��-m��,�����iC�MAO�Hy����C\�47F�(m���u���,�Lt'��r�;('MيqF>�����Ϲ+s������fq*�t���,����A�A������F��	���	�����T�xqyC�n�n%ꘂuv��@wӈ�A��
��g�X��(/>>n対��|��We~]˯~�[�o�e����˕�s�1ZJ���)y��*{�2��~��2o��5HfwT$����K�s�bn�Ə����_�ۯ��p�xr����A�����Ly�+�	kHʭ�N`�#N�]h�LU����� Ϡq�3*./#Ӛlv�G@0Y@�+�JN-ׁ[�P�i_���+�:��=����5���}��������Yh*��r��%�$1#sp�����rM��b�%s�H���5Ƣ~���k�O��r�3Zؿ~���$ĝ�4�ɑ��C�8c0���1�W���J�n����������u�rI�+��%&C5�y�x�X��Gw�Č�c�KhHI*�.2u�N ���X�|ԿG��㠤��q����{V�=��ٓ�J�\-�1�s�0А�Ԫ?3eӨq�������Ε��Q���꜄�h����n�����Q]4�᪌C�7,�:�q��A�]�hi�����Ĝ��"d�б@�A��J=�r�n��xU�9Gu'm�[2%��T$�3�N@�)c���;��(ȸӏ���)��HF ���J������;���e.s��-3`.s��\�2���e.s�j�M����,�P�Hs�B0.��G�O��dY.T���4�А���@���-���-m�SS����h�f&JX�OU���O5'9�p�������j(��c����JH̥����$?'�A�������r�#s���d�e�(C��cP7(0y T��3g|O�nŐ2����߫f�tVk��f/����W�t�-}�jU��O��!�4����Ѣ9h��{*�ݽ�?��w���������<�Q҄ɼ�����݀$�lI��? ��B@.��xX	�'�s����0z�%����-J�M���G�ߩ��ԃe��3%A���`8c81-r����{�~��1H�����.�+*��B���!<��8O���3��.�CRL�������rO$Wˉg_��4��	�L�51�`�������] �܇�,P�>�����������A�L ؚH:��f�nN�)��J� ��Ć�:88�n}0��P��s%9�!���I��tX������r��_�3\��$�dY߇>Y>�꼓��%4ϑ�7��F��V�S�f6�p�ۮ5f%w8T�U�F^����s�<�������J�X4��h�Tؚ� R9�rr�7�x(Ll>�{�9���G<b%� �np��tGuٰ\� .��n�t2��+h�e�w�R�e����H���v�.}����+�_O�R��Y&���vX4���9Z�p�4�O�8R<�`O��1����h��.0v�-��P
A�`���Z�C����(b�QId)7b��`���&TI�|�M�*�Tj�II�� �)4��}5�V��b�U���Ɓc�Ȝ����a1'%è��)���d��k��|@��Q�]�n�I�lD���������XU`�x���懒t���^�ߒ�n�z4�zW4�u����T¨����	����yֱsyu�� i�� ��a�kזbd��4���S�� �������g[���[���ߠI��R�F@�j�8j�r�����t�)��F���}4����(�O���㏄7���B��ql�kH-&���1�.���z�YA~z����������_�����3��P+{��$��k�\=!���� "bI�J��>�kA@�5��a��� ���}���:�����9	��ɻ��E
��k2�Tɜ04tD{F������,�~� �P�@q���[��pG�f�K܁�1�{�3e�����0؃��!JJE{����S��A۴Ģ�d��y�=���`���cuA�>�w�y%���X��U �W�,}i˗/?�_��7e��Z>��#Y�é�Lʈa`쳭J{��ao��E{�A宬�E  %E4����z������G<��b��������MU��^�6���ܟ��0%eZ�u�
�������o�ɉ��k�� �HPW���k����4�Y@��|�s���/��A�|W�ͭq�c��Q��NP�nۍ�f���1�2k�JF$�?���cfs�mLA�_(�9.թ	c���� ���s%\v��f��U1�#�d�QIi#7�cX<�k$��L[Q���r��H�-�:(�Ȇ��Z�;��Yug'���e.s�K)3`.s��\�2���e.s��z�-�֞��Ԣ�U��`�񒂁� |Xo���v�8���x��� ��|���)�#�����j��\� Xh�/��gM�V[�0��m�w9Vp׃�'���~�\�v�j�xt�#��Nm�W�!R�������K4W���t�C4 T�Ce�S���y�ay-���<ܥ�pз�4ϳ��:FZ80ޔϭ7�p�����R}��@�ǁE�8�*q�b�|��5E!A�N-Cq ��_�G����{~~��C�M�FPb�C� g�z~��*a��]�8;[��奼x�ڳ�.~��Gٛ �۷o�)�w����ii��60�s �����	T�i|q�az�WVAU��Q���AsF�0� �^կ�B��W�?�?(p�}�TKh �˳3������wuOP�\��N��Z�v������E�[�EkMPgk���lV�y�m��a�`d�:$_-����,vM�,z(?��x�*�Ơ*L�݁�� %��\�nT�ٚ��e/�<�{~����
,���xX}����Tպ"�q	Lc|\�C1�$x���|�_�$��$C�	r��֥t����W���=�B�j��ڠ/��F<ќ�[k�NSH�k���h��*?|���<yJ`��
�.4 6�~��]K�@`�\#kp�?��e�|���BZ��a X �8>h�p�C���Ѯ8)X@��9���p�_�g�{TRAR�R@��ۖq��$���6E�lԜ���l^��PQ��a���lP�nQ��D�9s�G�C���F{�$w���	(U, b ��*���x3�z�h���N$�dq]��7���FR!�(0g{0W������[��*l������"m���ZW�Z�c�In�BR9V��7*��8	�ԑ�ց_S�O����@U�W�MU�[��\�X�+	w+s�I��q��<��=����(�
s��Ìo����˳(E[�e�_����s�/����{���r���J]po�s��(���H2���s@��`)�BQ~Ƙ A�N)JFd� ރ��L�x:���p0��`1Ks�|�$��$�w�ZPS$q����?�K���8�U�5M�ﹲ�������'��S�Ñi�@d:�ׯ��q�m�I�{R��%���=�q�׀�\��h"|n����mK;�t�Ʋ�)���\�|�Ѯ����Sy���İG���6$P͎?����y O#i��}Z�ĵHw��3{QO��Z���e���b�"��~dO 6�:$�h���و���T����4��u��QJ :p_����A�~�Q>�t˩k����o]w4>�]H�9�y����̇����`"�ӧO	��]\��0ݛ�\p��z��FW���cX�-?ȗ/���S�V�ᔘ:2�p�w�4?��F:&w��n�'Q]�ih�S������F}�8( ��W�A�4�C���):a|�8I�ҵ�� �CM3{u-`�4"�!��d�Uⲻ� ���F�@���\D�!=�����rǖh�(�hs>U�3��{"nb�3��-c���5��`ݲ�Ƹ�#�Y�ڲ$	U��6��O�䧲�:��{,��146]�V~n�?���l��?l�±?r�4+ )��[c�9L�F	;��W�2���e.s��*3`.s��\�2���e.s��R�1Zw��O��v{KӅ��9`*с=+�� E~M,�ȸ3[�$r��\��6�v�G�	�=��!��l�q�4�My�D����㇒�@ZO �#,�o߾%PN[nM��Z<T�w��]�&"'�_���#���.����u�#��Mj;OU/A����m�Mن�֕����.�`��g*�7۽���r{G�*0ԏ0i����Q����	vT��
�Ҿ)�¹We����۟���}������`�}R��.�F�Tv��!�@P.wvq�S�=�̽�чʳg/x���z��C���������v��UJ7��������G�r:[�1e[�s��&a.$@1��?iq�;
���ҏa���cwj�
Ku��. ~Z��#��ui���?�G*�(��f��w��R����vۜ���:[󤆞�A�Հse�����{_��|��� ��b�c�PEJ��;��l�i�.8^�v��*Y�= )Y�(�ԺZ��B�b��:��Ħ:�j|B��Fw0��h�q�ofK@X����7�!�E����Ӕ�c����x0u-���)�Cl�-  %%>@ź�ž�#Z;��q+w����qs�D�<���:������+��)*����3�3<<>�c��Wȅ^�^\]��>�D�?}�\� l ��x�v�r�]�zg�ӣ�e���,@NhM�P�
��'`~��>r�e��oh�����	�7P��S��c��5��ǚl�/�fqܕ9%
�$J��9���Z5�X���H��Du.Q@ xo6�#�s$�)�m�Ib��u�<���Y�{ڐ�5f�����{�5' U��R_ƺӍ���	�?U��c��`I^�g�n��>[j���ŕ� �+,��JE"�F����C�V�V�n���o�������*�+Lh�����u�uc7�u��eu������YJM_sV�bM���T�����32�( z}qN�\Q�~���[ڏo֏\��:��{ls)�7�ZbPWe/j�FV�Y�Oh?��pd�F�i�˳,U�=��/���[������r��NQ��)(�ld
�h$%�( ��\zM W�;�x��<!��1i�S�k�0<R�|D|������Ĩ�zK�̛��'$!��v��6�����{�P���"W�']K��d�2P�� :biA�}Z�����T���oՂ|� ��Vn߼��b�Oɨo�S��7�!� ���d�~P�bya��#��좌����M}}�����܋�5��#�q��U��$��qI�u��Տ%�%��]K�g�l�?�$j$�-m����[�� �m�F:N��?�����gy���Ϟ=�/���d�-�xFR 1 q|8��(��0MJVg�������e/�q�?�����������c'��H"�����|���$N�g�x% ��7��RL9�)S|7��/e#�i.y�"֗l/����`��p#�u
��Zh\FM���깞i��`��'|���`��N�j^>۱#�Zl�:�W�[�oy���m���%�Hcv���x��5�7l��F�1��x48��b �
W��a�*u�� �=��xٸ���$�-�����gaq��;�@�!17:U1ɾ��!�O���Nɼ�Ev�w!����е��_͹�v�ַs��\�2���2 �2���e.s��\�2��\Y�Z�lU�U�ʔg�
���`�S�Ýi���^�Ž<y��_A1Uo+�v�k� ��t�!3�i����k0�Zֻ�ָ��M����8;��wG��[��� X�Y'�F�:���[?�S"� _��R^�x!/ ��rqqF���G(���E~w� ��_��8xƳS�d�(s��N
S|T���@��N��T��� �=�e3��v��jBS +�BE�,���� ���y���W�?o��[1���b�	-�
tyPr�3�2�byA{h��~��<-�`q8lx��=붖��{U��v�82�����:�%4��h.qP ����B���_��k0U���jc�)pH�	ԯ3�m��R�¾g�ҏ�m����-��J�rؗ��?A܀�<������Q�9�E|u��3i4%�H�ZX�"�, �nu���d� $�i�L�J�ho?T��阀]�H�2z�끶P�
p��,�� ����0����� �|�q��H��$0^A�L@�_� �\]_���u���O�X���Rw������Hu1@2Q�1Eyg���>� j�g��r
�ׯ_3�:�RB�pg#V�l�)Eb�����)T��'���p� 1���RS��?}��{��ˏ囯�����ߕ7w�O}�%8�灕1�f���&��<��g��c���`3��{�A�>������?_ܢى nu=����bl�[��o,�Z���1)00�`��,��"&P�;���͵�yY��y�g��W�}��<�ºƖ\�U�R&sm�sB�I�:�[4�bO0�U��@W��ʯ	H1C և����ƪ���������M�IwJ�x?��yP��2G��a�qp�7����M�f]���X{ ڃ��.B%+��� 8v�j32=���X��U�B���Y��s\E�:��_�W
��v��J�O`}@ly|x$g�;����������� 8��Y�T��6R��}#� 0]��ڸ/�@}u�k)�m`�hH ���w�������n�d� �%u^�����u|j��2w͵�cĴό���,+iJ�=S������/�?���r��yB��~���?�]韅�˿�V�����i��:m�T)���[��EP� ��벦����3����J�����+}7ʯ�y��H��}�m��������0�[��F*�$� �9�\��k�ASp\�8��֕���؏�М�=����C��U1.�$h�]��p���'O�g������o�q�����k;H~ �I(I�8��6bd ��7S&M�;r��M&����%����.k���~*W��|�s�l%�o�����O����6`x`����G/�����?㜂�˗�M�$��7�`�������C��/ɵ��:����H�m���:�`�`�>��S�X�p]>�
x�G�g���T���]P_�Oؓ�z-M�0�4���1���4^��s�hJ�Vt�Pw1���a�8�X��X'�0���5͍��'�n �Jt%�8���y^q�`->g*�%��L���5$Ot�Z-5fg%-@L�3q-������geOt�1�=(��8�~�;�}܃@�o��V$��.,�@�`|��4q� ��֦t.s��\��g]f�\�2���e.s��\��)_��MLUy�Ý�����"|u�?�*�������p�Q���&��Z�9UJb
rm;S͏��]J��Po4U�ZY7�w19(�|�I��I��wTw�t����/��{y��7r@>l , �Gv�$'��'�S��M�o�r8��w��A�͓'�qh��S�C�P@+�h����s��8<�B�eF���>8��z����j���[*��\�(���7n9��a���֜�!U�R�hσ|������d�<�������v0��Z��QY�4[P]:�-./n���g�`j��a���y����f����A��=�*��I��oquup@���9 �ݎ ݶ;H��!a�_{W5�kΚ����y����M7������y'�..���*�I�#��	�u��@z����Ge}Vp ���dDJ�����3 �zZ�B��� YA� �pnt�0W�>_����.�!Љ"�����Չ����� �0Er��G�� ^6�]��j_.�,t��WPuҋ�� �㢂�W$� �޼��g/��2��ե�_����=c
�����X��#g�X��+���t�:q�9A{���@��۷��ߔ�t��zd���9�	��R%<$D��9�c�
A�I��y�pGPmq��3 ������|������3��o~#�e��e�lܫVٖ�C��j�E/@ 2�a�@��oU��d';���lU��c�8bS�K��9���v�ؑHQ��Y�,�$�����<�G*bb`�G��ΐU/�1&����2Ӽ(������\�9���b� !T� ����L��0s�1N�V#��K���	 ��R9��IP�D�N�CVp;d�O�d��\����yYC�d��ٗJ(!��xA��ۊk��`:���v�)5=aN�����1 �kF��>˅��B��)RTɌР`�Hkx�G ���Aл����K��%V�j��d��\\����Jmձѱc���ܾy[�O���g��i_�yTO�!3��bN�}
�Z,����*o��ѮOnn*�N2��룂�5'�E-���¹� ����ժ��,h��=IW7a7�y��{�s/)�� \���m!@Ǣxm�pc/�=���oJ��я,/��=�_������T��KL�ajxp�IV��q\���Y��@j"��踦>�=�zQḃ�_�ˏ_�/~�E�KcY�2��������_.�ͭދ��4���g�D�i}|u0��f�`�E��Y*9_��ä���^��]y���m�9����Lё�E�#1fsa��V�EcU����	;���?W��VF�}H�qd��o�V�iw�$��^�T�;����A�@�F�J߽f�D|��]8���_ɯ~�ks~9v1��.	��؏�>�����o	�����O���������d�o \��I�����?k��AI*}����	�
��F�u�+)�S�[���r}�#���~�:g�����JgD�%�ug#�M����������AS���5!��'��JXE%�z�8o<��o�:�S�`N��Q�QG��{�o�7�ed���\��FRd5m�!�Qe��K�%�S���Qv��w粌K]OD�����R.n.��ߛkQf��8?���k~.��NYo��C�y��V���4��A�P���lMۯ���d��M�Z��_-s��\�2���2 �2���e.s��\�2��H�B�L�������a��y����*hS��rR"z	@�d |�e���롸�ϼ�ی'W5�)����E��ō�SH��M�V�._}�J�z�5T��YWդ����m6�ZO��)&��n/`�Ր[��?���R�Ky|��o/�W�j.����t�P�uf��RS����H!��ǻC��Z����۷o���-�P���M�v�k����UK��Z*����Z�Pé=)�a)���?��������hq߽��cy��3����r�c=��t��nO�>��	jU  �w�<���@������$6�~=X�|��.S�B;	���*2x;��o�\ӾX�E��NS9���Š���<�͚xV�'�^����~�6�5�wO��'��\��x[��4N)'|�$RI�:��::��~O+��|��Ƙ\o�<$��D�O��s�Cǉ�I)�$����َ �1�FU��g\�:=��e�1��蔌I��O�չ��gc�՞��1���[�f��2,�/�.��;W�����G����s v�.(�V���e��mG��������;y��-�uV��p��V�B���F�>u�Y<߳��"�X�_�^[�:!sn�~���B>|��lv�$|��)̦[�N��=���"��L�b��Q��=����G�� O5.dmcF�������ju<M�-�?0HM��.p�Ĭ�E��>lJ�ɱfh��Qe��C?�� ���GO��1 ����x��3������_��x��2�W����
k��<�b�%:�$Kg����.����ig*��1�d��}�iQ�m����7|�*8=u��rX7b��G4��
��͚f!�c_�؝�x�]S����b��˅�3 ����S�P�l�>�}^.�/{������x~ڪ�1��!�^��	3�E�Q��55DgV�R�ɝ�}�.Lp�q2��-'���k�s3縒MP���+*�ARA��tvQ�p�3�~���6B�i� ���Ğh��*=�J�Kp4�q���Q���\���Ƶ���as6)�d��������N~�7?��:��//o�gϟ� @��_sN�0	��3�b.������k�n$�g�({!�'߭K�e���7�$9(�����yµ�
��	�t�3�$�lQe5s�#�T鯞�d��t������}l��q�|������E�[p�i�?~��������h��p�<$s��`����q�ݫ�j�|^��B%(�����H��u�ܫ|��'e_����o~C� �+�C�˨�5�2_��_�x���sy��{t����$�u�styƵ�/czod0�c�;Ms "R�yu���:n}��:Z�2��8�� Q^Cl>�4 �Pc��;�`��4b�7�m}��e�#�+G�j$*�Q'��a����~ѧ ��Cf�E_n�>	��Ҏ��Li� xҚzLwP�����R�ٺG"�X�X�3Y�
�;+�r_�zѩ�{�7�I���0*ً퐐���|��ӠS�G@���*1�)��O��	ï߽%yw��u���l+Fv#�� '�h�0c��<_Eݔ��b.s��\��g\f�\�2���e.s��\��* �!��nΡ榮��Z� ��Ń2;�t,�"Jˏ BU	�
�V/�V�\.�������<�"g.�r��w�  ��IDAT�}�|�ݒm�����@�r'�������
�իo����5��G[U!�Ϝ�\�ڪu ����E�u��|���?���K?�+>?Ԙ]��3;g�3vŐ�0p/̓ �є8��Ȁv�!��흼}�F޾{C@`��A{�v��M�����l�Z'�˪�xSSE���>�L��o~*���At@;S�&
D@}�,�Z�_��U-�{�x@m�i�[*������[��A-J=v{��u2��U�8W4�Մ�ԁ"��<�U卷<�7�OP�G� .�8�_S��l�W��I��@�\�`����7���7oޘq_ǀ�~ʚ'��v�cS�U�Nб4I��r��o�R�� < .��xO6ea.�P����8�v�?U��<�E��կY����*��^���w�r_���aMǰzQ�,!�����%Mԟ
*X���o�\���&���R���x��NA���M�/_.�����=+���z�� Þ�� v ����5��K`�E�Cc���>�T+�_�3���ӱ�.��vWZ������;%4�=�?�)�>��G�bu��g���+�
C87�v���jV�-�}��IRU��h*��]Zz}G#�t���1�c**I*���<�m����'�˶�Ͻ8ƍq�yd�k%����Ÿ=�u����z���nCwJp�Q�(�U9��_:�B"�9�?��S +*���3-Ri�s_b���c���F,"وy��� pr�4G\�+�X��&�=�t����2�見���k�#�E�xZ�%�S�X��H��a���PS������HK�R��6\����)�kţ����)Q��E�ѕ�nC��O]#t��8��
'��h$�iE���Q���4:<}���i%z˱,��ZxÚ��A���� �s����Ñ����iTB��:��p�ڠ�/�C�-L@XU�י	��4���~^�������k*�A����_��@;wZ� �����/SP��`k�+_�ב��P1~ܯ��ۯd��-u;V�4�3��˭��m��5]s�Gg��}%k*%�4��B��1�;t�P����� 9����<:b��`i���R 0N���?���HDP�;S��rL�l%���Q��)i�!��. bkFpb����	�8MG�+�b޼~--5��͓��_ȓ�O��s%��������ٿ}&���T�������'����������s��zG��,��a�95%'N6,6f�4 'EKu�{T�P(c{�`����#�5��.g竺���������F�B��!�I���$�0��Q�L���/�S�;{h�����=�$zFQR@2�1I3�>([\�:�}/���@�
��I��IDA�1����ْ븥I�}ݮ����b��ry�1�.F���>b�7o����t�KlZ���\SA0��tj�������6I���s��\�2���2 �2���e.s��\�2��`9� vQG@������KU�U�@���͓Ĥv��f����ANN?���, j8��v��`��ք�� �����<�x����Q�ؑ�JwO��?�2�KUd록=_h���)���.��͢`�*��z�8A�?~�G,��_ɳ��x�	P�AU**�������)�E���' ��j�
���[( �y��j���Q2�ڲ)�] �h���9��w�U����5�������lw�G/?�����*,��R9���0��V�r8��V�G8��K@YW��Q�
�a�}�j�
�U���(�N���:Oߨ��G�]�N�Ѐ���p2 ����>ZZ����Te�-�D�ぇ� �h�;�2ߣ��[�ԗ�4���q�/��l�$��WMS���,}Z�o+��1������'�V�x�gO�TǆU��d���(�u�ya@.�Jϭ@�@�����J���I�#��?�8�_���)��xݜށg ����~��/2���ZPG�B��z�@2
�q�=�,s�0�0 L����}{K�T�t�0k�5��Hp-�3I�����F 
��&��U=_����g�#<�z}/O�>%Ȋ:`>��_/^<�������%pIͭ.ڟ�c��:\������Y��ʼ�b$�N�aڜji |�ZQ�d),�%D,��"�,��'�R
m̫�W�%��%��}���uҞ�:yh4u< |<�@�O	 ^g����2!"�9��TCd�?��J��=�I��eP3j�7s-[�����-����0�FR@7��]7s���T�C�jc:o�HF�����1i���ȶ&Y��t>D`��&�ڡ��!h*���!b��ե��H%+�G�⦺�>;��� �|�[��rU��ô8N���҆2fm;9�m�(6�䬷����W77T�⶘oe?`�
�j��X��П�y��Y�we-��hښ��b���Le�q��� ��Xo����9٦���50�{�P+�������Wy���$��O������+�����U�l��t<g�������L�,�N��v�~�������}Sb�c��e�2�߇T��'f'�X:��ڀg��8�W>ƚ�
���0A�%�_`<b��.��x%ƒ��J��TIpC��P���{�i ��� �����1�)~FWEk����[���}���ӵn��zz�{O�;��2��A�p����yv}s�k^�`�XQQ�X�� �����?|Q�7O�?���Kc����_hz��o�_��({���9ga�	�H"��N�GX6��d��� ��<�c�i�Gۃ���qu�Wĳ��,//�I��-��x��ۍ>�b�$Is�tR��89�)EzU��n{Sȃā��<4�큧s
��ݒ�8��'��%��8.�'�����ywh{:z=2��o����+�̀��\cG�������7Ѣ[q�������_\^ʲӔ[�;�2A�y���\����ۣ�ű�����t6��Mc���8�6bb:um��\�2���e�� 0���e.s��\�2��|�J�RW+�� (V�$�ť�q8��2���Sn ��TҢ`�aG��xP��$��J=8��xH� IcTp`,��'�J� ���8�M>��w��~���$���s�@jb����\�6(׬��5�@2@k4�����/���
�^��?|)g� ���6� ���=lHUu�I�S��uN<�T�x'wo���6j�n������$��U3�{�,��Z7t��YN�JX<�Ž������wH;��J�?��n�Z����^]]I�2� �{�O�v��	���sICu�pKe����\�]tlJ=��M�Y���	 ��X��6�j��-��^Uap,�a�v�UX�A�D05�:� 0� �h@�`J����Jހ�.ꭠ�*�\a������@�� ���"V�׵n��5�f-������x��	�^������@��8���XST,�Ƶ 0��. � ���^֥������č#A��
`�'��l�̑�<�44A�+8���᳁��N��{wK ��^~ /�?�my���\,���<?�Q�r~v�w���>S�쾼���W_�� $�_}H��; !;��wS3zx�ـh;4g��O�-jS�ju��T�@���� s��bJG\@��p� ��u�C�	�!��L���P�m��86P��S���q�?������A<'%վg}4�,�`./��
�j)�`5� ��8Ie�y�ͳ�l��t.*�Ô�������,�'��dM�N;q
0 �G��T�y���A>�k0SDo9B��RrT����0j��L��tM#��|��bC���U5�<�����@U��qB�hDW-��u� �9m��¶�ka=@�|c�xjJ?��1F�������`��Ti��P�KYkJ�:6[�'���+�+�F,� �hq��!Lb��18�Ϫ�N"-�u�n��I����O�ų���^nDGIF�5M� t�9��:��|񃂋:ߔ<��d�#�����gͧ����}t�J�ɧ{	W+��^�c��y���D�c��}������<��;w���'ߗ���e�>��3}���������?b<�dN� 'v���#ƀ�Y~g��V6�%~n���Q�C]��Ń$��^�JK�sW)��h�vu(PP��$;�	�?.��q�=Z��J��	�1v�{�qnY�S�{r�1��@�]�z#0�8��o5�G��,uS"��4a�SNLyn��܆�*�ߒ��asnP�׈Ra��Al���93�={�}:�  |�W?����|F�����	W_����/>��;]��δ�s=���~gn"��h���W�8O��!{X�Ftr�smQ�<d�s�qZ��5���A�
c#�<��f:)�,��tt���= �c|�J� ��SSj�|<��+Hv�iCݦ��"�D_�5��T�	���ku��6��w�SY_���rR��)+�;�d@�`�B��/.ϯ�<*��x,�[꬀=��
���ό5�|������#ݻ�y{����^����^p$�(�~�����hӽx��� �r'���e.s�˟q�	 s��\�2���e.s��w�t�.kv� ��LϛU��g{S���F*�g_�f5AU`9�|�x�b���j%�*�uُjK~ԃY��pL��1�C�49H�0����z��u<��C>)PX���������U��o���z�����I��E�����7��Gߓ������[ �yh��ǃ�M��������Ue<���Ö �8+�Yq}D�߷�u�7��r���.�2Uǃ���}z��Ο��l�����ŋlZ��H�[�֗�ΣZ�h'{4W�[�{�����~'N�h��Fv���2%A88'$� �d6�U�����?� �@���_�rq^���E�N��Z<������[��E޹��l]�ș`���*��0��k��A�x�r\%�|Oc�?���.�|��CS.&�C���<؅2�6��QG �h#��R P��č�{y�_ӽ�`nV>�Lq��Ԛ�"؜�Չh�(��9ɓ[F�i��L��o�[y��W�O?�� D�k�Ċ��s=�/�֥޸Ӌ�%��>���[o������k" ��@�p5���L$[	g���<Z�d�:�j5�#��$N�:N�U�9Ϩ@1���LQ�T�4�:@]����@,�h�s��R!��v��@T�?��w�C_��&�3h����s�Ӧ����z�m��&��I�
i�6��s�X��ͪ8������Ǧ����%Z�M@qn�g���iu���u"�0d�|^�����4�I>Sds?X,�|�&jKi� �1��Ε�i��JȦ�w��$�Lm��٧�$�J�hu3�Gp�O �}W�¡�O/ ���7h�����D�]�� �J,y��C�F� �A�	(��O�e�ۛ�Z�?ƺ�H�1��<Z�!'��0$���2:�[�qM�:f%� f���?D�k������o��.�������d�QI'��`k`���6n��a4z�w�ƴ���	�{�V�̈́�ɜ<}��;bWD�2�yoiT�rQ�b�y���[Y�.�')��AW�[��J¹���S�tK��g�9:2`���#�l��u��x�[��h�p#��Ց�����9�[�)��Q��u4M��
6F��Ƽۗ�������#v*�&՘���T�2��[O�1j����xT�t���Ř�q��fc�d�8!��>��Ck��\:�vk�c���� Z/�Vt �Ï>bʟ��'r�z�qwy��D�*���٥|y/<���K=]��r�#@��)����$}m����6E �$�|��k��l|ִӶF�@��<�`�=bEx�n��+��@��R`�2R2pϑ{�{�?�o ��A:f%#�i}��&;���'��t�N��F�12	_k\�q3����<H����*E|�dѝ\�_���E�_�� =���q����B�Q`}ǘF
���<u�W%��X?�7��W[�����3�T؃b�=�^W�:Z�����J>
Fd�?Y�5n�.:�?� �2����/�����e.s��\�2����;WF=P�y��j�%����@2��q0� ��)�kV�Y��#�#�ac���+*���:�/���HyU�	��
~�gGS��`ź;*X^�P>��u��.ҽ3��%U���O �?�����}�&���j!�	 _8R<{�\��<��k�<Л�Y2��e��"*�� p`���r�\�:���#E<9��v�ճ��8�������`��o �\_��gO�>C���r6�)VUX?�->�Gq8����x`j��U���<�S�թUw�[��

:�� �L�:XNp�7�^��-nX[�J�����vvPڙe*gm��ia4����;�����S`�S��Nڰ���@x���zhM����P��}�z�����˻�[�T`\B]
%|�'Y�-�:�x���8��A��f/w�Nw��$�l���p���ᾒ/:S�N��tn�:�'#z�'q[d��	 �GZ��z�_?�������`�M�w��~��	���~P��U7�<��^#��݃*����T��뀊��
��M�[�P��-����v��y'v���:��%1���Ǝ6#l����7���b��JNPg
�F\����ߘN@�l���y��o��j�	��֕Ȑ:���}�X^g�gD�J̷i��斺"�%���~L�*�G{$>���8V����|�l��rV�I�7�{
���?!��譯�8�gR�dL��,�^��X�N�T4b ��W��W'���7; ����ag�j��nZ��
�����̡�: (p˧�
�/��������vԬ=��T�E�+������l�~8H����J�� ���[��,V?���6�g�����JT����+�jJ�)�
6��H{S�%���� 6>�y*WF�B�����I����K��Bl,�\�`����/M�]s`�����a�ww6ДJ؜���Y�c�`["��ȶ_,����VK����BR0���١�f���	���Rǲ��=6�^G��D@�i�iK��Y��o��9�d�;����E��qO��X�t)��ԉ��k��3ٺ���qH��2�^��k@�`�����������8���-�֯�Ɲ9W�|�[��Z��:�}�<S�w�6�v����_�e߂�O������g���^���7y��-�q�ߗ:�1����N��~��9MX��^�g�N���[�bpg���o�$�����/h��Y�^E��g:��׏k��¼��ʶ�Ƭ$��k�������q#�co�W�����%Q�I]��V̭Cܵ�֢��OM����d쟞f�. �dA��H'���e���ryƽҞ�>����`ߑLU�����=�]i�wes[�i۵�GO��k��{mԑ�H�͋d��w��������]3������e.s�)3`.s��\�2���e.s�����MuU��Q��z+Ҕ�!��h��{�Z1��F�+�A�q�RU����rq8R}�0~-�-�����<x`�C8S���x�\�j'��W�f�9�v��#v�'v�Ń�09�
�MA9E��W}�#9�"HL!T��jP���g+9[�Ѳ �f��z�ܫM�^���Z[�� ����� 2u-hŉ ��)�bI�5��4@7� SP�3�Ro��գ� �F�g�X��:l5��=�r���J�`���Qp��@W������sL�I�L��魜�&U��X��%%X��Tm.؇��(��S]Y��R��jAp��(�^�5O4���GS[�Ҋ���䱪�8��1�dcj,1�_�C���6�j[&��E���[
��D�������\@qvv.7O���&xp~q���9�eC���v�b ��Úu�{��� �wY��:O�D&�a�n �)�� ���w�JLQH��hJ��SǆA��e�w p w.��}�eb� |�h?L���P �A�\���H�Z<�(��A�`�T8�t5�+�'��+1����33uL�΃�J������:ȑ�"A�����tphy�ۍ�0şś4�u�T��n?���-�����W%%�j?'W>N�����.YՅ��J����l��ƍ���Q�c�h���Hi��L�r�<�T߆0��~�>�^�*>AA����������� )�s=D�G��\�q�c�������5�.�m��O#lԘ�����}�k4�]���A͞ݓ̈gF;���q�|B���a_�-	�cm�ہ�o������Ӟ����Gz����4m���6cr�q�n#:�N�C�˞�G�*�I�a4�}V@��c�W 8F�"�#e�@���'P�|W�tM��;%��A��'{���X%)����ؑ<��vKͱ^���̶��5a�-��������͖N ]�"����l8�����wHi���4t�9�<eN$�A�x�<�:W�}n
jO��{��u��\�<"����@���y����˞�h.?WW�%�D Ƚ; ��s�e��荠X~����$�8ɦh|}r����g��;��?ל7��*�6��Ս	ϛm-��ú��k��%8-������_��S������cJR[�1g�l.��h:�K���V�ip��aOS=����8IgD>ب)y�jJ�G�9e1�R�'CF���A׏$,"�Ie%�h���0�;��1L�`-����-�hम�����ߘ�ǈZ>���~5N%�@G���8,����	 K ��P�����*s��e�V�W�KWe?Z��Օ|��nS�K#EҦ����)����zq�������qUI�Ff��8��i�O�W���^Z�t���\�2������ 0���e.s��\�2��|׊�=���4\��Ͳ\�F[�VV�]ljL����3�Y�K= ��&MP͜� %�u��=p�\(�\���Ɣ�xT����,Uw�,���V�X�p~�j�'����ˉ�\��,������_Fs�S���تt���#Tƚ�Y��R�M=�sU�*�0�٩Bp� �Tխv�[��c�Z���4���P��rs;��o$ W�F��BR�ow 81X���Z�����ި�
��%k���d��ֲ�4m������rR����(�S�r����G����&
 {[��K�V���P�T��W�~��=( �ɑ9�����o������X���"X[9`���<�:��8�TI�d��:�xĮJ�Q52�b�����ܽ��l�3Ac*��D��d(�k�,M�XA.F)��c��ݠ�;��j��?7�G�z����|�,E�����H��PKtuM�kO�(�ɖ�~��d�p��}�Ui��ݱ!�]�7gCG��Baci��Tk� ��Dļ�N8��赟����B�,4O�z�.��q
גl`J��kl� �t�90�q�^Gj����@]DlLL�c����N�3YD�>5{��bS`"�u��J�i�u�N0��~�I}�X=�������6�_�V���>3!�eS���wA׌���c;6r�$�7S"��o��6���6{=��G'Us�������eZp�8Z�z�{�)��	 ]?���jw  ,�1%rm׵`i�z�� ��')�Æ=��ٻ�ӧ������):b]��}g$'7���8�4�2�gUʗ�`� rs�G���}�QN������5�����>�q��k�"��^*�(Rcķ�06�r>uSq���1 �$�U�sG����d̳3��pA�U�?�t���ʂ���CG)�΀��CH�srB�=nt2Mv�w�u>�+���t/dc��Q��g�9��Ʌ�/��5E�
<���R�#��شP��Q���=����I$��'����H��9+�r�����}O���1������Ⱥ�A
����gr~qi���'#�;H|$��<Yے9'��u,�:cp���o$Ow_m�M�kш��k�+�m�k�:V��g��/s
~����7І ɞ�V6gF����r��3���+���)�*)����D[��?���߉)b��;#' F(qYɯ$by�aJU���IcL~�$�l9�6e�uLI�*qS�t]��c짻�B.���[ܒ<�tG�K˘���$nD@4�VNC%�����q�zG|O�kY�A�c��)c�h���e.s��\�|�L ��\�2���e.s��\�CʍH���\� ��1G	]��ܒjmnx�tQ+��3O���q=<��'��~(����8VtA���<�
�Kā�D9�`�8n�;�� <���{�
d;�L�̃h^/VU�G�g���V��Tخ���p�S���Q�� X�*+�O�Ȧ�� ���J��U  ��������b���Ae�� ������&����Zi�h`�x����h�Sp/�!i�L�_=��Sh�Zݫ�J-q�M���z{�=�A�c����)��4]���z���A,�P}p��c��}��N}��m�>֬`�J�����)���u�������)�5�n\�<��P�U�e��)���ChGk�ࠤh���q�Ƙ{;O_ �Z� 0�? wgw��O �f����~�yL0 34z��H�1fk_U�9�5Me���
u>a��z���Ƹ�����%���6���������$��XD��V�x�h�[Nf��H��n	�$3�Y�g�뎺/T���F���J����*ySo���m|�FhȞn�fBv��H;scp4Ц�uL��0RMк6����VA�9�c �܁M'rL�r�'�Y�6�*s�;s��c������a��@����5�@/��,�fݝs�w�}<;�+����8I2�k�f��
r��=����m|��=5пB1�}���	��<�����H��r��	Q��s��%��c���]�s�Rd������Y��h�x!�)�A]�;S��92�2,J��',�H?�^(���ke2�5%�ُs��T�]
������Ϫ������Y!�c��K���St]���S���`�K�o��m���c��`įQ7nX�:#�9 �ǣ���Rri�s�3�����I�һS{]�I�z�;b��tql�ie��Xc��&�ذ}Sv+�\S<�=*�>-��4I�j=!��j��:�$��Vd��.5�p|�h�� �E*���Uz[|O7࠰�w�F�L>O|
f�R�,�#����V��c��>���^Y,�>�MS�[�C�g�#�q���f]�>�q�{:
MC��h묃�
��׵��xcI�~��J���Z|-��:I���L�ߥ����iC� p��c���J�~WWW\g���$���үk9�L��)�x��T~?����'��n��C��mv%���!�b�"��%�`l%�,t
ׁ�~G��`{�kGR/b�2�s�H� h�H��*�`��ց�	1���'D<%Ǭ�5ځ�l�p?aCd_0W�8^���h�{�)_�q��S��00 �"��h�.s��\��g]f�\�2���e.s��\��*	���vEk=|7���ڭ(���9X���~�A������0/0��y>�N����!(�ù��C����VO�z5�2�rk&W� #���)q�g��s����x��?_O*��9�Ȥ@<��^��Ed�J����u��U35�h�|	�;X���>�Q;��ϳ3�DmB{�f�jD�eo�4A�p������	>%��?����Ղ
/�	��mtK�J\����1��G�T����ET`G\]���Y�����!������V�a��{4�~W]=�֨
��+�x>r4p��c��Gw���X��;�`���mk��9�=!F��Cx��	�v1����Ȫ��~�|�~ �9�d ��F��>���%i�#ٕ�Z:�Sg�V��V�:�2���07B�4�@���n���Mu �5�ꪡ�u ,$L��$8��&�d�K؝7�{gw���<Tr@S��B0�<l��ԑ���ڐ�4R�bi� J�LT��
2@A@�0���#�[�(�)7k��� }5���P>ڼ�]��T��O�l�_A��\v-���t]��Uu� �d��;'L�͆��
���M��b�9x� m#7p.��s_�]3:�h#=�����)�ؓ'�uK�1)����4 �i9�1Cl��1� z�BL_
��]K��k4�%�"�qK0�l���
�喆A��c�Vߔ�vR�h<�P��:]׮�m�Q��v]��8�>?�&�����,��������E�@Kѽʢ�Az������9�n�4�$.�:��4MI6F�S�2:�!�Fcn���6�:�8q�����.}u|(����=���j������W"wP[~���8��0��~LҒ�X_��{%�b^�m�+RU��ј�u�h�џ�m��E㱒2u�9��F��"�� DW�K�'���+�6'g#8��`hoH
p���E�:�Ʋ���� �df�H�	x��eZ�v��γlq&jj�g�\b��A�C���,,���T������7n�_���S.M�_-�M�n$Y�Y�� #�k3I��g��D�����rЈ_�к�y`��Й%�wukj}�!�o�������nnn��h�f8��`�����$��D�Re��cl��$m/t����wǲ����k˳��+Y��z8Ҳ�:g�!��(\vK�o�EG��@�Ŕ4�����-l�fK��-E�@�X�8��v��D�͕)��@S8X��:��������q�1�����#I*}n�F�fk.s��\��g_f�\�2���e.s��\��,�q�~��8��֧��Z��,�mU3Å�7gȥ���,^� jT�s��`� �Z4�ޅ��R�%wF��e��UT���s�ZVP��V��6��!{7���%�P��Y��֏*P�u?e��`U�jD~���NR��ځ��֬G�v��`Y��k}��b�+��!Q�Q��f��;H��z��I��[�&�������7:��@wS7�[o�/�[�G���Oᰘ��&Jv��>�pX'`��/W@�s�*X`�gv ��#�C�ȷ�iK���f믙z�U�!��WU���M-f��g��h��*LUd*�<y'��
����^�c#�(V*`��E��u��^���M�����	^,���ֿ١z% �����!��X)N��I� -�l�Z�k�8�zF �J�C�T�
*kǻ���i��:�1Q}cW���\�W2	� �of[�TU������y�ru~)�|���͑B�{����x�&N��@�=��0��Yⸯ�%��ު��Ҷ����c,��9�P����y�����6���L5�6spǁ�����ǭ!s������m�X�	q��'��43b�w)%�Hp�g$��������HuR���;eqЎ��b�3��橯��v�qdi!|��|��H7�Vฎ6���R�grsq;m�ϝ���^:R	1�^%�	#vu�up�˱ZY;�s���F$�E�ր늽{���@u�q,u��i����/A��5CH�ȕd�|mO�y[�{����=��3*dAtA]	~�F�[�y��
� �Q�q�5�3�B����h���T��r���3���!6��� sr�L[A�Qub��ރ����w�!�,�(u�9٥�����%<�ӝ��ܑ�Ʒ�5�J��[�Q���<>y_;�菿
F��Nkɒ�}҈ON���m�3��!F��XX؝�9��Ǌ�j�x�h,�t:��A��͎����i:#�b_9&��iu^a_���m�|}�x�f?M������A�,��k�Ƶ`��\�So�k�w(� '�����SU��=I���"��o����Z�fqu�ȴo|��C�^Li�U���!�:��&s
�*�$Q�.��ܝ�#�线���3�#�!�v��c��
�}dP2���&�?����lC_ɟ�9�)�T���c@�	�{�wb]ϑ6�
..��+�ɑ
���c�ɓR砓��wM��}�����޲�����l�E����Q'ƴM��ӣ=����"����I@C��%-T�'c�)��4
�?{z& �e.s��_P�	 s��\�2���e.s��w�t97�����MT�,��r��z`�M���Ƴ�������K�����a@UH��ԩ�[S	:���ܮ���~@����z0;��`��a����0MI�k�P 䢂^�p�ӏ�rS��jz(WA8q`$�����]�K����?4���Di��9�:0�g�J�@Н���`���2�3�fpP��&��>�H�I���|���0W}W�)p��?��j�a&UNb9�"v�^-祑\���Ӻ�s�.�-���Z�N�*?�U��%�M/Մ�宮���z�I]�(Hv�����Ym1׆�ɘ�9dm�`����E%$�E,��ɵ0W�|���x���:>\5�s8	'����L��IV��-��R7{�W�������37�;LAY�g�qБ�k*�J�p@Wܵ�@�-&)��w:&L�xd�G���rq&�Պ����)�=��A	�s�j��{��lm��m�c5��a� {��Y§h �8���Eǽ�1֎�}2�oc���Z��l<��kM$S�������%���:k��P�E���9�A-�VGs6q ��3��4�Q�7�[�۵�^�CE�5�����,n��[��B�P%�LK����jѴ����	�}c $�hN��&����t@��9�f��q
G��H��c��N��es)h�	fX?��5�~�
fs����m��ť�zS��=���b�񢱎��2>4W}���Y-��� ��s}���o�PÈ;5,z�EmGc�NGOWSB�~�㱵��ڵ�u��^�`)��v����d�}����x��$�N|��K���R��d�|������ڑ�#I�F�
�s�+I.A�c��[C��%���X�c����l�xl������a�1�����m��]{Ms��D4'�8q��������RRI~M��o��힞R�1+�|�:NI����妒���Ҕ�b?��Ms��t9$�_Ǣ��-���}OF`�um�FИ���.�~uEm䖠;�VW�����<ES�k�^��"�Bc��!'��N�P��X��w��rQ�Yte-^˚��9� �XI% ��2%J�{�9�x�;J��4:��P��u�rV�|�8?�^ ׼����+$����ϙq�x;gu��� ��j�s�[.ٟ !8��{:F�P������{���ݘQ
K�r��q�k���$��u-n#q�b�y��\�2���9�� 0���e.s��\�2��|G�0��s��欇���f���`l�����\�=}ʃ#�Q����D��^F�-����%�L����������{�wv �`�h�\A?��XAw�n;(��\����յ���9�S_���TE������HmЦ�
v���c��+��*{�N&>{��d�A�Z��a��ꏮ��C{C��o��q!��1�\��X��&'���^���.�������L��\'���k'n��W��~h�.`O^����&[O=�Wj/+Pꠎ�}wg�2WTN�&	��bw�n~�cX�r7[�\i?� �<��3�Sg��l��U���6NԶ�j
�)����d�6.�@�ܚ<W�I`�ؔ'��)�G}�zm\��n  ~���`
<�Cs���uw�l%_�����`��]��:��U<�{�l`zÙj���>UU�����|бֈ/��8��mܝ_\P1���ċ����,�^n�<��y��Y<4ps��n�L�%|)P�k_V�[系��ӺZ��7e'�45�46U�>4�����c�͚eI�31��:�.ݍް\�x�12٘^4A�?e�!2�^4FiDb� ��!����S��p�>w�����v��oUVfd���G\�|�h�^1K@���_�� t:�!�^x+� {�I�pSL����G
�Oā�,�c��JF�RTOK�B(��$1�3�;Q��]��Y�xc��t�,Zg�o�#\gw�98���]���� �G:�uC�u�%�h�v�&xJ�m�f'�cA)� S�!�Ʋ��iJp��e���,D,71"o�l߸���~���gK�>�����
�(8z*!�����߻x��Z� ��������1�_:�̡�� ���N���/)�9�d=y�./�*���	�rm��hr���uNkG�.7����W? ��0�s��բ��ķ�i��B�s��=���J��N\Ü�HQ_|�8��Vd{��)�V�s����nY`����Fm���=����{���yԽ�s�/�1��w,Pʥ�G$�?:ކj�5_�\����e��\��z�eS�F��u�b}�۳��p�Y�) ο��X��Hs>[������q�Ι���e�=B�V��pr�~1����}>{x�ׯ^�݋{�ۋ��?���+��G���������Q��\��u���ӓ;[S�Y�g��|m'fn�Sl��p��P����$<q��͢�8��:���BQ=�r��_]�6>[��;yx|����Q����FI�޷���Y�hѢE_xZ �-Z�hѢE��%��.򳟽�����h�֞�O�l�t�0Do'y��4�u诉���6WCA~�}C )�����H��	j��]"�mO�I��j��Z�[D#1B��	|>!�&��/0��Ʈ�b4�2����u����.��0d����i:Ak�
u ��p�����omFb�	�����: YzDl73BHF[����vo-r�XL#���(�y�� �i�����(;����c]z��Q6�7i��l��bi��=�]�֛����J�j�4D�G���_uC��D<�T��y�^%�.�!eN ��Ѱpt�(ԭz<��5����%J)H��j�ќ����?��;P?�x��J���J�:���9;Xփ��E jP@a�4��L*�q�$���@�X��2g�H`.ȝI2��`w��!爚����eF����a�+� �R1w�����G�����\� (�ԹiG�vOc!���*�u��,@/����P$@l���a���� �:�PyĨD3�pf�  k}���Y@$�J��T�1�����v�O$9��� ��Q�����wwHۙ�Z��9#�|{Jin:�c# [� "�	|��SL��$�4t'�!��<@xOQ- o-5�~��kt��-_+����d���'s���[u�T�W��$Rf�Tyts�b�F��=/��:����:?�Td�":��5T��"�e�΁c��ߏ��/�իW�ч��_�X^�za����g�'�������?����'��eO�Z��Pu'�p��tf����-��Ge-��f{��3j=�(y�~js��k���lp�@����i�Υh����Z�����:āj8�L<t�Fۻ=�t퍵��w��|��,'���<�?���|��j�� LÑ-�T�@�G�:��R��J��F̗��Xj�Q��Q.�A��o�_Ӻ�M:�iש?7���֠��;�����{�H�s��VϙW�y��&~7 ؜1{)ֽ��3�r�g+�}*�H�7����aԿ;?����˙�pH�Nڃ뵱�^Ζ����!qOY�e�ºk\�5}��ec�o=eH����ׯ�ַ�%��������o�o�ߩ�����.g�8VLFL�ع��S��$;��%�-��E3�4�����1������R����m����ܷ^��W��z����%�l�0�8_�6�Ue��E�-Z��� �hѢE�-Z�h�[D���^jm�i����-҇�V��������>5~��@g/o@�T�-n�ջ�Qߞ��ڌu w�N��(�D���r�pv��-9�v��ɜ�ӧ�V�ԣ�5z�X�x�8��nx��9�����M�Q���G�#ꊀ��L�v;��)�0����`)��f��{R:Yؖ�LLY}�9ͯ�g�CM����Ds"h�ąi�D�X�g= ����n�G�I��� Z^���I�ܙA¨)����3�y)�K��#����6�E+cF�'��J�K�h0Ú���pH0�79��r���\��G4��|����x��F��4�LO�]c�����������R��{	"�?TF�֏/x�0�k��%����a�;���|��3�0��9�[�8/ �Щ�ζ�����}�mD��Ȑ�6s4��s�@:&��8A �� #m�`�م�[s`<�"�:zD����ѯ�z�u�9��k/�s��*�G@��ݧ}��*.>%�l݈�Q[��8��@����%�&�r�)�o� �^bO`���&��,�9��t��hﴰu�{�k�7����߻�^����t�Gۣ�'��`� �_�N
�k�뵑����|��7#[�8�l�9N���� �({�W̻��?��v�ޡ���5Ǖ��0��02e�)�y�k�־��:ޖR���}-to�s���v���Y�&��^w��4��[b�C���Iz�l�%��/��$)i���sN�;T����~�s/I�9o�{�8b����,��_��P�E�4
�:���Y����������
�����ˍ�"��t��<�����߬˴�s\ic�V�ĉ����m��μ��1?����y�(,5�����Nm��1���s\{�N!-���7bs�#kӸ>ڹ��W���^��O��	Χé����>�H�Y�g���߅��]��Yc�Ό���y���%G�;{�o(]�%�z�}�8Y��O�������f^���0�Y*��L��k���y�E�-Z�� �hѢE�-Z�h�[C~���!طz���Ո6��0��]�F��-�� �ŕZ���:�4�Gj�l�@%��W�M��a�H�eu|��������p.��@����[�&J�홍~6,3�3�4���Aqo��*��x��Gm��4��)m%�)&�ײC�
:�G�9��L3]�x��l�OFm�)�ɒ�>�p��l,�x�1o��'� � 3��#�7sg�c��}n|(�í����"]���0�9���r�A#�F�26��Q����+7'ÿ��������q�6+��Cv�<� !f~��o'!@^	Bؼ�Z��}��q�&l��\�	"��Թ�����೉^ �Y�j������?���}�y8�4��3�t��=|����/_���y���e*3-�c�Y'�Q�S� d(�bp��n)�' �D�i��J����H@�39}�X�l��6�D��w��j�x;(��z�y���$4	�o�;:�&���R7�edQܮ�UMs�%��6�٩�H^��}�C쏡'��wX_�|����#6�$ �+��g�J�i¿ƞ�~
d~_j�S��:[\��h�z��ᠡz��l����vB���� X+c%���cͣ�NG�:���a�o6����qbX��/Գ��Z'=F ,�br�:�����}����C�)���Z�k/g�	p:�5�vv�1���*�/&�1�T����=��Pb��<�sI>g����N��x2��M�wF�����^�3��8��
; ��n����g�i���"�X!�<�k�ϊ�9l�BfY�txF�l�B��'hl��t�����c���r��SLrxM��>���خ��s��"tJ�2�F�N�u����h��c"sB)��,U�/�O:���~SG�>��q����AǠJ����Ȗ�9QP�#�;>�.�)O�Q#��༇l�5u��'��,�1��� �(;?�<]��ԡj��ғw��ַhѢE���� -Z�hѢE�-z{��z���^�����}� :�k�].��o���A�<<hܑnW#�`,ې�| ^� �5�F��)ASz�\��h�C*���B3hqp� �h�F>���:<J�U�^�9��v��ndpH�kfU���#��
��P�Vi U�xV-�l�h������6�#�-�T/�}�.��NFd3rhA`(g3�
�6?f -��g�$�b��@�Q�H� �0�����N��l��O
�p��e�*J�� Uz�GK%�mAPM����a��wYq�u�5͍u5��{�u�$��_���l��G���}����.DM� ^d2�Ӹs�e���i�#շ���\��_mc������E:S��l�6 `D���/�6�>f�\�ק�hr�(e�`�p~�$ �yi������SGzlD��j3p���|�|7�F&���1W i��5˓̔4�h�����Y���-��A��(�I�T{&�v��^��;��ru��qa��v�.K�.�|�{kA9	�����X0o��6�K�Wy:da0�V������R��1�)�W�s��@���LY&�5ϗuI�����2!�C��P���{��:%���@\瘨�Ш�f�k��uĻy�kv�HYF�讐msb0}3@���dk�!�Qr�|iv�9�5������ t8�]e}�9���j� :��@b�Ҳ{�����)�=����V��c�3Jx�ì(�C�>��u�BgA���4�}d0i.�t��z���@E:��������ȼ�
��#I���jZg��N��%
����3�sa�0���2�8���G�us�c=ֲ�����`��MZ�P���N~=�o1Gs�E�4����lM�5�$*���!�<��l��Ŏ�Q�G�ɶR�
�J�|�X��c�=,��埩��;���s���Y�A��Y:�yWS���g��D��K��!��s�2?gٝ��Ϛ������p�ս�O��B�uk�L�[�B��3z���60�?������?�]�{ț�u�f�����޵��Yي��Y ������D�W	�E�-���r X�hѢE�-Z���ޮtW��N�� �i���/E��)"g��?�j�%״���:��i�O;bݍu��YT� ���K�3����4�ۡ� S*#�Ta��a/���p�|��6�D�P'ܑ�w�Lx�Sa�e�o��3���1#b�Q?�?����@|S��\	�H�� ȿ�ੑ�R���!�N�?���V�����^�4�8��~�c�Ծ�y�a��hk��n&���[t����U���љ �=��'
	�A�|X�'��3tG��>N�c��� ݥ�P�[P�k�С=9�E|/Yι�J <=@�.���L��b� 3���$X�#���X$���w^Z��� x��Zk}ϡʐ7��J5D���u�7���n)X��:O�U�'S�y[�רn���:��)0��c8�f�~�s���#M���|�h��Og�vu��u�[���Rv�� tb��^ ���n�����/L'\�-��JP�t������N ��X7�˦v¡��������8R�o��]���O}�D�G���٣���k��&�)P���޷c0T?oԏ�g�t ޕ4�g �������¨�]LBP�m�WjB��[O�#.�q_�9�FY��f��{ꭨ:��K�n'�<it�~m1��a����5�?qSOO������?jM#�=׬������j�������z�$���q�� �K8�ؚgjh-Ϩh��r�Q��a]�M3n�Z��3���C�c޶�Z�6�i�����Q��`��ҢC�s�;S���E�u��|�򨜔���V���Y犝�Y����� �6����(�2"���߯zj���Q��}�J�m�l�7��������Q��������Ov6F�k:/�˺��{��I:=�P;BG(��د�e>K������g_W�>������+I�e�	�e�~.~��۠����!������rwR���-֫����:�/�;y��������<�O<��!�2��K׸��q��@���v]��M���� �P`8vK��b#���U�=��Q��:�N�&3��U�C�GͺFyS{*+��?���ǉ����Rb}g�����2�<��Y޼�L�|�F�|�����ÛWr~|�T���E�-Z�e�� �hѢE�-Z�h�[D�����V��S���ྎ:�����N>{s��>�H^�z%/_�he@� ��a�i��sY/���	ƙC���Z��eU�L�2�%�aIM<����?�m���2TC<���~{�q^�AR%v3>�hc�؍t�n�4��ܐ� ����s�o�[��Z�L}��k{�im`��~�����$��"���} �I�������/^�q����2�5�5���z���
�m�1�[}��ot�������3>T��N�cr �Q��bdOg`���R S8�0�6a�_�����u��~4�Z�iX�m�ˎW[� �#�V�uh;�쵄�����e��-ʫA���ѤD�� ;dOv�=�+� ׻��Fr]P��cďR\T&�z/b(a�T`��:c�k��Zɵh�=����B���!�[?B�������
U�hD�k��0��Ӏ����d���a� �S>�9"��9��r}�b�c�c�����^����~1'��S��4�f�rڶ��uنC"H�O�3�MQu�R�8��e�S�g`K��u��� �A��F�Z�KT �NZV�}����1�` c�9q���+��L-9���6Vu^��V���@��WY�2(��7�]$�F�6���n��h�#���6@^���Cg��B�����R/q��F�@%�]ci4��!���rv���k�R0���our�~S�ǜ�v�A���Ҩث]���}�B�����P j��z}ӵ�&���v����������>{�E��?�_����+��h�W�m}�	x��a��������>	�]/�o�Kw���h�o�:`��=2�;�R�1�lX�.�0f�N[���t�x�j9���g������1��T��zܯ�(�l'E�#��G�/�8�?�1 �����#ֿ9�Nw���f��0��kc�Ɵ׳�~�/�y��~w��Ƙ��ܩ���ʓ^��1���?�����z!�<�>lm�	-���2kt�-�etz�K�{O�w,��~V�ZL� ^6����ډ6��wų;yF��.3��,�rv,�O� Ncm�w��3y.V �#��T���u]��۵��V�^\ߏy��p��3JO�߻�^��	1�N5��xZ{��#������~��Y�l��3"��mC������@g�!�<㍳	K)ع������;i��]�A��â�ӹ��j֤���0�[�KX�����s+�<sj�8rr���_όO�'��O��3�������ͧ�O-Z�hї����E�-Z�hѢEo���k} �����S�j	V1��/�����y��
 owwf�F����a�ˠ� ��#���*XT_²�g��������� �/L-��4���'c'����6@7R��	����g�6�p��K�N�&�xv��'�T�-��\��=O=���~O(ܦ���Ğj�@�D�_��� ��1/̲�<P`	N�߹�7�
H����%���4���#�5�gm��R5b��a����e(zJ[�7�ȶ��(#�� x�Q���ޅ��qM�6W�KP����1�ʂTw5�F��ua�1r���
Q�<�� �����h�ӹ-�vR ����@�vú�U��(��q��"X	���	�H��%��Q#��_�HrШi��}}��Fs>�@��d�!
�5Dт��C�+#�E=N��E�x����-6�w���XOj �((G9�<����@_S����^����ڨ	XYԱG���=i+ I@ ��4 �r
��G���nC�1+;�IA¡�?��ѩ��^�L��LOl�~l�w8�`��F� ,t�q�:�li;�ࣂ��oMߩSŕ���ٟ�O �V��"��\D���4��(d��Y��w8ب�T	�d<KG,��Zva���T�$3@���"8����Н���Rd�	@R�cP�8E��r:�soga:g�C�6Ms�;��tظo3]��b��3���h] ǅ�2�}
�Aۯ���Uføv �'ܓ�n�'Ru�d������]y�7���N�f���p�u.`8�����V>��y�٧WY�������8ZJ��z�Y��k�����{�WzBrg �m׾G�!���N� ��܀�z}$g֔{���Y�7x1�ٯ\�;y���ݿR]���w���W���+s�z��^eh�k"a��}������'���ea���5����=������dt��s�;z�cQ�)�{?g�����6d�:oOO��uO�r�^7�����#`���E�Φ29 J�޼_��{��ZdH�s׷:-��� ��|qG�Z�p�b��p޳ePqβqW�1�#s���$��p^���׹��{��v8}:�].`i8�����]G��G�;�4���l�A�~h����p��;`3�~A�����vu�,�{�����tW��)��耀��N'�|��8�꠹>j^��:�ug�:{��t��^�Mȫ9Y�>?�ūW����eP��;t�B�ǡ#�qm���96�Ӝ�A3�Wd��A�ˈȎ}�9�:&
�v^��!׮!�@��TG�p.��W������<>=�g�~*���;���3�����������-�-Z���C�`ѢE�-Z�hѢ��z�J����T�60-���0�[��'��|�����F]fC�`P���� d)� f	�DD���V���=�E��G��n$3p�%�%#��|�GP�!w7�� ��`m�X�#kpf�>����69�2��Ĺ|I����=�3�
0 ��z�lAɃ^<�rb���(�AZ@� |�������ั+X�����[��n���+ F��j�sT������I�O/k����?�����q-R�Z�;��[�y`�禧��h��N��\�����y�,p�-�Ѽ�9����c���L��)�z�L��$^UG�h����<��9��`��h�)�������|����O����ˈ�c6�K޳_���n���� d�����g����x�4�h��\����\�ԧ`s��Yc��K`��,�u�����qd����輮+D�6�2�� � #�a	@#,��3\��R���^�6�͹A�e)1��(�H��
j7w裈�&0�����ڤ'<�I)S{F��wa����-�b��@D�&?�� UL����4ӌ��z����ב�3�fk`du! rO9�檥b��9U�]��:���m ��d&�_
�(���)���1А�2<4�q�U8wXs���Pk->	�z��ʳ JL�M3o���;�_��->�O�G�{�����q�r��uD�4Zf�>9gܡ���2�>�l:^�/بk����,r�
�4��33�p�a�>7"�?U9��~��Z3�\���|��{��g��?���
���9>�W��xՐ����}l��Kc�5�P�g��W{V��b~���m��@P�|���8g�~�J>��3u �5UY����r��Es�R����[������<SS���^|Z波�U�l���\�#��]Г��Zg��D��8҆Ӥ;u
"J=��#�֡m�Ω3�e��r7��t�b�8&uf��<[S�6�?����	K��q]7Fsb@�-� ��ѢcM�<�lO۽�R�#���mFa��T���ϛ���O�Ncg���W��ݘ�.��<�e�ީ�d�; ���T�Z�4f��ٽ:����נć�������g�)��"�7H�~_�$h���Di�v�)�c����Du8g"�b��V��E�-�r�r X�hѢE�-Z��-�~�V���7�S;J �N�]D����܃ȾuK����Rs�.l�0�{�v5>�Y3�Kk쀶L�m|%��M�/�0�E^�`vkqcXa��hT4�� v�� � ��a-�/��i�tX��jt�����v�0�OI@�8h��Gk4�]�+P�%ȓ����P�P�l��ӛ3�3BZ�sff���y��c5���l��*������� "҄��{� ppρI���`Oa��;H�W:l�	|Cpq9欹aQT�#.�ɂ>��n?�6>���k�1�T�$�K!���4E�&�y�E���&�P1j2�]A��p��=� ^؋t�$s��L`�/w>'��:��s��G�;yYݲ&����g�@f7�����-�v�����;@P��u��Ӿ��}���H�њI��c�� Hh�Ԇ^K�-�}��3��(x�kQ�M'*�6J��'pmx�a����ޢ}�^�ܝ
���u�2	"�'���+ln�gz���j��=�w@c46��x��/%��ŃEB[�Q
� �B��w:+�]��}�d�`���?9=ʂA�́��Y^ԉ�|A��:�t@W|?01���.���r�m�l���oڡ��_ԉ������n���_�k��a?Cj�����"�7\�X���p"��E���CVGi�KE��N������Р��l&p۱�l�d��*��@t>\x���z'�|����o3g���h8lɫw�!?��A�^Rr�ś�/nq�/X=gz���Ha:*��s�j��Nż�$6�O�~�g=�؞5��[����7:��^�}�Q��3�Ank��+�.%��B�nk�F�8�&Y������X��3���� �ۃ]��J=�y���2���s�9QX���2�3c�d�}"<[���s@�uiԝ�L����
����s����<9 ��7X��fcB��|Q�mCR��>'R'~�Zf>��"<3K�k�m����Ø����^���ƅ��5�Ltx��,��5�֒�M�o����G.�q/���>��άF��d�˘p���@�$�7��b� 2���mW'��t]�w�L]U���Y�-Z�h�����E�-Z�hѢEo�m�z-�G�=F9�b�����F^�ð4��_�� {�͌1c�Q��Nr��������S���7�v�#�͑��8����83��a+u�Es��;��Z����4̙nߥ�,@7ZxK�D��>4�	��e:R��a�ь��̞���F�[���=�%@�b���<W��RÆ�0����f�wKD�k/e�P�N)/��	ߑ�/ ��N�	h"�A����l�vC��x�s� f�p.tF�����3����au��:g��,S� -��4���5����B>m@�Ԭ���#D�>���"soM�t=�lt9RI[�e�����|�A-�| ��P�u`�rK���Q"%��;�0֦��b�Ǻ[P�;�/{�R ���e�y)&�P�ٸC:/�(!���\(���[�lw��@���	��πY����p�|G[Y>)9�wq�ĮU G ]��mŁݼV
#�K��7�0�wPJ��eը�|�Rw	��J��'Y�Z�1�~�eM@S�eQ��t�9�E[,Ǒ���|Js�
�- ~��	���ߤ�	��U'��}�|rUP�р��ιG�6��w\�4���'`��¨�)�B-�i���oV��\�����abG�ꈝ�-d��qn�g?�;��b���-�"�z�4��`��U��6O�n�yOrj׵jx��Y'V'�i�K�ӌ��!Jz4�g�g���{���Xo/O�o��1�M��>ϩ����G�I�e��:";��ǯ{�;���I�m��V��O�㝖wxO~�_���}mDf�g�Xt��=���$����AgO�ڒ8C���"������,�v]I�6� ���2���TGqS������AD� ��x ��g���֡Tt�f x�ѥ�x_V~���w��-.����C��Ͼ�Ĺ#�w��_[Zr ȧ1�8;�m�O�s��2ݓѸ_��>a��3>�C���	b��S����{:gV�X8�;�ۄx�)��U��P�g�"�sF��y0�R���e����y���ZI���
6$-Z�hї����E�-Z�hѢEo�֚���}�~�t�w�"�:"�����^' ^�b�؀ٽ��� l�mk�5<Cb��e Hf�Gd�^
S�~.��t�
�t��7 r��0~����5����((�e��?�hr�T�n.4�Ԏ4�Z�\�GEy�Fz{��"-i��4�����A@��'��T�'����nQ�f؇Ѽ�7��"�|��G�[T��	�g{����j��Y���p')��d�p���v��h��dqφ� �w)�;�����Y��ϱia�B`���������R�㻂m�\R�_�0��Z:$�,��& ��0ew6$s��Ho-�,�������/���֨٠OUS�Q��
 �87����a@�2�-;%S��M��a�J�N(X@�����`��S).G�֩cD"s�g��s��A
� q9�Hg��+
"�@���f2j�?~4����v#��C&՝�?�F�}A�	*����v%�-�h�n:�X��;m�����P:��6ѭ��&�ǵ�3���rC�
Ǖ��BH"8�,�>>�pЯ|0���]�$e@AƓ���{ʦ������Bg��������\��}ߵ�򢘜�3EE$j�^0��s��t�x���H�t��3�z�a�v��� R���*^l�"�H lD�;ܓ�vDB�(E����@4ߘ.i��}Cy>
�a�)ѳ^+�<a��Ӷi�������(���_�e�h ��!�Б.O�^�% ���#��R#�q�����^��sN^��)�g���8�7��u��/��{|<Cw�YMݠ���\U����V'��	��/֊�?�$� a۔	fK@�Y.T�!<�fIh%�k�4~p��G�%"�z�z�L�t��%�^̩c�q�nq��W����;�E����D,�U�A�:1�8/�q�<��xo<���M�ag��a��k��MImp^���q��qd�Z���AI��ym�4���ة#x.�|��{��7�4�}��ӻ�ٖR��ߕ���d�3��*�ǒ3H�1�R`>k�]����cL$����Ŋ��~��"_�hѢE_HZ �-Z�hѢE��e42�^���@��~� b�"&%�V0D;h.0�U�"�Y�:�(�
۽��h ��
����a���[��<� 
��FjN�F��
�d�zk�g5�D�4�1b��Rj��Սx���X�:!H�=m�o��-30^�o�`NA�[mes��:����a�n��3 ߁�x�XyG��.��wJ����A�T�6�v7�6D��T��RЂ����豧����M�!J���e��@��D�K�o!8F�ټJ#��)�4����fp���d�-k�V�bln V?�0؇�I�u�`�Zjş��۟-�و���y��%[͋bW�*BC��Z�@��
��E�3\[�V�ᙢ�m	��D=`��@<12���#U����l0D'<e���<$]���M�D���䬃���#fY/��c�v:��>���D�h���!TT�şv�B�S� �FK.k�,�l[-������ ��pF�Jҟڵˌ�P/�t�mg�PV 8Џcc�w>��>�#���l״5��9et"'3�o����	\�� �EX����	"|K��Ŝ|:ACMKS]W�:H9R0[��Աj������)�~0-�,���l�˾pyD͛cW���#�������7/��3�z�~�hfxu-(����?�9g���q���#�#���_�ƽ� �v �tt�h��e�����}�:�V�] ��9�r�LNK��vy�G�;�*�y�����������h���A����8U�4c��ߙ�Dw�p�1��S�G*�$GŸ�q�f=�7?�&TP�O�8���h���?�7���Ͼ_�t:�\�2>q�sN�t��U�!���I���(�,@��9e�&�](�.�x� ���3��Tl��E���3k�E�ϻ���mo��ݭWΨ��>�_�ƥ@JȾ��Y��� �ӑy�k)?G9::v_KZ�����r���\� �t:�NL�����`9��W����N.R�. ��=/+�.�z�L�}���J1�8�ᝑ\�:����o�q�cNw�h��
Y
}��/�S%��K�b�5^!����S�L�4:(ӱǏ!��-Z��O�`ѢE�-Z�hѢ���md h�.9�bv( "7Q�n=S ���	�7��ki-������C����E�� �$Yd���U�����4f22�3�*6�R{qbH7@67��(ʈ��Spz�dK���0��?!�6V8�ล����+O�=ƾL����o����N�1y��W��p*:�5�qq�
_�ܲa����8vO�N���������}��0�)�Sjל�g�d״t��G���\���n:ȯ�܈~������k��5��l����=b�<����QK�s1�� �|�ᑧ݌�[�N�[��l�U�v5_k�g~��9��~{����aD����	�in�|��-17C{���x�-���Ӊ�
tDwYdJm��m�=B��Ň���[��׉��Q���������U��.tB�T�@���Ţ�����!�i3�� 
T\G���=o���`(K��o2�uO�$���b��o����Δ�xOu�����	.��I"���D�H/o��]>�nz��r2�L��1�'Vبl�����Hu Y����O��?�>��뵍�#��|����.�hJ{8.��*��/>Rt0�ɿ�_�_�r�Ȧh�N8�]:�3<���|����4W���Y
B7��w���H}��}���7k�I���r����Y�S:��[�p��S	�Z���a[�uM4 k��!#�0�ä��l_��5�-�1d̿�p҅=�{]^���w��;�ÿ�;yzz�6��9�ó��գA��l�7�~���}�x '�2�Ĉͱ-1��6��<l?ew��TN���M���{�_�����t�_�sA�Ȅl��N))��\��05Ai?Y9��7��w{i�e��{׈9��YM�N��U'���Dq\���PƩ�\G�?#�;��gs��\�:��פ�o�zA�Xp
a����},_�}V��%$B>}n�ff���-C���Hށ�<���>xx��¾��z��l��e �C��<Vϻ\+�0����3��7���n�87q��3u��s�`�����s�-�^�p�78�8�^�8� ������nw	.���m�qvO�����&�ҢE�-���r X�hѢE�-Z��-�a�9�^�y�r�t�lmj�
P�*�Ө��M��0~#�0��iXtr˰�n�@�>F�Y{N��.Y�)��^���vK���Ft�ؚ����w�����=L~r4�ug�<��Cg�|�!��/A��5L�G��3DY�J(��&CΏ�58|HD�� cg�qgOalU�]z�.4$۴� �}^��K����Gr����@����UF,��9A�-2ʒ��"Λ ?���e ��� ����9�R ̞�sݼ� �;A	��P�}�a�ǳ)z�Q�6%���e�3:'x�>���x�����L�p>n�E��{c� 3+$�_�Y�1V����Ir��r�����d^݂���Y�M� ���4ȃC J��k��nC��T[�q̻!;>�������0���1� 0��y�C
��|����xb!��[�~Ij�m�:�v��Y�}�O�K]�	p�)s
�I�X6����>9P�r.�[�J�1��Z�c�,z�$Ǹ}7ǲ�v���l���T�H��5L0�`p�a��VG��j�_�.�!���1����!�;��T��+�.���>h ����1"�|�4�y�QM�kl��,k�pdIi�G�4_���}n[�gw��A�1RsL���ݎ��G��X��j���o��]�����ɔ��g��L�W��,vmkI��ʿ�w�������|��7XV6��"��؇
��������G���X�2�K8p���h\�9��������������7�������e88�q�hn=� ��p��� u�PB�~�u-<�`M��������L0,�C�ޙ.���#ſ�����*x@��e�&t�{���{�2���Îp�L�0�	3-x�w��q�mO	=l�n��Zsvk�_��&��[b_q=˳G��*VZ$�>�3�p}T�m�=�{��,�<7͒VҚ���Y�{��<�.�R�).��y�1�S�{zFz�7e��)��I��8�8ę����w��ɪ���A�T/��%pҮ����5��L52��K�i�s4<�3��z0���h7���CݢE�-���r X�hѢE�-Z��-���d 轵���E���0��^eDcA>KΨ~��;�k���a2\�U�q0X��'FLz����0vz4m�zO��
�0�m���F[X��%��d�S8ԍ�4�����T7��� s��Q:� kM�h5u��\fލ|4�a*�K��#����(s(���Ss���|~��V��|Ń�W�kO�Q���|E4�_�p�j�4�1�
Ze�]ܰK�í�^�>���"�f���r��iIW���� �Y��B*4�� o�EZ:�⑔��;i�oi�����
�
a���(����KL)�a�Ш8��~M��mgp�S�ߝ�����8©×��](O3XC0&;L�}��M��1a���������'�ˆ�<K5���ދ/+�Pq��Z�����r	&�H �<����p�x}�<C�G�7�`!��&��`��hI���M�Pnޏ�rH�� 3��Ϭ��í!�z%_�N$�xR�ƺJ�FLW�ac���m�_F��&O�{
�a�3��"������Ѧ[D,gu��b,i˚xcs)޻��`a���eC����8/B�۸�vV��$��C^�WB֋0�z��Q�ƒ�� �V���PF郝��A�_�"9[��[����au�^�jpT�ݴ��Z�S[����LȘ��������}�w'����� u������L~���Yvk����g
 }:�?���%gJ����"���˙�tCE6�����2D���[o���Yf�@z���������e��aC1ɔu(J�u���tJ�S&�b8��c�@ڡkG&�Б:�u:�β[��$j��0{�/vn�3HK��`5��q2C�o�(�B�X�{��t��.��}�~�6d�-x��-�}��o�B��f����g��R���HR��ez�rV��u\���hv��� ֳ�-�г�@����mQD�G ��p�'j^������࿥J4��x����p�����z�HyHqQ$�mg��{���W�E�-���r X�hѢE�-Z���n ��ZG5��/;��u�;")Y���E�;x"�ʺ~7��x�lj���`b���ү��b�b���A�b�$�&�5�v
R$�c���I�JE^�������1����A9%�`|���a0��Fo	�c�Z��J�t�'�; � ˒[DN�
PA���E�O���+ B^.�GY�i���[��У��t�O�#[ s��tcj2h:Й@��'�<O{ ^ �$��e�3Ę�1����v!R�w�/Xl�2��R�݁�������Ï(g�	6+�q?R���Nc%H�l�."�b.À����>N;���x���9���<�s\�`c�)��|�Y�
o��)=} V���ߞ��u�0o�,��WG������%~��c~��`t�E���'P$�葉i\�y~<�2�F�EC�4_�C�i,]Aྖm��n8M����!�c�<;����D�nΘw�W�)�I]��Fd�`���[K�9�K�u�ip�ib-��%t��t0=Q\w�:�/Z���Ğ2�d�e�e� �~���y�E&
׭X�u�}�s�q�w�I*�����t���y$���)�OaWg������)��D&�©��&��^���l���~7�8#˔8sj�	g".; �`3�>@H�H��.�a��	��LP��Ji?�����'�����?����):ez�����P���u��׫��!k�Aڊ�L�����Or>�\���j8c�k��&��_/�������<�'_�� X��ᨹ,�)���ٕ�@v� p& ;9$Y)"�p�����M�|�r �jF�+���\��U�FyN��Z+e*!�|E��>h���/�Uw8q�����B'%f+��BWs��#]��L&��Yc('I��p<��Z;�@G0��D����82��۞%nИ�@�mLuKƙ&�ݶ�DY��LL���X�����;�ŻG�[O:)�Ir:���B��4t^s�&�g-�2�c�7f%n��ԉ��-Z���C�`ѢE�-Z�hѢ��z?i	 ����-�)�����"ū�g��gL���vć�h
�	���`S�H��шL�n��.Gg�.u2pi��$ncP9D��xT7:v�'ܦ ��X%�D��=}j��a�lR[�^r�&�ǨFԄ�K����0?�'z����"t<�?9Ё�����	�K�3Oi/`��=�U4�`�^�o"9�-�-b�z��J7�<ӹ��g��G�et���1�g��{5jo���n0/0��4E+����p��#�Z�)��  L�T1`��
~���34�ls��u)i�=��ld-��yw p�@0;���χy��f�d�����X��*�4�ɹCk�S����pN]Gp��Fx�L��w�_DW���������,O��ls�c86��L�B�r.����t��:"�y�e�}��T�d{7�C�l]�2�:yjuf!!�@���p'�Npy�F&��Ph'��,��/̴b��	bQ*�(18֜��$��օ;FX_�cF:a�\��ni���3"�K�\�����%Tě0j���U*�5oT�)�P��������������о�Qn�����h��lsӦ}�����5�m��` �9	��Ya�K�T���f��y��3~?m �5���m(J��~����%E��@�fe2lb���*#�Y�X���ߕ��'����2V$2դuK皚ךL��;*�pd���+�+����1��0֙���@o��69$������+м$��>J5P7Щ�N��ע>��8�p��w���um�7�w:u�v��tR������i�w�5�p���>��	�Ņ�t����]�����Y��q�y*3�����2���Fg��_,/���>>}�R��5�g0g�ў�՛҃���q'�4�����:)դ��i/���m;�1�e�V8p�sdE	N
���9#��`�}yl�n� <uV�Kd���t`9���N�+V:lC	0[�-Z���F�`ѢE�-Z�hѢ���}�ԍ��2�=ҳëj�f%�F���>��� �H�~	p����M�i��� a�]7��t^�L�x�v���4�l��?���qF��pl�y�G�\���H�<ߓ�~����� $�u�i|�E��l��)A�KF %{猩̽>�|s��0.�Y�L��#SL��%^�+�Ua�&�%�;�@� ��g�$C�_+	�
�΀�d�N�~�4	�6T���iq�Rο�� U4�r0�����Tk�U�k����΋gl��NhH'ev���R���Mf��*�� �6�'�!3r�L���,�o���â�9� $|��D��`��|��Q	�{��Hl/���w0<��">睃����u�4�a��}<����%�>D}6n1F�S�23� �j!��ک��=�v��F$�l�M�m�� ��*�?}�gM��a\!��T"�3���.�!���-5��6�?�6��J�WPn�q�N�:
4�f>@g���5�'I�	芿�s@���LԸW����G����-J
 <�������d��~9�g �5���W�Zя�c�����=��%�~82uR�[�s�{��5CC�T�j�V|�L��5��Yz�k�N4�Ot�4��{����o�˗/�?��ӄ����{d��ؽ�H�y��n�,ء��K �����T��'��{_��Z#��l�ϗ���q�Y���O:|��z�{���Z��w��jf41=� :Um7խ����ӝqƏ�����iqFs9s|�3W�%fq�-���`�9����U"��4�/�\�����1���}���rӚ?<;'
=P$g��2���Q���"G��C��:"�d
G��CMI���O8K�$yMI���_�ueM��Bl_�cK���3�/Cy~�>[�_�8�t���k����{�����aݤn����:�g7ѢE�-�2�r X�hѢE�-Z��-��� #����_?g�[&���?$�A��[���.��8�&��xΌ�0x���zϹ7��j���k�-��l.E����=��ȷ"l�Δ�4�;����h}�ཐ��S�Y�U��&��<>�9h�h֏(Y�A�D�Z�2�*�$��C�X�FC��L��q���..+}�9��~��< ��}+�9�IK�%.�]i�ɳ��s<��8C��9�
�a�fb�z}7+�/!���<��D)9��k���3��҈g�����^:�L����g�,�� y����I(EV�|:�̀s����
�[�k9�d�/[���pv8������"���ͮdi����3�L��4��m��c@I���Ϻ����LV9R\a*h:"� f�:��e�W��Š��U��vW�z<_h�4��l���z�d�r���T��h)�9�	w�6��i���}��ձ@A�N'*q}�wO2��:�m[��i��Z��H\�c^]'�:�)�-9��m|=�Z��/9�ED2# x��i��_�@�/�SN�~?_�����)�:��r��`P�5�A(�$��>(��C�i@m��@���1c���%Ӵ?��C>F����dU~�=���ַ�%�_����Gz���f)��L4��\eݵ�D��"�\��{�Z�6yk"�%tT?�3A	��H��&�M�y���ݟ�rޕ�OOg�NѴ��=��Rt>�ЏG@�<{*z��K��p�*
��5f:�������aƜ�ץC���C�p^;Ε^������Iyt�N���Zz�7�XS����[��-�"5΢Y^���>�nA�Yޝa�K���R�<l/�צ� ���x"}{>��|f�u~ʤp��n��޻%-�I����՟��ߥ�?��#�N�����t8��ٲ{�<�ts)�c��hp�G�E�-Z���� �hѢE�-Z�h��C}8 lۦ�^{/��ЈH0�O|��g�����e6`E��5G�r���]����#vh�m��]c�1jP�/I�1�i>67�Ȩ0��:�ǻ�Xp��|�W6 �&@�)�N;D�K�#G��h7p�L��$i��ŉ_-9���O�=��h�����Y��&�D<$����3=�̻ L�����uc�a��C�GL��/�y�xi;j�g#��;c=�����#(EC�`l��38\f�?cVw�Y�:����~g~LP ��:>�#�@��ʩ���?g)�=�Xʭ�z��L�^]o9�UO B�ۊ�����Y�b��L��믖�,�y.�pl�X�s[b8t��1��0<Dv���>?G�������-3 ���;�v)�_\v����9<���=[��&ƣd�+9S��PkJ���^���r� �{-:]TJq��
���>Yk~�+yN��{krc������Ą`�g�ho]�S:d�����v���J����[=��	,��JAgKl?��um9�qGg�R��w�Tb�}-h
k+�m)���M�im��u��G�yz'�V�98�'��׆�t��ؓ�G'�����}U>��}��~�B}�/hG�Kp��>E>q_g+�Q��v}����:9j�>3�"�-��.1�c�LH��^ʫW����Q�K����8ϴ��{�i#�)�G��g<���6�`�G����kSdr HR��"p�{����\b(!�*ϑ�� �:�p�� ��촩�Y��2ɩ�6k���1~���RV�4�᠔�|�{6_��c�!W��v�,�����r8K��Y����_�af�=���4�s�gc�Wda�I'������]�u��c���:��7W�;��e�|f<Ӊ1-���Q��W ����ajѢE�}Qi9 ,Z�hѢE�-Z��QW�iWll����U�,���0���n`�n��'�۞��Q�֖��5� Hr�w�4H�@ �d������cH
J��Q�Z׷7��lX����?��������|�1��hM�@=7��:	 9���'��D?��j����!OS| ���s̗� c��%x�[��Iȅ=9����x�lԝ�VͨI2?���>��MrNp�^���#d'�6n�� ���!}��q�ѥ5-�)}-&���9l�8�n� R�qL����� Z|����o��w���D��N��|~�^�Q���a��y�!Ȉ�=4�����2���Z�^*)z��Q��sM׎H��X��i>J�5U3���w3:Z�K�<��t6�p����2n��-�� Dǳ��'y�w�[_�������N�k/_�O~�S��������O���i��[s�-t��N�eQ�i.��=�OF�������n�KK�?�]Y��-"Z��c_�J�G���B\0ځfr���;u�}$ҋUD�S�(�� ��Z9�i�ٟi��Q�%�YdNݭ;6ڎ1�1D�f�,��{\<�ו;��؛Y�{\ _�J*����;%��iXg�}�ѱ�]��4`�1��mp��=�Z@~}����~,?�ɏ�r���u.U۳���^���i���j!��Ē �ڬ�l��N���f|��sO��_Oww�����%�:N�PĜ�jEJǐ��
ef>?����ٷyN�ӑ�2U�{���ΦL�Kfg�:�=@ِ������k�:��_��s��{	���%�"k�[�εe�̙$뚩'���������t��7}�tn��r[���YRzI���L�H?�����O��Ì��p6��0��N�Y���������������;��@ޡ�̳���U�;�~���ם��كmѢE�})h9 ,Z�hѢE�-Z���ӓf ض�����0&�ɺ]��� 5+���K볱X�B-�1Ϡ_@u�����@9KZ� M�3�N�Ɉzd�[9��Zy��}�w�M�����S��kN+�:�x�1�1�Im�^e���O]k�1K�[g�YAZo� �}	uH�쬡#�%#��ԡ���0����ʶ�2=筃���՗n3@�i@���*1/fK9��h������#�*��N`����E�9K���5TR�
v����Y�:���`Ng�ڟ��3``��[.;��<c��=Gb��?@��L>e@s��KI#L�HB��c&��{D�*\T�ޣ�y��i7����O.�sI���[��l����s��^xgQ��T�h�<���c����8_�!��#�5� ���\k�×/������|����H����������/�_�����?��_�|V�O�!"eA��A�ď�:ڙoi�p��;�ҋ݃�:��G}�N|̊��&�,#����ܗ}���܍O-�S|nOW�>�k��L\�$�����oֶ���Cv
�6>�����	v��υ�7�i�����ݗ��=�`���[/?g@n�ټ�=_Ƒ(v̭����Y� }���$\��Y��w�{G����ˏ~���9�cP,�����]E��p^��[h�R8�e�0f#�z�2���=ʧ5�,e*Έ�§+�>x�+�t~Ҳ秳UT�3z*EB,����~Iǒ!�Ñ�& <�ev�-S��U�����g��#ӌ�3�:�����\������'xOk1w �9��������='^��	�u8A���4��M��Ltp��t��#�%f/	��k�ѳc���ɇ6��Og.�uε���u:��Z�9jT���d�'��U�4��8W/�s���.}gY�����=+��uM�o@P��r�j�����ZN&����3KߢE�-�2�r X�hѢE�-Z��-�����?���ضM���"�X\Q�ay�'#{3��Fp�'����F�ww��1�D�<��@��$Jav��;�� ���}�3���Fqt�)F���F�\��w�8<���'c���Ɔ�0�����5F�ƾp���6z�Z��ZҌ�����q��n5��̾5'*ez_n�g��a���������l =�@en���n�e~6Z> �4,����M�G !_c{�p�Ø|0e�o�K�[�W³���0�1jx�;���2q5�M�"m�-ޞ}n��	���.��O��	,��\p��@����|��%)��e�	�7O1�枣9�xn�3��>�0�qѲJt�*�����|��|� R�<*s���<O 4Î��	QWXD�2�5�T�q��I����T#��|*?��?���-}��|�kߐ�O��������w��� ˒�� 
{����>�M Tܓ#>��/���.l�x��ix� k�j�J�n $�e]�}Jzz[⿔c)�� "��1�܁d�r�ُ�Js��R��,wޖE&O��c�KO�c�w����������w�y�s@pM|��x�	��8p�`���gce:� `�;�F���(ڊ7�Y����g���ݦi�����O~�y:��`)Z/��� Տ	q��L>@Y'�������oY�:��8��z��^����n���_��~��r��m�:G�~�˱�Lپ�[r��]B��)�X9���x_.`e�{v�c���>\����IΗ�\��,NQ�ԩ��Еʆ��%�w㢞g����=;q��X�|;�3�X�Cw�/��y��1E�|n����E8�;��$���i�pX�>u=_f])z�h~o>?�����c�Y�1�������%�ԕ�L�*��A���T��͎e�T@�Mk�v,��p:uI�Ѱ�Z��PJ-�΢E�-�"�r X�hѢE�-Z���!5�mmk���|ڶʏJ�0<u�i��F7��%�!���#�0��4�-9}t�����`�KQ0S=X~c;��2E݄u�MC�5DG�|�^#J��{�©b6ʕ㳽���#���� ij�uԻd�c��v��c(���+99h/z�]��KnT�Hy�������.RZ�˳�M`��/��c���M>��X��h��?�o|�]�<?w�J�</�z$�7@u�Z�4�^i��Jж;%8/3E&��G���K�'��(�݁�0��J<�O�K%���J �VO�~��ƼV�F��o��8xᐌD~�����Љ9�5~;��?9 p��}w�6�pӅ����z�/(�<�ۦʁ7�4(��2�	�KC��~��ſ�syz|#���?�k���'���/���*��η�A�����ޞ,�84���Sь�J��͠K�#H����@�|a[�Y�u����E�! ��M�uܑ�(;o�L�t��b`�%�oDv�.��,��Y�d��֡)��-��X�{�RB�}��&Y>���lM|�>�}N�|��io�u]�9�Ƹ�����e���\�㼆Ӎ�:��<K��\��0��m��v�����������|ޯk&@�4`o�ʈn���yr$�`�����Q��#Z���`��TX|�ל%F��>�@������x�)>v����<�tB��!�x_spR���s�/�h�?�GڣJ������,9��u�9�L�9w�5��#�1���]d+;�VœW�������[/B��傶��r��� y�� ��������}���'kI�����q���<Wh�׃3 l�9Ig���s����6�}�9؏'�Tۓ>zFo�\���q�5�(7e�z�p��d���y:s�ab���kv�B�~�Y�hѢE_0Z �-Z�hѢE��etww7���Z빷�"Ƈ����>���k69�=݂\4Ԧ��Kax"��=ڈw�`�:��*5�N�i$�e�#�Z�&�DQ� �0��/jm��m6�~�e�~�[y���)�E��x�y���C�.�����6%p̂L����w�;b���{�>��0�F���)�<ɿ��SȚ���������,��~<8>}y��i����ⰇA~r2�s���R�o��n�����o��5Pw ��C�w�����%��2��Lq <)�Lfg��Ԭ=o٩��	LI��!�t&���k�W��u��>�}8՝A���a}<�u�8Hd_g����h�~%�D l ���?mc/�o~�[��'���Gy��k�N'�կ~%���/�ï~C����������,e�[ٖ���5X���.�N;�4���q>���N����P#���%-�F&߱�d�Kӽ�����Ab�R_7i��}t��-;@�W˦Q5�>��J��l8f�tx%͝��C5w`�"[�vi;Aj+��4D`���"�����0�X���J鹯�=k$�xF�A[==[o~�͇�7;�P�z�!�ZY]��)���� ��ۿ�o��?���y�غ/Zr�J{i��)a{γ���#�>2Y�kl��;
. H''�Z��>�P�����t���W������u\��[P��=�s�?�w֯z'���~��S�s����~��r�/�!�>E�#3L�qT��Nj�lq%+87�Lǖ�P����>�dߧ�_��,���20�}����%$�;��7JY���s��Ye>K^���w����S->�t�{�N}�s����N�~�d��7x��lw�~��W<���Q&x~f���X�E\o�c�@�b�][���>^;�<p/Z�hѢ/-�E�-Z�hѢE��.��i?���v���[�u���1J�����OJ4@%��\���¨@����s��}WP��娝�@��$[
�����$ۍ��y��-�z���ɮd@F6bs�u~��w&הt-���j@������� z��2��C5s�W�������x���@c���i䵱�tF��s��~c�*S��gC�E�7R��.Q�!�!;8�@��6�z��z�N:���i�b�#_
���5���J��Fe7L'�� ��l�P~�Oп��)�o�rvw��V��iDb^��[���!�=���pM��x�
�q�{H�c��3ST�.O���Ӭ�;�
\��Q���B"�s����[i��ǆ��.o�yn��}$�50����뼋��,���ݖn�n��
�,��b���vM}����˻ﾖ�������������we������|���������婝!Mޥ���
�u�0���Z����}֛�y��f��|�O>�:����'��=�ؖ *�KM^���e���u��;^j�JZ���y	ù�r1��X� �*��F/�,�9�|����Ϸ�/^bj%"񹖕�{��F��U�-t<`���Ǜ�o�� K2��{��Z��j�s�｟�v|�Ѓ�Xy^��N��yɐ�=j5�9'S�Q�n��݋�����J��O?�LFi%/E��������Z�t����#�c\Cb���]��ϳV��A>���>ryzx� �����t}��*
չ�:�[}�1��;?k�����.	��B��@�9)�%���-��/̷��`��&�ø�d����@��`���{��ɒ�>,2O�w�����pvf�)ɒI�� ],0 A�	�U0��X��	�od��ֻ),� QW��%��.�6�3=���.UuN�2"~�Y��,�͘���;uN�������Ņ#�L �+�~Z�c�n�k�'�
�<A�ϙ�%;���J�wjxx�5/��N�>������~��=��8�$ϴ�sR3/=�n�4p{��̏.�K<W�?|��d������<c�w{��#a���#(�̣�r�)�D~ֆ���SC��yz���L2����!x��;8��:�����p0K�4��H�`РA�4hР����e99[_�V�&�4��`�g�,y]h���AV����d���Q�yj`m�`�GS�� Ub�� Z �a�#r�^�E����ç�C�j�~�{Q��"s[Iۅ�y�'1ݥ� F0�R�.�s;�F�l�^1zj߃q֍���+%�~K�#Ѷ�����������A��ؒ|$E��Y�u�/��m�*��8+ ��/�/JG����B���0g�%^6/m4j������o�q�� ���~xD}/3yw{�np�րr�f�f���[|С��/���}D�j���n�'�����PS<��QS"_I��T(������y��&\p$D��8�����2Mo������D��Z��J6�S����Ť)d���7T�cl�Z��еN�ݻw��g����NtyyI���]zp�]_����)�H�T���sP�<i����@&�@��9����`U����KMW?[;�Eytٷ�5b�g%C����3QB ���`N��� +����x4�|��@��	���sZ��`Q'�����,���"������f��("GAG���Zg>>}n|R��抒ɖ�0�k{�P�T�F�?A7 �g��`7�\��g�,
��ZP:�A:���ZT����e�t�g������?�>�x�Z���4�����:)�F�.���W�i�SY� t%�e"��8���z�����q���f���N�=MU�fwh������?��a�w�%�X?�#���ƛ�{&o\����d��?�s����ٿ��-�#�X��'^T����z�a���`OA.K�CƼ`�A@��g�����ͳG�A��s�cǁ�.%�co�c��Ɖ c�#󎹴}�yU���?bF8 ڙ���8^�2G�9�k7����Z��s�WeD3�1�r��J����M�g�n^��%�_/�=�f'�6!ǖ�~]y1%��a���4�kJ�`РA�4hР��ʼ^ͧ��&�|]�B9Y�S���JF7@`�>�_+�@��T��2�=���hU��j�㎖tCukXH8�͢Ŭ3��o!Z��y5��p��C�N n�4L�x�ޥm� �����mo���o7l�I�,u÷?.�W2
ۆ(:����ӱ��1ȍ9�f�/����sG���#���E�w��2k#�`���9���c� �ϩt(p�ّ�O0z�!�<�@@tD�4)�z8�+CU]=n3�YJo ��R3;����+#����j����m����3�kށ�B X�"v0�,������l�}��*�e�~t�p-����7%�������9nc�jd"�y.�d*!*�޻(�a�6�c��(����#���N!�����2 �dq�mw���3zp��������œ�������ONh7�����{ D�撉Q�������)+�2P���^ܹ�ِ�M��) �k�~��&N��Itj�H��-�W�
|8u>�d���i��� �wk���d�������e�L�#����/�3�S��K�m�z�I#�ysq` ���C�=���J�@���ki/и�����I-,��Lg�W�7�_��П H��X=�
����G�n��D��???�o}�[��ӧ����Upw?{�W-;b�0�|%:�u1xA՛�9�gu85]$#D X� f�ٯ����f����������������)�9Ԩ|�a&l��O��}��t>�O\
�vxU��D�@??�94�L��'u���w�pY���9�*��{����Uާ��f*&��?ۜ�~�9h1>&tΣ	�W,s��3����)9h�<�џs�(zJ �?�E4���8�*���a7���ߎ9:B�x�D<�;��#+_����_{o�(�#	��ӟ1��ɧ�6�W���wC�n1�}	a�Xd�s�ҳ��^]9�2hРA�~>h8 4hРA���PJ��6N��rrr�Y��&g ��ǌ� ��Vd�E���2�7��<g\�>������3���l��h N� hG�PH�����(5�C�9�%�Z<#�����6�=���e�Q5@(�gdi; p�V�{���0��w[�h�,.+�z����\ ���5�(�E�6mJ�0�?���x�v��WGE 	c�������rj�7����}��|>��Zׅ����P�)m��m��hЈ]�"��F�)(�r�o�F��u���g�ocoi���3HL�g�"k�DV.�A���d��n4X��qC����)�S�9��B�u
�h�=j�_�ra	�*���M7x��F麾+I��I��s��
�o����z��!ݽw��D����hZ�8Yӓ����>��/_qdtt+�3��ծ/�����e��ߵ����h�*M ��� ����N�k��q�|��h��h�r阥T6��X$*]������e�9�gd=� 3 ��	f|3O���Za�
��J�� ���O�=����)� *^�`��y���y&�b� \N�ϫӴ����|��rݟ+��q�)�J��<4��!�}Н���'0Nߐ�Z`Y�&�^� �
��s��Y-{�~��.?��j���RG d�c�?��߿= ������)�۷hi�Y�e+I$��_(N8��}��CM�_� j]���s^�Q�m�%��ީ&�nb�s��(�Uv��p��Y%L��X/땘�kƂ��ў͠[Z�����N~X#���)]�:H�W���ۈ2^�ss6����~���F�5���'��2&��余���b�s%um5�/ʖ	�]���@��t[G�CG��5)m�g��~��f�a���a��#�?�A���D���H����X���M�g�v�3��_n�6���%���(�D`����4hР��A�4hРA��2ZN����i�RN5Co�)��J�����h���Թ�@SC�^�]IG�G�*�R?x�̈?h3���Bt��u+Z��-i^ hḷd�8� ��¨� Hߑ���L�Z�Ѧ���0��3�vO���3��FW�s3��r|��`�QƘ�q� ��k�<w
"b���ȣt(%������%f;1Rz�oM���\�p�]�;���B0{4c2C�Sf�A�`�?�⑁�?9��xȱ���}Q�X���B�����E�˖鉾�}]���r9���-t�uiY�c�$K�39�e��B��N���c����PE}õBezg2 ��lqF:�$��N��H>���%�D���S��\F�u������K�����@�������w���=��>;������g����t��f��6i5��@�k����Vǆ��K�Ӌ��?F z�����7�;XU`@^�=�R�4 ���;�yZ�6����G��R��w����'�������y�A `��D����ú$�ۮc��Uu�� p�����$���~��9��˸�8���.,.�̗�Rt����꽖k'{�zmu��o~�]^���?�煖�����9n�낷u�}ߨ�v�9��i��s� �Ԭ�};���1�w���p���p/���v�ey�}��~��<ɚ"2@�7�T�'28�����>֩� ꚪ�d�l�����o������V"���tA�|!��V���';mi��<���a%0�8u�:�-YVrv0%����e`�4{	�y϶̈́s�����"1���ߌ���@�[̅�%��[ͽD�g>(a��I{c��xn�(��|��q��)+�QPM
y���Sd�����.7����i{�����liR�+/X-�y	z&��(f!CF$�֗�u���_��0hРA��64 4hРA�z�謜��ҖRޕe�l:���5z��S�؎o���:�H�v�}.�-Is��ZYM����� �Jۨ�|@�hFX?K���>>׀?��x��,Z!30t'M��,�p�zu�Y���i��������bi�u:[� �7<��Ȣzw&s��Q.'�?3�i��DrZ�"����8I�j��h����VV`XQ�<�<�Ø�Z@�sK��&r�;����r����]�̵hDm��#���]_��.�k|))�X��(���y^��j�;�a:���zKD7q�jw�>C��Ǟ���G2t2ˀ+q`��w; ��eL @���=�@�u��ۂ�w��pb)���c[��50G��_ p�![D�0�D�W���q`������eV�#3]���_���?���=z���/~���}NO���>���^W��ǟЏ?����̸� �U�
��P���h �����H��z����'�M���_Թ@��e�������rW[;O��Q����ё̷u�2'����\��wq_cٓ��M�d�JY��g������bmQ 7��]��]C�,;��� �]<G�o�U���z��/��8R@a�Hx��q���:�x�9�}2, �2�IJ�h����>��=z��%}��%G�WA�䞭,G�� J��g���k�����ߢ�G#g��EGʾ���቙�������Eow]]o��[w����e�Ӱ/�r k
EF�c��A��ϳﱶF�߀�EaŽ�
%�gVe��~_�n���jEg�����jN(Z �F��ȇ	��d_�T�q�u� L{�;�  >֕�Gf���sɱ}v	�Qd{�N]�c��t���y��# y<+�~����w
2x��g|B#o[+R�Z��8�ʙJ߇�[�_���%bY4R��ʁSJy�B��Ϣ�������\���ޅs��_��x��iH����6>��ẅ��$u�����kM+��z)���A��sB�`РA�4hР��JZj�����Df��{��!�VA�������D�`>�d�[.���-z� \�%>OvQ4J��G��t5�7*��cI�ǀp=)��,G���u�ց!��@����E�Zt ��x ��{�>�LM�r��p�E��+ RA��vv���9���36~"����^�����-���5���|
��Gƶ�n)��.Q�<"��4�k^��y������3a��G`���lcn�&�iġ�}˄&B����^o}� ��H6�(oL�px��d3�M4����J�㨛 8[4#������SA�f��o{6>�{�,:��h�K]�>[�QA���tl������{�K3v�> �^L/�g�t�aPzЉ���k= ք�-��~�Y'T/�RS��3}����O?���{�>Yq[��n�$����/� u~�\��s��\�~�F�-@��~�T��G4���'cq`ܢ�9[�:��S&�O2�&u᧿mQ� <�5���<	VH���#+�Q|��[YX��E�Exc%�)�k�7���>�R�bBs�SE��S�o��9�3����)��<G�nNQ_��6s;� F������w9�3�9�|���vvvJ��}�3E���ۍhAy�:ܡ��"��cԨ܄��"�u�4���[�5D9�&yb��RPM�꺛2���Q���ݿw����綻����~~~�e �R,���e�i���i�5BXe������;Nѡ,,&�䕒���XTWm����x&+!P�k������3%x�|RL�Na���%���s���8vȉ�������N3G�uF�k3�M??��q�����)�p,�߇��	}�XS��X��9���99q9SX1'��v:Ƕ�\��ʜں������̧{�$U���bƚ��-K ���
z������8��m��k���|�ʃ7��pРA�}�h8 4hРA���Q�M-��06����>���ݐ��&���#n�_$"3���^3ޙQ*DtGj���. ���E0*v�4`%����֚�	cL:x� B9>O��C4��;ctR0zdP|hO$5�"�>�� �yucm*q�g�@�� ����ݹs�n�:��wn3H��;v���x�|���|�..��%3�W夑N ۺ�?�}J�|���4�.��`ؖ��<���7}�� �g��k.
 Y���E����U���M��mf���2hP;
p� �� ��*r�9"����0�~E��>�ysI��a���c�s�E�T4�7v��<�p���Kc��~DG�ݻ�%�(�����^^��� �__�������У!S��Sg ��V ���%MWR^d��F*���dC�w�N�H~Q�g� �^��]�M����5���^�yL�?�eDt�j��@N���&;�o�xj��zΝ�T�{��JV� -�0�L������Dp����<�H�C�n�u�a��٥��=�_:�� .VK�o��(�#�3�b��i��,���vl��o�?G4�����ݻwY6���K�9�?�󄗄i���Z{Pg���H?���M��ιd'�u֫��'��Y���}�������:,� 0s��Z���w�ϊ�W�:����Q툤FҔ�E������~�� tP ��3��)m�}�UuH����<	��XX�`��D���(]j	��s�9�}�f��/%/CD�@���#�ǟk0Ƚ��v h7�52t���.�S��L����ͦ�k'qI��ե���]�������X����vw��fTӶ����x�~��O9�#�zs>�n�2?�tu<��WL��=&���3~f8x����.��笔�4h���A�4hРA��Jک�q	a���J�D��w ��Ҙ��d2G�`lj���d[J��톦�3 �i@�#�۾��,�ݰ�/�C�]j��.6���}0b��I=�(�u8�~���+���Oѯ%�	)�aX�@�e�g���i���(����	}����l0>=Y�٭S~d=M\W��������xyJWbЕ��eMO��Pjp4K�ɣ'�d����٤/�h�R�o�26�s��sG��H����M�A5 )�s?7��AtL ��F��{[�f�u���=X>�:ܱ�ָ��g"8 ��t�X�>��66���~�z�f���L$#���GC�I��F���K ي>��&����mƮ�8�������P�P`0�]A#�����d��G�Fmf@	tl����Z��u��� ��3Rn�.����,��#�=��S]� ��YG�p?!�:�T"Q������γD��h�7�L�xt~��� �I�=[��e`b��I5�~J�����)��=��<�@eFM�.�4�k��`�照����6sJ	:����ٝ��}�r\R�}�_�� L7g|��,���|v�@��^M�	b�^���wy��}����"���l�v��/���y�G����"{c���b{C!�_��#�J`��B��F�7�i�uʑ���%KG�og�s�]__��xm��ꉳ �)K�w��Η%����	���Ϻ���i���᷎���
�\yGN�G�'��L(���噺8��*�g��<�@w����yFI/?bZ�����g��@t�[�;�����/9_��O\�c��b?S �/��?�W홭{o�� D���F,��N��Fs#�X�;)�.V�w}fg�At�mϡ�$ϔ�\u�ԝK�BM��V���fc���q�֓d�YӠA��y�� 0hРA�4h�[HZj�Pv���J�{ ���	�3���V���l6R�!P���-�q������ȍab�,Dj�;X��@Ģ`P����Gva7�)w�k�23�Q�7�Ij�C�� f�c�~�\<*�&��8�D�Jn�f@�_`~d�i)��:��b���-�$�N����z����$�8@M�]�U����k+���\Gx����*{Ėq|f!wۥ�ٍ�d���,�.���� ^X��iץgd0� �K�׏�7��^ꐍM>G�oopG�[۷�A��@dE=��F� ��5���}�Y�K��7u:=�k�↭�|���&��3�8������o���f� P`�/s�p�0p\#zS	��������=ſwUq|L�� ��ٝXl΋���ń�O�"1u�P�	�Z�A�Xà��d��V�6ʠ�n/qZ���3<_k� �Euv�}cѨQQ�X[U'���;h� l�W~_R�,)�A!�i�Z�E#o���2{D22���lp�%���A5��T�>f-� �c�G֖+H;��$��ǈ��⼱x��)!+�Zh�9�K�d_���z�\A$j�b`輠f=G���!���s|�zNu���9�>�g ����	:N�%�)�v���~��u�{�z��� ����6��K�M_�<j}o�9 9Tr�*Y�x�4���P�kÝ���J��LXSHy�)���R���;w����˫k~���v�\�n!�`.��}=,Ǩ���A�c���Q��-��N��V�A��=�������I�ʼ�RDܲ��|���]����]��G�f��DZ��0����,���@���G/¹��ԟ����@{�K<M�D�d�g,��-�?>��<��p��c��%��e�|?���C��:<�5M���ݸ0?7:=�{;�Ao�:q�K�H\6��	^��L�h�3�Ф��g��H�~�{�vQ�s���
ux�:8hРA���4 4hРA�z�����Z����PsTl�9 �n��mj��o�NꌋG�C����tC;�͖K!�>È���bO|����Z�S 4�UDz7��Q����:�-`�l{������,o��� "��OHT����L�?7V�>p� ��̉����j�8����>�''��M����{�C�������>�я��䒁��E�^���f��#^9:D�ٴʋ�b�q�!KKg���#x�*��A�K����H�ն�/�|�>Y=��������AX�B�Xz|������6����tx�]���Z�֌�I΅$��)�?B�)�5u�n����|<�U�0�@	�"�458k)���~�T@{;���C3� H�w
l �TA1�{=�������S�'ѠE��8Ӌ�:`�w�5!:5�����I�<H�}�a����V�x)%DO��%�.���r�M&�](��ȗ��C�|G����Z�D����J0d�V�۞����u�jZ�}��ܡ��K����ߗ�H$z*6���~'�c��Z <����fR�ʯ\3���G��v�����\��WQ�u�'��/�ޜ��lj���ݻ��?y�t�rPz�3C(����.2(1-YıC�\D���pu8ྦྷi�jP'vJ q&�w�.�V��2����E�����N�]�ʼ�Ò)�F�&vL����Ʊ��}�Cs�@+�=�^�TR�٦�:٦XC���K(�6ۍ���#?jf���ֶ�Ov�s=����)!��x݌)����;���5n���KU�VK� p\�n�������{Ÿ/���>S�������0�w���S~o; j��X��+P��@� {��E5Iw�4'���M2ҝO���Sc�`��8S����I�.�����A����� 0hРA�4h�[F�"�e��RJX]�ѪA�뮗̚@E^5��4c���= ��D�����R�e���r
F���qiV#@
iinh��\'��� �A��O�ѭ�l76X�����C $)0!�)��4msi�7�x�:"x ��bs��ϜNw��zU��D�����z���nݺM�ܧ�����'�ke�ҽ�5��>}F�NO���R��9�& pj;����:a�"������p^x�����\�@	<���4���SQ���dֈ�e��7���:it�h\�E�P)'t����
��u�7��G�Z '�W�B�g��ࢴ�d5?/Q8]Q�r`���DM�h���v*hu}��S!�Ac8��Џ�w�5~C���sA	}��	��`�ab��P�]��� ŵ-���xh
Җ"�,xV%��N���'D&�������!�`�༆+���>�IjF��,�v�.P&�kj�L`�ȧG�b2�����<���JV]��:��/A��W &1n��=��+�\[�q����ט�ʫo}�1��/����]z��;�w7�-��?������~�c���ҹV'.�����Y1t�,��Vu���|S1l�7���0��Y[���`at���ߧ�F����z�t8���b?kە�6�#���Ā^��>��<}��%G�/�̊�2�Od�>�tn�=D��}\ ���2�`����I�%�h��:���{��)�VٶW<s�z���f��F�]Ķ�'��3�K���4����v/Ԅ�c�:�f� :ǋ�!j{;���yUˉnݾE���j�_'E#�K��>p:<A٘rH���ޖ
ʐ��5��1Sދy�y����n�LXGXC7�qn�����Ԝu����eZ� ��� ���!�=��}��^�>8���l�����������3�� {�WT�ki�������
�}-�2t`��+�Et8'v?��D����K�Y�nM�#�n?EO�iРA��|�p 4hРA�4�-��n���uZ6�4���j�p ���)7��J�V9!�m��[z�"�`ڂ�R�@��P!ISkvt�s1��X_S��%��$f��۸F��I�"�X@-|u<��@�����}6�����>�j)�'g� �<T�r��c��6��^;|\���:�N��n�>���ܧ;�oӫW���򒞿|Il���5�_�COt�:��ݿs��NOi�ZU�Tp:�����ć˽���<b��O�m���@F�����bu�����~�'8dD��3GU�'�5ƽK7W���n� ��	x����d��!��  t`f��尤zC�b;�t#���:y��QD�����9�5�:#Hڟ�d���á4GӿЇƩE�\�"��7�]:*SS�G�1�V�����+qu�����v]a |����@P!� �t��W	Ԕ���c%y���M˭M
���MI������8� ��Mq��)�v�4�>�S�؁������w=��g������	E���B��Sߤ��W�
}���t��]Z��trzB��J�ܿE�?����=]mvR&b��6�V4K�~���n�|�G��7�.�"��>��!�" ��D.��-8�:;`.�T�6�����z����2/_�fp] ���*IƆ�g$q�b~ ��㞏 ɐq�n@h�)l�|O��{x%/E3m$�(r�S��]���l���
���U?p��
�r�L®��5c��at#�����7�����y]J ҭ1M����z��-y_�w�=zD�?�T�g�k�y^�N�?8� �G0��t}������$2��:6&�ý���	ߧ��7Q�������M���9�Ӂn>��a	��}�����Љ�|�1��3�����)��k���g��Bq��o�}M��_8��w�1A2���[$�WIe ݤ:hٚ�B���Qd9�;hРA���4 4hРA�z�(眶�]��\�Y����;ak*�H|2(I�+��)��؜���-ڊ:��G��z���X0���Kňz�X�C��0������>�\a��S7`�q�A
���� ���∰h�H�D~�/bO�7�A1��EkH%ۢ���.��0�~>?=��jM���ur��gO?'�Nh�[���V�%�B�f�?iqp&%�gp� �Mi����D̒e`H���H���t�Y��1�+jף޷�;��C�����o������H�<��nt@����!B_�Z{f�� �3f1������ ��Qgs�Y� ����M��I>"�H���ku�#8�X��yU/�@q:���ۮ�x-�{�����Rd���5k�JR��5���� �X~g*3l@�C ����4	�����ų9$�ߒ�'��v�X�q���}g� -@�flY45��4�2��~*@²�/7E��땃N)�O��1���� ���[���+^uo��d=џ�3������%Vj	�
��H���{���=����s���s���=J�<;���"#v-�Q���l$a�P�=pv���M��+ۛ�qG��A����h�K����QF�Z���ӞO�N�}���ݻwh�����W(������f�J� ��;������U��� �2)A��<c:Ie�;�$yGm����
��ܵ?k6���_m6�߷��)���H��F1�{/��m4mj3a�Z�>-�9C���
[�%c�9�����s&+ib{+O2�}(���x
r��67�l��:wm�(��cf
�M��O8������m	Nw�z���D7F=:��e�����MN p6MG���M繥ɢ���?L�n8'��Z�����ܖ�u�������n��L��p<�'��3�^�@��������4�kD�`РA�4hР��v���^粔�i��i�rl7�)���_����@M<K*X5ޚ�Q����V�d ��E0����8�s��� ��}����p�P�Uxa��{�~��� �p������r�J�̈�x>0tg 3���7�	����&7���&n4��ʒi��ߧ�^�v�����w�֝;������}�}���~�₾|��~��}����&5j#�1CF��iÑ�6�<�Qn�нus�Y��Ay'F#4q�Ȁ���e�Z�`Z0�f%�>��TlC���&Mn��VR�%p�x��7���	p��)�0ou���]��'S�sՀ��
Ŝ(a����-��z9�}Ӫ�'��$M�[H��ߒ�/�t�= f���?@:E��R�$�PU2'c
�.��$J����*��M��j��ת��]]o�*�D�(�-�z@Qp��PYֱ�,���X- C�Y?l���I���0 �Iuh�Q�Gw���\ X����^v�C��d��`���I�$,��H�������;@g���}i�7�:���'q�"��I�2dq!��}�~����]\��y������~�w�^>Ew�o�����gw�/��/�~�uמ�rXR�5�%���n�!���k�����J��������^$h��j>������{]_D(_��l�+��9�\/����~}����	���mW��tyy��?�`ܴ���D�kA'���c�Hw�ΙQ�D�����q��S�|�hORp�����/��N2�v�D�/3���s6��I�]^bt>����g�eم����|R3dwr�N�3�B^��yQ�L.O�w-<��g_�l7�J��*�UD��!\�Ɣ\>�U�t]ƍ'��fޘ*i����2�D��{s�з�����<�������A���~�;�\�yn2�P�'���Q|��a�I�����*���=��8�؞�eK�l|���yowv�Y&����=x>7��c�?�5��ӫ���2B>.���g�����`}_ٯ�\]�V��54hР� �4hРA��e��eZ��߯/���:�֚O�:5���M���p��Ka�L-^��;<J0F��w� �%��hhe��B�l@.%dP�F������Fj�=,|,�� 7r;8#��I| ��<���n�W�Q�`���-�L��G�`�Ђ�5D ��������'��J�_���)mv��ѣw��^��v�����65��R������g_�O>�����)��NNOp�vcJ��P��G�3�o7��o�����R����a-pxMڇ�ʯ9�&2Zq-�W�����!o)�4R���$�rt��~-���}\��4"7Ч ���.9�� �4]��mx&�g�� [����	�b�ix��͘����\ ��S['N@>R1�3 �(�,��"�Y�u'b`�>�R��);���'��:��T(F~2�⑶^֭Aқ�\mpߤ4�WU*"=D 8Rt��u^�-!�vt���+�^�S �ʠ_J�|oq�C���8m�$mǈ���cm�$T�
[���?�W������g�y}�Na��g��������t��S��۷�������]U�Fvu���!댌aQ�7�S�c̼Q�� �A;����@4�~ �}�.A��G��~�5wڲ��52)��y��u�^�y^�� ��ګ �� pp��́Lu�9����H.�%��p�A|}J��@��^;S�O4W99??��$ zm�:�mw��^����夲�#�<�Y6^�{���)�$S���2c���R �� �q�֒+ȂP99Y�y_d.��Ud��)��m8[�u��:ל t[�яr;��wpzН��pf+6wG����"�;�Y��v��+/��~	�g;W����U�:p�+��#�����o>8+�z;<�E'�8�����Y�7ٞ�P</��#�NR쌁�k�o�V�g��G!���6�s�#J%S���'�A��V�p 4hРA�4�-���Yͪ0
s�ON�QP�*M3Cx46j�#�'AF���4c"g5R,�TB��\P�֍��h����OAԤ|7+ ������q5�����oh�G�D�%�L�� ��E���M��nyܒ�^kl���$���w(�ȵ�~�/N
Ɍ����p�$� ~N3����/.��;�����ҭ�s�}�.]]]���%�~uAO����~�}���������kfV5�����ǒS�
g��rCx
5q4���:>��9Zr��6��P;�=8�������kq<�:p#]�$�w�����]��x�	�i��v�9Xtt�ڱ�XHށn�`_|: ��>y��������<|���ʠ����?I���� ��Al�l
6� �BdzQi84�)����Q=�5���q�&��$2G����pj�y��j��}�5yqy��t��!Z83Bn�NR��*�5��Iz1�-��m�"��A~L^]�l-��D�"r_ԧd$��a�@�Jʹ��@��=c��Z��\��]/#%��qط�� Oɜ*�i����kv��׿��oӇ�G�����vN֧����Zr������zC��/�/�q!ȗJ|�u�#b����=~'\1}�g�H�������{�E'���Q��[�+h�k�k�i�eR2h��8sd�:�g�NOi}rJ�^�f��u��2��_�H�3�{t��)Я�rɺi?�����C����w�#�W���?+��@y�=Mt}}��?W/�7R���Y0$�A��3�x��WaN��2��	�ђ�yG��Y��\~����z�Yf���My�);!2�ۿ���޳y��.�w�	��k=�d���/b����~�&��1�����u�;�|	󉳡�#�o�L�6z��������;-4��]Ы����Y�f^4�����
t<�[���O�~j�?Wc)d���v8ߩ�ZL�k����;����?�y����q�mNp�y5UY-_��A��5�� 0hРA�4h�[H+���$�ܣ1����<��Z[�TA4hM��گof =�XȊ>� �I�f�1@k0./<����ޅgHS�B}ـ��-���ѐ��-y� U1#p�f�q�c8R)c��s��W�߫��0+� �g����uԲj��֠��ۘ/��o�h;/tqyM��|F����$���nݾO�yG�^���5��g_p����/�y�����M��sV!��K.�$��z
��`8���x�LX�����D$�1��,K��Jܣ�Kw�@�[�?��c��M�@3�8|}�a V��Di�g}�D�����-�n��x_ .���i�������h�$5m?�vה��t��*HNlsa?\�O�{���N0+���aI���sr��,}�w��~}�O����NONyN/^_ҏ~���1-��p/R�%y��D�\&80�3�(t�p�!�Yd/q l�8����?`��O�x�u�Ѿ|(��z)T�h��u�������>�O�?\Vm�M�^��4v ��)oT�j)��A/��`������^�n8��������׷����?yB�P�|[�����LB*��uS>�u���M+'/���U�JK8������(� ���hu_�95�( ؗ~*�Y�N�������[�̯�l��Ƴ}�mI������rҧ�����OqN�낍*�rP�3pā�,|��i���{G�!3�{v&�v�����5��5�v�����2�)/YM���.�v�g����p�y����:��y uS� ���{���3�/.$���$���-�&%�Q�;#&�:�ߙ�l�4�8�g�xL���PN&��\�Gb��;+�ǌ'��k-E����c s�h� ��h��v�6^�g#���'<	]t�le{���~�kǎDΫ�]��4���?Oc���	�q
��,����Q��ر�;�Qx�9n٢��"�A	���7r������4hРA��v4 4hРA�z�����,eW���%X�̾�܈���x�ߚ�0DΡ�m��mz\��I��!0`��j�)5Z	 D�n9q���R:��Q[�qPl���5g�Ȗ�!y�XeLn���k-�`+>�}����=".��C�d�(��,M�����6�9��3&���'`XE�հ�F�:[��L���...�/�����}�.��N�z��'Ϟӓ��8�x���f���x�2ʬpI��q������M�c�ؐ�yn
�a�%�>�h��9`���_1���an!����`���.�t`�8��)�_J7/���2�����9��,A�I�b d�8a����o�I�0ЂU��T[��)�F��o� �4�z7Z{�-tr�L׊�6�Ȭ��+տ�Z ;�3IZW��d=��i��޽{tzz͕g���~�|}Ie*V���lr@>�)��v@5� �2P�BkM�o����zW��*8قa-x�ٳEu�DpG�,���&}����'Ţ�}.���@JQ��5���8�v����S(� }���x���[>jf��1�İߟ���l�{]���+z��w�.gS��������'��~������<d�YR�3 ��*�?�K�?)0&�|v�N�A��H�uȒ��z�Tv��;y�� zC�?���"�%æ�s=�){��?��f��W�������+��~]����Ĕ8��>e��O&>��_@��6A"��H��,?V~"9�Y��/'d�DS&&Guh���Ν۴��H�oͼ��-�2?O;汜.��$3��:AT����FS(�Da|���2��Z�_e,A�0��t�����'�\���[Ӌ�/u�������i��|φ^p�(�|k+���B�N:��f���-��^Z�q�|)s�U>©7��_C��.:���}��*�w����ٖ~{OЕ�R9�ܟ��&v��X+�ksN9�Aϛ&Cw^AW�	<Z���]V�)~�>�ct���]QN�j'�v�s����;���hРA����p 4hРA�4�-�jo�����>6P�/Y�?
�	1
f�N���ـdP}�z�I�Қ̚I ��C`��Ide⪰h�ߓ8�۵(�,���@����nÖ�5�)�yH9/"H���� �g�k��"���ޕ�'�~�M�!����QQv�;H���l��= J�@I>.`��jVoR��K����D�	��1W0a�N 5u5�rI� I�+�@M=l�N�@ �?5�7Ѡz��c(nL}#3����<P�1Y:��7�^� $����E������u�!^�6�s�o�	#��Р�ߣ�8~O>����e�.�Գ�F��y�����
na�5�*�1�P/��5�JΧpSë�5{,��>��`�KjT/�� c=�ܠ�Jxi1H�"����&����l��E,���ߓ'�SӘd� �Sҙ�?u=�Zߵ �8_��������g4��X���̇;Bqp2+�:/ ��Y�P���}�k�u }>x��R��|�q��,6�/���<3�v��S��f(3T߱�2��@=-L��"Ҏ�R���O3�����Q�������K���5��oZqv���~�����[���^o���%�η�M_<{F�%�\�
c�.�^[=���u���և֎ֻ�6<�cA��#�
2�{\�(��a�����3�L_�H��I)�a�!��4͖r�_��W�_��I��iN�����/K7��T#��;9��6>�χ�¸������X�� ���93Dc�7�-�_u�n��D��^H0yq�����K��>c�I��:	D�ړ8")-U�V��;���\=�)���=H����~/�Ҹw���.5l�J�G�G�Ɩ:U�d"�{�M���ȯ��ޖS�s.0К�R�!�M��#���X�����W�`�`��4�l>>tc_㭮���=f9�?�w�\�����ވ�տ3�]�:��3��Ȉ�������q�֮I2�k��t��Yby�4h���?hРA�4h�[F˲���y��<M����0��ui-�Ț`2R@�ɒ}�A�\�߬N�hT%���U@�A�e�]�^4�ȥ�54�U��jd�V+:==%d/��8�`K	�	fp\��ˎ��*U z�N�VKpF��s�i�G��sZ%��mSI[Ok5���i���{��jUTCp�����-��V0�oH����D���%�� Oth�DZl �E����n@Bv�<9EB���Q��v�?��A�bk� ��6	`#����L�����Y��#��m8 #��f4���
k���w��h�ȍ�Q6���c|_�}p�Ȩ,wQ ����rnQ�1-u��,��U��D�h�(��6d�x�?  ��y�f�*5���$1Ҵᩫ+gb�:-�R�H��������Hj�p��;W�6�	��������XjV�ιJf�S�'�*딴�t/�7�(w�]@	HǴ�c^���⚦���k5�����!����t������Iy�l����8�Q�2��o8�.�D��4�~���Yw�I���CI����= �Wyj�M��@�Q]���u�X���}},�#D�g������!Rnj��|��&9��e��D�����n艁ӓ�d�W����~^�����@Ϟ>���5�߾EϞ=���SN?^��<
r�Zju0A���Tg�U�x>lmj$��wG$w��B0����U)(��
�ӈ?�דf�PF�..: ����k� ~%��ӓ���ͥ��N8�T� �=sq�m1�3�Y8�x&����(���!�[#��H�ޟ�>|����y\]]��w��g/����I��Q�4�@�}Q��D�D!��g�0��� �K�5��8��Zc�\�u�ž�W�γ~C��K3�g+`al��]�1�������C�`�3��&�z]p���KdF8|�07|������9�uD��D�)�?��^o��8�.8v��g}N���#��������3F۵���s�|���Y$2�s^��6s����be" �҉�(�Nm�xt���	/�ώ��q�,��Τ�����+��:�]��<��gРA�}�i8 4hРA���Ѳ���(�9��� ��ڈ��1�M��_��
��H���$��L���͆GY��� �4�$�0�)pUR5=��G��o�ݿM�}�﫠�I�[�oK2L������s}�y����P#�* R��o����?�	]]]ѝ{���o|L��ܖs�6�w��sb��	iI`6�n�c�ngz��%=y�>��O�;���:g��������lu4��9p�(-�Ψ��_(�I�[�CA k
� ]����@դNnz����m�A�I���`l5�P�����$* A�>�����j��l�DR�eHq���-�	�A3��xN�3t�� 
��Q �uC9r��,��b�lc�h�|S�E�����ţG{Z0g�#�6�e{� H��'�OZCy;�%6o�PN݄�$ٝ �̕�+�
Ԧi��VtzvB��NO�HQ=v(b�� �d2��݈�g����V+�]";�y+y��}�^1��z6IZr����&qX��8*j5��[��m��gM��Gѽ��8K���sz������}��7���<���_ѓ�Oy�5�<TBD�D�WZA��v��?֫5������^����^��T�ę���U�߿w�����]�ӕ�U�__]��dMϞ=������c���d>rv���8P���옧��U���U�v��q��}��\4+�N�/��\�d����������e�<��󶓽.��M/ P��Y��
,�jT�uX�DR!!�D鋞����!r��,  .�&j�˞Oϟ����gO__�O�׻��1* ,�D��$�!W\�I��L��}Y�'��t�3�}�յ�`��l��"���;���q�._�m��/���@  ��IDAT8�4_`��"8��@$��D��t�,�ח*n��HRg/���y�W��+�i;�:�9~�LH}�utt��<�� L_�������{t�_U]^^���y�:��ߟD����"s+<���1:��qfП*��>�PJp,@�� �J3��YrK{~�;��!�d�/_�Yg�!KS�LB�ȳ���(���w-��,C��v-aE� �7���{o��o��#�8A�/G�����������/n�I�M]?�1��2�0Бuw�\r���y�����l��e���Z�L����<+��]��#l��@���D�e������ǩ�\m�	�5hРA��V4 4hРA�z˨f X��������<%�0,nm$I�
�8+�' g�3��8�'z������<|D��)m6�t���/���H�}����&C�-n�-�}3q�o�*_�W�+�������Ig�~���M�+��.��E�j@	�w��l��'O���|����_��t�o)��]g����ٰ3y�څ�������w�[��[���K�����fѺ���>��������C "k�5�Z�������kM���r�ؚ��о�$�
�9�
���]�����g-�Ф5��^+��SZ`�q�5n7c�_��b�� �6v�+� 0i��O
��0#[y�%�{)0�{�a����
y����G���m�h9�"�F��`Q蓽�e�Z�,�>����e�Ӆ�ۢ�yрC�<Q>��n���sw�Eg�M�=���QĹG@\�T��Bgg����������θ��=4�3��7�i�Z�"K''k���Su�j��3�$mG ��_uh�'%O��w�V�q�+�^�|E/^�`�v~~F������t��=|���'+�8�̥VE�R)�Ff�c�[|M���s�?m������mi�m�c�����0��D�#j�S[	
8������A��,��L
�3|D�j�1���k��6�\	�-N��]%�w�oiA!D]C�$ ���zu��)��޲�߫͆����K�W��_�w��]�x��j�re�E�V��"=u��T>f��Wp�׈��,
���Y�9�8�l1�?tU1݌9�l��X�E �?n�X��5 yُjQ��s�G�%ߋ���JQ��E5KP=�����ޙl~��E�b}ۨ����v�G��m� @1�GtP	V�: ��I��B�U�QuA�M��R8@uv�N-��B��h��ub��sp����C 7_��$��ԡ �7c?Q����A��g7���r�x��F�l�m�y*��H��Ĺʹ��aܭ�;�6{q��~��l�S��JSf��{B���㑧K	�$���:6�2/�r�m�ýsܷ��~<�����2.3�S��'3���38��l����r{L}��LS��P���m&w�Yq ���l2�LH�	M���<Sy�9L!��zR��h��H>n���rjn_X}Dp��=@��t�؛`РA�}�h8 4hРA�����۷K��.缫��
�V���bP;����V��;����@N6�f�`�Qs�/�%�s�ɯ��$qj�S�����?�/>����8��õ���W�=5������ՊV�^u�h��P�m�K��T)ф��84�b|e#��h�������VT*(��R b�V�	6J'�O�X'�������꿦���c��{N֬�Z�j�����#�Y�I�ڂ�����" �UjL�G(����L��1�-�K2�J3�V��y1��=WB,Y���������YD��	g\#�����Q ��g�S�@���~�fն/7;>��$�� ����[���(Dq��u�V�>���H�5�ؐt D-6Ѡ�9� �8��q!�5����̲Î3�AF�W
R�;�X2��b����N,|�Dx���N*aͧ	��>Ϻ%�-��jd�_���)}�s$=��GT7։��#���ɀ�
y����5�mXL�P�i�\��k��mE�]�s^��q������o�;vTx��Gt��}zu�>��Cz�λ\�����'��WV��]���2�ht �2�l31�YR� �;�;��:+V�AH���@�@�t'��=�	��J��\L�]0Z �B�y�����sD",��,�S=�*���,� �R>�f��𚝷[����G��'?���[�I-?#94�[׆����"���&��
;��l�����^����
�լ?��4=~�}O8C@= "W�=��C���n���U�5�<�'�'/1P�03Q���� ����®��lX�V��^�|Od���m��:���ѱ�GT���H2%k[F06-�U�E����h�9pM��"sXu�;����_�����fGp�w�X��3Ɛt�A�?;�d�A�n:����4��;��z�<�l*?��A�Z��3F����:��<I��]7yI8�����œ�+s角Ųg��k�<ю���4��� k2�C�˷�N%#y�|mP��t����-�2SO�,�N(ro�D#���7����z���ܨ{�ꤓVbc��5��s�A���8�QӇ؞�ע�= �-�{r͞��`k6œt�5��*��/�CxM�K�|����Ɵą�O��v�*p6U)�ʈL^�N�t�Ϊ�J�%��QJ��A����� 0hРA�4h�[FsERV���YOKJ��(�� v���tpQNb䗟��jd��銍л��7^ϝ��E��V�2	� Q|I�_&5fi|y���
XU��#�9�r�8K�_�紐���q���~��?�o��e�o�ݿ�ѸY�f?g� Ӡ�60��S0��}����nw�����������ǟ���)�!O"���x�Z�iQ띁�0� ��8��n�鉑]��bLQ�j�,��7�m�t'KF+�S��+�o�(LX�po�R�#��9�x���Q�Ev���\��G#���s�d��ҵa���_M��h� �N>;�[!D��\[_KL���;��q�g�r�aR@'��G�� ݔ��ls�@�Sx�d��Qǯk�"d���)p���DVW����¥F4�S���8)��'���_o�E��#�9dc�-��XǹSL�H������cvR�+���O�_�s��$�����֪���|��/��� r�(a��$�� ���{��}��c.[�ɧ�ң���r �<��-1�?5@D�׆g�t�\u����1�:�|_ #
|�
ވ#F�W�"4_��:�������RVx
� Б�e��_ѿY�d��A2�2�d�f��R(�hAj#yCWMO�X}%; �NRR�~^'��_������]ov\��W�+ä6}�R�ᢖ�A���R3R���\Χ�$�B�]�����v[��EK��2��L�-� )�Z�^o
0�SM�5��Ct��@�!��:�d�?�	���H)��3P8%>_pd�nG�6����\ܡ���F^ܡ$'8$�yJ����x^�34a?�M9��7$uJI��;�g�hpy)�:D�$S�E��pQ�S,5i�⠀��F�M���'�ф~�\b�"����m{��S�\�O{�2��/i�߰C���䳜C��C}Ȓň�wƓd ?���x�S��� ���(�cw��n�wǏF�g����Si0��k����V˻���,�/z�p���4�4��:x?^�� �yM,��������$���8�?����Mݎ]+���,�����Pv�HQ�z��l�V�j��Bq6�S��u�~l�����@4hР�����A�4hРAoU�[�����ds�Z�S��u*y���P0�RkO2J�������Nj��5�����V�'s��Y���p�������w^)�%��ͼ�����;��_����O?���?&���g �Y��l�̜*���z��ǟ?���	�����W��ԁѯ��~��	}��O�ӟ~B�_���w���}D|�=|��}&dj��'k�;ݡ���ߠ�����LPǛ�d)H���[_�����AwD�b�Z �P�������H6�%�GL���  �5ƶ: m�08.�~�MJ{;}�O�"�Zq���o��Lv(�dF�ҦĕȪ�(ݴ}̸�}��Ҍ{JY��
R�nT �"8 )9x@ͼʑ���,x�Ð9��:��>ǧږ�E<�gϥh�@�C�%C@�Nd�![�=l��h�����Y��V�$�U����F�J���]jV���kɜ��*ب_8c	f'��d���]�\O~7���>��O~�>��7YWl�>��A6R+~��܇Z�� �Uϵ�gqL*p&؄4����2T��ͩ��Kq(����Az��:�EjxW]����^�z�@ot��{���*�ߥ�����(p�Q����[���z�����:���������ȒR��Z��3;o��<==�[����٭�}���?�[�nѴ�VKTǊ
X^^���>�l��]�߽��>��Hd�^-���ye:S�tE�g��R����^*���6׫~~��ŤN%"��9��j���C�	o��C��:ou.�C���ꕚ�&���ر������[�������׈�u-�Pϒ�[�6z�_��n���tM����5�'���"��8Vǲڿ��3�w��9??�w�?�����H�ݣ�_|A�r���~�����~��nfz��%m���}�J��o����iuB�28�"p���p�)�U�%�@0��� ����b��M_��ԇ~@~����T���}��9!^V�}ݲ��Lh߀��~
���~��]���A�w�"����;Б��XI"�=z�����⚝��{�"g�%�� M�N�f�Gp\`G��|  �=K7w�	�
?�� �E֒�̉�"���
�IR֌$� ����a�r���n6�=�Y*t���{gU�u�g� (�f��t'���bM� \峘g H\%���y��l? ����9NHkA�����u��̀�8hؾ7��q*��i���Φ�����-+b��Ov��dI���IJ�ɻ&�:q��R�B�B;x�|/��p�����*�ᨢ�f ?���D��~d�^�r>�9��25��੼ �*m;E4hР� �4hРA��ET���<y����7�y��_X�H�`j#�5��̈�M��� �$4&5�%�����f�:�Z��HJ{���H�I�h�O��ͿW������}�;�a��v�a�Zy���@Cm`�҉-f��i�+(WiQ�ի����G/_��w�;Nq͆Լ�ޡ����������f3�*I��d��_�5�?��?g����$3�۸�=?��"杚������������ $FuD;:��эѸ�3=;Je���jg5 !a~�W����<��5jGI�0P��{�d���1ҿ8�c�����-����;�4�M�)�*@� ��N�6�1��p=���ҁ�;�7���I@�:��i$�u`�k�>�%^�nH����&�Kw��z��C��_�z�އ�uz���ι�
J>��}��O����'?�)�����n���g����	hf�j��j�}���_N�^*0}M����I�?!Uof����3�þ��@�f��$�[��S`��Û�;���D1 :)�ɠ_�R������_ٸ�Г'_ҿ�7O��UWt �EYD�.p☋Ej[�� ��H�
_�_���Ġ�8b1�7[�d�@� ��N�V`0�	�e�Ǡ�s(� �&�!�:��]�����ۏx~_˔�~��_�n�c�4�X^�Oai`�վ�:�&`��,���SKf��ӳ3���}���ݮ����^F�L��#84Ԉ�S^C��}��t{�n���^_m9u��gW������.D'�a��w��yM�$����5=���<}&�uU7��sPK�V� x�=������˳����C�r,{#��3DG�yi��&<�7(֪�fA���� ;�_�����&r���c.��N��Q��}���w�}��9U�\^^�Z��5d��D�-Z�z���H���L� �p����1��/���P��t]f��la�R��%A�a����P��|LR6����8w�,{�.(�����?��ߣ�Ks|u�<���,2G�B_�曾�����e2�y �S:�)M[~n �YG��.Y3GA[��-�n*>w�E���"�̀������龴X�
���@�,*�{�r@˵p��E^4/[[�,�Måѫ����s)����O?����bРA����p 4hРA�4�-�����d�W��j���e)V�ь�b�ђ�DѸhv�`�{���J-6Q��H�w�y�`��H.�û��,��m1�!��W�@q.>����/��E�	���'ۤ}��Oد�VC�٣j_�z�ƾ��V"Cw5j3�z]A�����}���aPW����S��􌮯.j%d"7ɍ�F
����� I�<��;�$��(����ڢ�iɞŻ�}�_��g��3e���_��$
��<��uN&
��Ox^��.��6% ��;J6��� �D�F��L`$�mrXI����`P)H�!cR/��B g�l4�W�h����_���@&�qe�;D�-e�( ��CG �4�S��d2pv�y��&������+��i�5GLg�k������>��Gtrz�#�k�7���ղ���p$�?�G���z��9]m��:(ֳD���T���۽&�l5m6�abǣ����}k�6���D%T��AMw�K����!;{^�� �{��U�p�JV�;����M�̀��2,�������RuZ��p�����^P��/{o�[r���̽����N5�TRI�$����Hbr��mh9���`��G�����#�~��n��a�Ơ��n��JBU%��oM��;��v�s͹�-�{�vVܺ���޹3W�̻�o}��o��<1r? ��WQ� $1p��7�!; X�]]w��:���e��ʌC-���b?�Kԟe�Xg�D���Lv�D�ÿo��r�,<�(+G��Ҝ\Ԩ����N�C}�i�|-"�e_��� ��8��js��%����W��9��,��+!��v?T ��؄;�>����3���=��݇��_��>��B[��8.k�+�bW�K�r�T�@E����2�2�Qt���9MY�im� e�&����恧
��M��h<*R�]o�-���D�d�h#�R���4[�AC�gh)�&l��o8�
Z"�ñ�
(v�[�vro�۽�s�<���|Q�"k�2�T͂y'�1�zЬy�l�=�����3ٞ���VQ�[������w�3�t>T�]7o�z��A�`Ź��U�*C��V��OJ��DY˫ۯI9{ƽ���7�5�\���Z&�Rv6�S��r���c�r�3�M�g���?��r�	�r�II�W����*7Mյr�_A}������"��+�Ȃʢ`�� g�?Ո�=$�O����F$Q`�N��YV�P_�Ϯ��{�����l�^K�(�o>g�ޖA�$�nY��A���d�er伦gN;!r� �����쳮��=#���QN�0��mhC{Ӵ� 0��mhC�І6����ZVT��u�1�(�VR���\/@�u�=As1�6kLa���	*�t�6@�����k2{����X�skGc��_��o�]����Z0�$KXN����V�K���-� @�E��D��H`>_A3*�sQk����������M�����V*�kn�� �x�X��Wg�i���ũ�3��С�����sķ���;x@��§����}�,� �����_�
��'�/ ^'�7r�o4u߭�g�U�_'i�߹��k�:@d'2��`QGR=�,���2s����#K�1 �.}��@@ܮ&�_u�\=�+G�E�����a������I1n��,�ș��7"ONu�ˌ�\=�({�Y� ��뿆�W����&��cR���A$�/�;�[[$�O�՚@}\�X'[��8�T�z�Q�5��:d�s"N��1���%�W:�2o*WU6��/�ƿs��>�m@�Z	L�ױ%Yo���:�J�;
#vaY��`T�>+ٖ� )��(�B6��أb�����C�V��.F2�H���)+a#�9s�̦�,
��J�F땸0���*������ɜh�o|Z� O�d2�9�!
���'�s�u͘�ז;_xU�̩���y.׼J�H����ܟu�o$�-kzK-l�?:�������{�G�'���}7�-*	Pn�U��/}�k�8=��{w²쉧�&@�
��1��H�aZ��s��A千�x��'a2�"(�04i>�k"��w�X��^P=�4x��y�5� �ٻJ���!�`=І���ߢ�iQ߬��#���:Q�ֵ�}/��"U�����`�е��ؤ.�l��/C ێ���iF�����1JC?uz2�s���:~�
��1��T��*�49���Gн/VcǾ?	�-��W̾n>�X?��6�����fh����}�L��0�+u+���;W*&�{��Qr�3C����{�wM�<�+��Jw��*I��y9�`��)B�H�:��{�ǹ�]�M����{}M'3��z;��?瀽��ٙ����*=P��յX�-6��px�"ŕ���8fp�U��9t.t&��m��x�����=��J�H|C�,**5:W�F�}�K�����%f�,�ȳX���1Nr�2gL.����,+fzv����*�>+��?����)xhC�І����І6��mhC�І�k��?�1� $���i����U��g�p JL�	� �@��T�pmZ.�٥g�{TG�ˢR�Ӥ�(P��:��B��fm#e,��M©<'�3��.Yl����8Q@Ye
dRq�]�1��^.a�L �Dr�x���&l��	zV�����~�,��������7�~�:ô��&	� ֮s�^�!y?�<v��<s���c�~҇��T�']� ���3a�p��gG��1�@�|f���7��mP�w�����R%@����ν8 � �f��A�j�[o*+0�0��̊��,�	T��/`[��Y�3���ɒW6ֳ������l�hc�R� +���l�L�.�,<�)��iʹ���1,�ߧ�K"�\�r��T!$�g(W��"�����@CU!�ү�����	0@[C�K9�HXw��(` ��s�ԴP��	�ֶrRйU�b�� j�4�;�} I��O�#ywMK�E?���4#�$hF,yL}C`B���P@T@��}]( k�!3��d|ȯHY����My�ر̽�a�N@L��:�-j�l�Q�D����ZuB�#���TzA�Q�e��,��*�%�t�#�r�
\r@���Z�OJ&(���P���K�+��cS� ���̖����|������aX��_��K/!�f��n���?Hvq�k��wnF�Ϝ���[��7������=�
M'e���\�\G#I�=���~>?�R벧.��H��Qi��9��ו�'0N���x��T�ۃ�}�ơ��9���JuG׎�#"X��|!���,�J ��bA���,[]녇��� ��A�R�Ν�3	���\�(H�q��'Q<J]�5�D$3M��dg��3���:����~6���P�d��}!�*�"&�{��-Zw�[�Oe�HJ^S�l]�J��	���	+��)���Fjp�^�����d(���b�G��g��q�����ꚟ�/B5��bf׮Ϗz}/���խ�n"6ջo}�z,�����صAǙuTB��]w�o��~���+��⫶`:��* ��Ŗ��M�R�/m\���s��Q��H��e-�j1�<��lK%{��c���E{r9��XGQ@FNZK�³�]�?�W��n]/�'�_�^��I�9�!�m�1w(�p�_|$����Y������І6�����mhC�І6���֐ �4��8�a-,n���p5s�~� W���;P ������P]b(���v+�>!ȁ`e�Ė�[�Q�bc��0h��=����'@&k�90�9��� �D�9�rY����b��|��vܲ�:�c����.��S���ZVG��b��`���f ���ρ�l�`�.� ��u ���A)��9>]1��b3�U��ڜ	��Tl��w6�H_:t� �Y�Y{��%6�����;����_�s���/������(�ظ�A�"}Ϳ�����*>��M�[��B��s�^�ڧ�K�lERB�x=vj�A����o�P�ޏ����! ����{�p鎋����F�\�)��\,��������5��ݪ���cX/V4������Q���%�W�ԝ/��ʟu���d<&�s�\�u1C�j���>��S�5���G@��k��J6�*@��n[?���ԩ���o6|.q\�A���d��$�/r��c�Ή;�)4<$��:_�w�f�gRܨ����p�4Ugb�؆K�?����z�d��Z���^j� ~�\XL6X,c,���O-a������g��1B���!yn��T_���um����^�^�9�EDR{ V�0$IWr`@VRy3_�S�X�'Kx24��������s����d
�|���}�%��_���/���/�l�	7n�g>�y8)���������=H3��>>�˯\�Gy�8�� B�VY�H>k�.^�����x���h2����7��g/�׿�ux��oPv�����R�m�� �~��E6�鷊b~��^j:V���"�L@� ��9�{!j=q�m=6�"�c��[Fq���l�:��(!��%��Hf�p�|���3���N��uYJ�G0�D�j��>�n�w�
���3��P ��,��Zv�@k���ϑ9���Z��%��L��C�����:s�;��/�G��_�9���=�����L���S���~Z�	ԣ\���f��_�NY|���y�"���+��V����������Jg�i�o?w��z�F�S��??Xi�?��~>���s�/�t�B�/��m�Qz��8%Ԓ���U:��f��� �$; /�A�$$�&�ݝUJ0U���%~�H3A�=2o\�Պr��K��������ϩ�y�S�F�yTJԒ$}�&��$���'A|��2=��mhCڛ���mhC�І6���ֺ�˫U�ڶ횶�$���\�˂���^�g �K���H�+pB�Y���'�6�d�R?����	&��A,��-�6�2L�)����)S��Qr��䘂�DcP&K�V�pDE�C�&�o"�e���5+� ��2C�" |lmn��t���ك��{X���5�3X�Q�.o��if8�_B�
��S*�BDPx��~�/I�`��,{ݟ�ͤ���H���<����#�`�K�,֬��G��\{�X�e6��g�$Џ<o�}��^�����H��A)�*�����S4��
TYQZ��u:��}F��3%	�J�Hr߅^=�پ]��g�X�B9�X'_��l<����<��W���ۇ_��_������� =u�[��I`�}��!+�'����{� �;�������\�v��v��mOON���-8Y,�������������"`�,��[7oP=퓓x��	���%�[&+��:��]ҒQj@ ׷׵�2���πg'�K�.T��r�%� b*�)}DA�.J質@4���̺��HӠ��~�}z4 � Xsf2͏(D)���Y�E��9�j���&��f������~G���づh�A�}U^�L�&H����f����D����I�"���zݦ� Lb��R6E�c#��=$�(�J��j߈�]̀�<0�Y��f{`��}J��@��(�3�����T����pQ�7"����b�?��:�Q��	����.<�����O`�6ǰ�9+���ʕW`�p\��i��;��ƽ����s�������8w~��Jz��u�f�T.�1���~�~�_�K�?��?��}rrD������ɵm�u�� {���E%�Z��Fe��v��粟O�y�w�o��_�I
�	!Aj�+�*���}*�$�j �mQ��L��N���?.s4O��xtt$�a]�'���B4
&���
<W`2�$x'��~�}�	�
��"F���X�9Q�,���\����\GWp�a�������@h뺎���SI��d�Y�1�Q�:X�o��(٨�3*�D�!��%T�$�����ڷ��گ���u#Y(�z�8}v��%t�������^[?S7U��?�����ͯ�Y--���4O��H.z�[�'�Gb_$� ����I�Lb�5r����G�ř�6�`���6�{<}�r���Cז���h����`���K&�
�#�����5Q���>�������p�՗H-E����>.e����_�F��ɉ2�1�ad�����chC�І�]��І6��mhC�І�lM�P��D*�K�,w��k\�cr^������@i�À�%��3����\�ɏ��F�5�o�a� w�`1g�P�=٥�'H�������9,�(�$��n���ׯ�?��߄��k��Z�T�;�(}K Z�c, ��|@ 
X����5űv�|>�`m��A� � �[	�a&H ���`kTN"�����6�s0%�<X�]0���3G	h*A�O�#���Ѓs��
�EP&VC��w���ͪ{~a�Q����6ZY'דB6T�Qw�^�� �o�[>	���WC�0@���j���@e���U�����it e�����]�e<[^��@k��Z6�r�Ц{4��F�_�	U0���.}�0��A�,V�FK��6�w�Ѩ��1L'3��_�o�ܹs0�Na<��Gc�gAS�?BL���/|���o�+�;?���~��|\�����S�U�E_��#�;��)��Y|������Ǟ���[���IY��[;���k���S"uD
``9�]w�Cd�J��0��d������IM�P;�A�ɐ5{���~�ߗ,eu�
���@���Jn!�@���-����́�3v�ݠD.7U}²^kpPל�/RƸk���D���#ya<�H�VN��2�8�Q@L":X�'��F�������hk�<�%!�I�?��xA�4�=��#�'=CW��֮�%�,�=t+SL�}(�f�x�66���Q�0���l���ż��	�m��h�&B> �@d[�q��<�Y�M������~���^z�T2p�C`�gh'����r�%�B�����˗_������+O��Wo¤������NY;d?�U(p~G��}�q�LY����Ԁ��e\�_����ȣ����d�x������ S�sgt��D����4(HͶ�c��_' ���h�����K��1{�~��e;8J�m�c�VD0�.V�:����a�*�_�|nll�����9B2�^`�Vh�7�����7\w	"L6��_��Kt��{Q��1���%��8W�@� ��_�Y2�2�Rrw�d	��_�N�q���=�T-�9IY�/�_�mͳ_��D�J�y���؉C�/�x+L���v/�^��d� �%�[?ݚ|��y&?��_5Q�lQ:����,"ղ2@�7i���Z	�WBB��/��׾h��Ũ��:��P~��sèe{P;�2�1�T���G�w�`���Ny�l��O��sş,�WW �3v���C�~Z��D
�[ʶ�w�>��76�p�����W_)�3WVY{�#ٿd�u	�3Q��ŗ�`�����$�����o�C�І6�7E C�І6��mhC�����<�L�d�9��X$��-C��#�f�Z
^sn���G%�@$���-s^2�%����T渠gg��4�[
�J�펢�ch"�1N��w~��~~�W�j�Rǥ��"�Q�g���Hr8e�)6��U�`(��
 �a�ϜD�T�q:�gҬ���0v8��%��J{�$e�\]Ɓ����Cb�Ь�h.�ʻ��H� �{��}8�gLu/�%��Q.�&C%+��`�7�e��h�����ۂ�,*�Lҧ:��� ��(κ<����h�ql�5�C�놨��
`���"�
"9��Pfwـy������6�6��<��fUimX@���֐�+r�`��G���O��p����$m��<��>�d :��������w:����<���)K���~�5)3}�b����&��������������L���y�����^���K�e�Y�S� 8����cB�e�3I�2�EYĔ6t|:�C%�#���֒�gHuFe���,b5o\P����Y��F_�%\חg	bF@��➥�d�
(�m���FF�J*�b��^�Te �w�+p��3�|�>0�����R`=��|����B�I����s�FU��������(�5d_�%.Q�;5��FHQߣ�1�	/=�\�����\@N��d��u���p���{���g �K���oXº[2�Ǥ|��?�q���h}��垻���_����������n&�5ݰ��h�٠�x��8m�4��c���aM�7~��}�g��?-C��1��!z��Zd/�s&ZMx��O9{f�nR�H��-KZOAԌh�u��G�=�d��J�?("���Hf��.8�.�/r�M�!���S��JX����n-=J��$�F���[7\��a�U�Ѝ8����_x�����;�y�kɀMZ�A,�}B_]�Gg���Ta����^X����W�lh�;���J�dg�r� �m5��62úe�.�3֓P�W�YQ&7]�1��WT(�`EM��]q0]�9�ˉ����ê.S��y��Y���ܨ��z��3���\��ͷ�j�BuR��	�=<�c��S�DeRc��X��*�ϏG�we�C�#�!\F_��ϭ�{��]Vv5��$P}6��g�JF�u���*���A�$4L\,����;�k@�n&�!y��-�h�!�ߺ��l,�ؐ*�k}����6��mh��m  mhC�І6��mho��R�-��c1^x�`fT2�QA���M��V6@��9x�Y:Z��%�D��(=mr�JI��2<�B���[���ǄAu����^���=��.\J�U9���.4��3Ĳ��b𾡀4�W%����٨z=��=J\��R�,m�l�k�-P�ΐ�������L��k|�(�)�$9�A&�������L6����v}��T� u��爒)j�[�#G{T��V1�l y='�g7�h	���;��+B�|7�ǚ��G���f�����e!�{vXŞ\��q�n��䠑�+����Z�2�+��"Kkf��Y��k`�/�r�����b�ԌR� еi`4����G���o�������G�9#'����'66f0�Lac�Ak5��H��J2��C���tF��������~���+��� ��Q65������WI 4��wrr
a��k*�������-�\��ng*�e�;U�۪����X|����jl:���3�9<Y��H�L�F����T�����맑�i�3_�Q#2M2?��?�w[<���*H�@03ғuVR��Y� ��� ����~�۵I����9d�E4"������$�Tl)؄Ѿ�@{4_�d"�J����f���,��=�N)X�f0�B���N �Di�����3���qD�v"�-f�on@3JD�9=]�
M�n�3L����/���=�"��}��\#�S���C�8\#{������;1h�0�|�F��� %�������:˼��rM
��������Kp��6�ėxm�@�-���|�UҨ�����&�YF}�:g��T���Q���l��|��g*�g��}�׀۰�ˬ��e�}��>�x:)s�E}l��y���}����͂�I<J�d�CCk*N�Q}D����H��q��_���T���'?�T4b#��ԥk0�B����F7Vv=���]�1T��I�B����un유6R�\7b��j,<�ӈ����נq�k뭓M�g)������뱐���?����w§�����3g���E?^&�˯��'c��NZ3���$&,���0����:�?KX.V�/�?R59��3%	�V/ӊ	��Bߖ��#\�y.�4x��\�o�IY�\��	Bk"B5t6���'Wו3T���)C�1���#i}��<��_�E]IN��g�6��mho�6 �6��mhC�І6�7`�.���.{ ��4��"U0��Y��,�¥U��s[�}BZB��3�)|�b�
Y�-Kn{�`��?��r����S��Y��<� ������~뷨$��AB0 �u[%H&�L���H���%�-�gVt�\�5�)�Ϡ�8�ɢ� c5�H��m{ ��o.�b����Oi@]�Aep����W5	pZ���_��h  �6U�4W��̖z�A��Bes��6� =�X��F�z�>� z�bw1;@%A}�ֶ��T~�g�J�T@@?�ن��[h@�{�����l�`��W4�~��y��u�dX0|&%�H�L����,��)�ϫ<���c�5��/N4�)4�a����R����c<+-���;��ַ�z�!" (a%����3�6r�{� �B��چ��/�{�����>�.]�g�L��f��˵��ʕ+��SO����-��G@b�D̾�ti%R�l�HVR_��	�X2 1k�?�'��Ub��<j��n"� X�ʆD�#�&.� �H��T'��)Mb��z�z���:9��(�<hŎB���HFh΢Nr� u����#�+a��1��#��~BI�1�1٠�r���\Sl8V������%��;ɀgUH�_�l� ���:��������3��̒�-R��R�a�py$��|<���l6��0�S	 �P>99�'�~N�.]�����e���I�.�c`��t��3��ـ����� ckh�SfL��h�Ip��1�q[��ɵ��5g0-�1��J[X�T��#��ؒ� �1QRK�$��іg�L�D2���5z��-��7��`D]k�]��H��|�5��<��L)���캿 ���A]U�6����Û��V�[up||b�N/�`�K$ɠ{Z"B��p|��l�lܞ���p�q2�D���$�g�z?2��l��_`���Y�/j*1AI1�Y��vֵ`l-���Gy?C�1L5�=����_�=7�_�n�]@�=@����Yk�C��>g�mߕ�7��lV��'�V��墴���B�~g�kW=�r���@���:��m��2�_�)I��&zL���6ZH��V��}�ѿ��^x�GR�:��~�d_?.3Q�N�dΉJԀg̪��MI��r9K�0���֝Y�?���㝞M+t����L�!}�#[3���Ex�[�F;��s{Ќ�� <�R�UM�?b)�:"�S�U�-�:���Yu/�>�P�O���V*�ahC�І��i`hC�І6��mhC{��i0����R��A<i9���b�*Y@K�j��cQ�;�Ph���ھ�28��F��d�B���EHu��)P�h��)���
�_�_���s��4�V�?�Z�kj����GR�ف�qs0S�h*@R�k��
Z/�8$0h���+���a0�k6�4y�7�*�$�+�`��f���~)�k�q.�Pg�����������f�Vfi�8�{Jv�4ַ�f�kwFMT���
�šM�wNJ�=�	\�Us��٢aN
Fj<�f�KV(t�lAR�ʋN�Ў6}L����kk��P��g-�|�O�$��4ӱ�5�%ͺnGg��P�"դQi
^�\��T=���l7} @W�d���=�u^�T�1���3�iM6h'9[��+�Z�Eq�b�TA���lJ�ñ�u�f�+�T]�������O 20�1����),�ʰ�Š��Ř� �������؂/»��n���q����8:8�1E�>Ө/�Q��UBV�$	�f� �� ������c��F��u烒:�ZF��б/�m�l��(*.x�(�R�7R�؂sX�ߓ曃q��˵�� �e��V>�"�X�/�2��!�r=Y�l0J�WA3�5s@	��ޡ��zJ ��:^Q�J��R��=uS�	~��Rכ�����_�6��l�*�����s$1�QF���6̦3z{�����)<������{�}hGX~��H�L���}�������;�ТoU�pL������]�'�}
~�>��'���o�Pâ�9�k��@�	�2�;;;����\���������}�۲/�9@�1t�`&���!r{چ�	Q����d�ZR�<��x%۶����7�/�z���gC�E�@Ku�J�5�/h�{��M(]�6r������/�?8:& ���M�'���䍴�<\'ݱ�z 	L�;�@h0��� �xGS�Ճ >MJ �����������������I21���q���^��}�N���gL�z ��ڷ ��O�d����T�5�R/w�|ƩT� ���P�{�
Q7�����%#i�3��O���N�xU7����s�:v>���Cu��kBUx-��B����_��`l�F�(��2��χ�{rrO<�Mx湧˙`��{[#Z�"(q1�V�W=��F.���Z��:�ڥ��OK���)YH��G+i���U�T��Dj`��y׃���M�X�@��؏ �	�YZj��9��2�����~��'v�ı������6��mho�6 �6��mhC�І6�7`�1��bR�a��B�u������?�	i`[[��~.�Z� �d�i�/h�XT<cR��R_"W�sтf���db������¿��~�x�g����%��,ϟ:�:�ę�Q��2�\-}P��IA�*K�;\��2��z� N秠�rƁ�`!ѵ��dYC��-'���XW�;��۔)��_���v��{����z�����@��>���@�$����5\}]��5�_j������� H�ׄ۟U	 JV@0���S(xـʣi"�k��0��g^�h�$+�������=[��l�e�������H��`��J	R;�~x�,q �m����lU;�Lz5����r�/�GfR�M�,����������u� :	�˽�CP��g����MR�hZ&a���7(3����,Ezm��)��e���i�0�N��RG�}�{��c����I�\�J?�a� �/�PUK�W&̮�AP�g&](��9���Ey!��B@��Mǻ�=N���W%w�k*o���Ł����I�%ɺ�dr�h������$@��g4��Ğ�Ӎ��5P�e <��_4��Mj�U+T�KND0���T�$���x�����ԗ�83�
%
��������~��O���lg��࠲A���l>�5��B�O|)~Ao$�!�>*v�^�`wg>���א��25dS����ry�;�	�����;.�<�|6���$�?�����n�,����|
��n�o����C�L�Aߊ`=~f���������r/�p}���ƥK�د�u1*�i�\�mh��T��"G��͉ ��ҡ���"�� >�a�����
u��/ �	t��er$0xxmf�2Z_����d��8-���׶�6�?�R�ãc�p��ɬ�/�����@`�~�ߒ�Vݻ�3��
�o�5.`���dۺ�U+a�gr�����3��K���ˌ��%5y�}L�^{�z��l�8��y����j���9����$2��O����J?��h�k������̽nW���d��]%�l�I�N���4�:Q�<�{Nf�,w���5��v�u�o�vk�Wc4���og&h%\'��V,ʚ��Q��TCTy$P��sțV�&���8q%~ֆ֟(e�gW�i����UiP������j�~T�>)�>.�+�3��gt>Y,;"@��;�֣��q��E�@6����J������=%��� �ې�ěf��<� �І6�7O C�І6��mhC���mr��իW���iC�z	�a�j]�A� ��1I�,�l]p��� ���`(I3���m���A��<~�@!斫��D�����G����&)��w��f���>�U�����qFbP`/sp� E�~Ct�� >V� f�&���?AD�}B�Z��|0�kP�5(�n�a�Z	:�,7R
�i��Ҵ{u��_�J��\՜B�*�[=4�L�ȩ�)ʙ�L3�"A^�����?�	�k�9H�`R0��+�Ϊ���t��6�s�ߍQ���"SW�1HVh�lW �{v����tM���UK�ֿ'�)�o�e-{Ɨ_�š��~.DHun,9P��ߪ��z����Aȳ�Sx�_#��\���n�d�MYϜU�$���m�^�����я~.]SƿJF�_$ ���F�㩘܎�s�#�y�9�Ď�wL7f���j"{�{��"=��U:_���%�2����VI��S��W��QB�nS����c-o��a�����`u�1���@p"Hv2rI�t~=�m7VY��gc�#�d����Z�D�h�n�zy���	��0S�{I�0U�U�6"I��S��?b�!7%� F�J��#�b۹zVu�ԏ��U�j�=a�{aj�J� #>��G6b�����D8�YU5DAR`�U�W��|�mǰ���]�'�'������ʜG��������vwwY��2��~��|O^���PV��t׏Hj��+�`�X�x��d�L��Qy���&�>���e�^�Q;-�[��5�	ܸ~���77���OfR )�p:��u��W������%�X	�DA��|d^x��b�©�~P�?K&;Ьp�OK��sDæ�DF��P愈#��z��0��L4BۜN�Dl�=���5$=9YG�	�:KEʐVRS�T������=�2/r�~a$��1�^����O�?\)T@�e�gUL�W���_g4�e��G�5����R �Ϗ[��Y�Y��@p%u�\]RA]�S�j�^��>�z���_�z�5��S���[hH�ߪ��.���g�vP_R��s�Γ��IάP����V�v�=�Ԇ�}����2>`��>���*<��qy0-�Ag$�+�k]Z�,t�Ci�NtHrvŒA�o��E�=�6�αHd��.�s��e�~/�u��Pze98<�o�����w��Y9�dX�s���)���ߐ���8B'��u��2T܅���ze���gh�27��mhC{�� 0��mhC�І6�������������͕W���r�� 6`��'��t@�)-S�L\�BŜ��fI;�r�AA����^7j0,��M��诃�h�`�|~*��K�C}풁40(���^�X����W�I�c�0�Y򓃚Q�)��D�9::�` TP��T�]F�z�:�* ���,�,�%��:����j�Yk��>��
�Ɵ�̀�ԏV<�ꓕ�x�gVPMdPq�	����#w�n�E��U���πW�P������ܓr����s�LA���5�M��e��ܛ ���>�*�{������e��dΩ��j�6 ���m4�U�$��GSg&Wӡ~ ��U���=oח���U���	�#$�
�$���!�9�_�(��������w�r���-e���y��r/���ڑ�H�>�̳p:�ë��
�;[�f�мM'3�q�&�fNf3x����� ll����s�_<�t4f�PI#ns����m$��`%?Y�z0��0e'�@��l`��1�ٔ��hL�v��kּ~]�b��������u�`�f�s�l�S��A��>�֪���}~�{00@��^���j��������GW�T�q��3�u�u+?I Tp�����%�X*���κ��u��Wu�\�Y�G]�F'�U ��p�3��������*�dL5���n�L���F.qAY��}�e���x�ϟ�����5�뚕���,e)��6fSx��Oh��/	�»��N���`sk��T*X���^}����_�??��~���׮� �o����G��{���
3y��kQ�XgQ�P��j���(f�h��.��x!�4���V�Vy�
�Ϫt��5Z^m�R��f��OB��6�eE%���*G��g�'V:(�~��-"-�}�ˤxTK��}�D�TH����F�0�|_���qB�W@Pb(p��*p?䀣*�����B����G�\�N��9�ZR`�A�:>w~au�'��|��Q�HN�^c��������LN����UA�]t�Q�/ =k�=��?��;���*�4J�P�lKR_�X�\��B	�_۝�oU���&z��=O���t��	�֗z����u����ǵ���vF��7�߄�t
w�{�/~c�X����,�E��(�t�cVR��ב�d���󤬒�Jb��BC��>�J��A6[�������M4L*m��1������yS��![jK���ɿ.'��Ʈ���f*�汬7��<��s�_;ju�:3�C�І6���6 �6��mhC�І6�7XC���R��r;j�M!�:8<#K�4� �sk� �`��_(��@`����&D�,�����Bk�Q3G��ə�\��* pr|�Y9B"H�[Τ��=gC'�Y��r��Ϡui��Rc���p-��J���`���%�%: �\����&�!3�����A= ���+����ϖp\Ƀ� ����4�ZЫ?�%Ӌ�|[+ҁe�i0_�b�Q��� ���8 �*�����N�S�^lu"�h�y��Ԃ��u���5u*Aff�ào'��
�`.�k�7LP���n7��R��eQ�e�L�"Iֲ�M���׋VP4�%�6��-ڟ�S^����d�b�=����:�:����e�)�����0_�%�!x�-_D�.I&6Jׂ�9y�_���Zj���~� ���}8w~��vxU#H�����1Ʒv6	[KP��k/ÓO=	.\�/|�/��O>�/����m89=���?��'����_x����1���s����%��cḐ�8�����>,�X������M�C�Q��,�
�����FW@q��U�p@������l�o�P�
'c�zP������r'�!t�C2��F��ā&y�Ϳ�AfF�������&��T2@���̦�>u���ˠ�:>[�@�1)_t�����e�g��sƴ��h��:�B��9��ul�`���t�E�%��z��'ŧ�-7�oퟻ@�>�� ����KY�������uR����*!����^�q��h$�}�������<��-�ڣ_+���m������H�+g�_�x��z�]�Y����˗I�g��%��ނg�}�\�����5��k��T�q+cA>�6�lc�#'�{f�{��ƙl�)"��#��#@�{*}'si ���d@OuE}��m+����:�A}��C"[�* c:��Y�ڵרDC��]�� Z�2,���I�%:�Nߤ���FI8��ah�6Jx�3�-��C��Ķ��?QJ!��	�G�q�ޣ#w�����D]wQJG�^��k�<��� ����Y�m�OM� ���~��BQ�PyF-W�^�o!��}I}������<
�4<+pŮi���9�	J��ٲ���X�\�9e>K��]'��� ��1:�ϯ6�!�����y X�?���Ήۀ슉��3�=���e,�9rF�
о�+�@�D���ف��M�����S���>�a���L���Z%EI�Kppi��T�I�jh�K�$T%�i@2B�vm%�Sᙷ[��ز��m��D͈�|��2ms9���7��.]��tR�vZ^[K�d�'�O���a�oo������D*�yoP[�І6�����mhC�І6���֐ �snrȔZݥ(��D�T����fރ�r���$��ڼM��[��0i!�1f ��{I2xh��톯�
"���Q3��e+g$�8�xpp�����dP�	�%� /P���(@�q�c
vb�]۴t�(D�MFZc�6f�@��`�:���C�M��h�L���`�����}�%�W�GU�����ၑe�93�Ug��7t��d�n Y��	,��f�=�k$���x�c�ۿ�����[�vv�`V�^�IM�|s�d�]�ޭ�$�L@⬯�u�s^����b�3I�i�ǿ�]/t]�J���K���j(ӊf �8�m����Q�V[+�PΚJ$KF1��Zs@����Zǜ��i=��ì�F�I�]���SϴN���3^;��'�u�$8L��!��D��~�h� 
�G���st��)�[�:��C����ANK��l$��I�AƦ|�����O~��`{k�����=��ف�����JOX�9:<<����W_��|��p�=��{����|�K_�E3�\��O>S����	���qTX��:��3�<���)������*rH�|���;<<��}�s�\��J�2��D��u4s�WFV�P�#`8$^�8��Q|	��ep�˝ /��!
:�myV��V��l��e%/$K���2@ +G�(�Y�#O+VS�fQ�X�$�`�I�J ���j�{B�~���
P�N<?I�)z-�M�'8�S�Bpu]�Gw�� �� ����������Qx`��eK#�o�d#EQ}�ȖHz;���3��ɁH6z�r!�������o�s8<>�QY'�:Qz�'(?��s����8&�QYW'�n�55�Q;��>�u�����r�<���
��m�կ|^|�U�ۻD�7>��/����''���<T�4��-�z�"�m�Ôm���`�?Y�?��ք�`u/О��2�3J�/�e���^]YϨ@���|�#!�/{������^Y�ʎ*���۸�=/n|�#ී�D���e4�%�s����,8�`�&ۛ���3 �(����7�uRP`�	PbnY��!�NT��ĉL}�z�I��է1�"�>��#���W1�8o-Oj�h4��_���d�u���LU���wN�O�/��LZ�t_%�9	6�9'J9�3f��3T�"A�eY���|���o�*���N�c�G�\�G�J݃���^���Q���VT�2��)�8�M��f!B�Z�;�ܪR��iZ��+�:��𕂁�3�L��5~���s�T�SI�V����L��r^[����6�F�Kހ�1P�8�z@J���NAc���o�2B�~�F(6�0$8�Q�c�l�ᘈ�c��:j���TS�z�#_�)�+8	k!Xf������������X*%$���<XN&�!�,x�����$"F�H�І6������І6��mhC�І�k�4$4��+�$�G6YT���>
TH�]��-f��GI�'���p�&e����(�0����A�2��$f���vL�)i`�S Yp�f����%��+��Ԡ�eq�[��'���v��1�`�:�������KX7�y�5���&���ݘR�Q#w �єᕗ_aPǬF��z�f�^�8o�9�e��5sV�E&�����ͨD���T'��H�:�� �f����\Wl��W����NH��!�jtoo���>�#�я.�qI�!��8I�3h�;יU��I+]��Wj�e�������Zܰ�w"p����Ŷ��Y���s
�F���A��Z'�T+�WDx�:�"O��k" 4 x��k�s]n0��D�~h"tZ� S��	{>)W4\� �T ��σ�"�H�:�3�NCBsGʽs��H6�>"����q�1C�d~L�/}�/���k�}�dN�@P����Nx�o���M� ��h��!�R���>�N"`��|�2���K�����{��k����}� �+f.ʺ�g^��B�srxnܸI~�mG�<���͜%K��
��ŵ�1��������,�(�vL�*�v�S ��r)�A�I��D�l\ʤ��}�����Dhh�T���6Ѭd��#�c����dН��J.���b����<&��	)���2g>�l����u1bvB|u;��e��&����Mt"@�l�+e�+9m��7�F��o��*��^
59#H�L*܉�;���Vj�a,~a�p_����]/W}�����T����Q.%���ƀ��-�5^��&Ra
~qV�k��.v�{*`���V!YgT�=/}!���1���>�c���g����#.awn�:��e�o�.������s���BWƊ��Y'�C�v�U�O���v�'pp��UT� _�f;(�c�-͇���2<Q�0%'�`g�I[gL����� Y�|������v�ˋ�2V��'�z�&-i��e������UP ���S��3���(k��=�2\���I�*{#��[ş���/�ի7�����y1_ӵɟ���zAc�^�{���D��ǳ˸���K���(�p:?���-�V��R6��n�&�h�X� %"M�bҚ��|"s�d6dr�W<q�����Tb�ZC'�i�06�]y����:#d(���S	�S�+��D����s8Br�8[�:SR���� G5�3���^n�S
�f"�LA���p~iE�(>o'g5�����]��"Rn յ��
ՑǻI6;("0i�ȐImRa]�-V�@!=�oM���*!	A�gų���)':�d� �� \r�&�r#�UR�B�a��(%��'B��_����5,B�Ϡ~|a�R��������+�U*PIKg)�Hm���|6S�D~1�i�L��ψ���\ť�X�T��J���`;T(��=[-�0.�Fٜ��o��g����t���k������%g��.7M�j mhCڛ���mhC�І6���ؐ���!i $ '�;����@/�\E����9(I9n-9(���������������C���	��,�נ��hc������78�����0S��Ѩ���!�_.,�R
 ���fp��U��i�L�''��SO�+�\�'�Ͷ��2lL9���NF�K��K��K/S�lX��ܹ󰻷_~ނ���<��V��<��7����J���0�\�5��D�@�aCU���_>+�
UV*��DQCу�NR'����.4XU���o
ْ�p{1��~�$Q3?�����z�m����/�M�p�Q[ƴ�v���٨*��I	��8D�֑��� `����|'���bS� ���P���H�D�;pf��h-U�K0[f\�^&�M}P��L���KG7TS6�����!�Ϛ$�M�y�Xea2�P) �Z2A=���%ؿJ`Ē5�-"��@�[@�;R@���?�����r% M'�,6&%�粖{��ɧ�w�y\8w�l3���	�&�/���b����F؟����Cz$:`M[��q�Nfp��N�o@�6�R�����$IS6_`e�uf ����}�;H�!���R|��xo�E�(XPMne�����K��7F?�$``J���U~ @��s�Lh/'P�z��6��~���o]+�Cg���M�X�;g�F/?@�]�;I��ޖ}@�6-�P�Ť� ���7t�|���8��ׁ-]'6�z3�*9j!W���Z����P�o��gx#i����WM����g���t�L�N$�3m�/��RY?S"�����˯w�I�mr'eQ�O' h���ׯ����(ϟd����'�ND�����a��q}����ǟ��~��'����~���;��o>	�s��݁�������~��� ���������t��K�y/^y>��O�L}Gd� �S�MG_C��Zؽ�$���G�Û-���{���޷��弰L���~�S�-���c��2��Zֳ7[K�������#��Il�l��6FY�8-~V�Y�~Fp��j9o�[�nmN��Ȋj��Oh/�����R��V������ZH�B q4����GD�,�Y�f�Z��9l���@A@���B��5� V�O��ݴH��\�I�~�D+W�?>>%����&����-R%X� �������z�k%�'��1	V�a`��bZ����|2BE��dY>o�6��8,`4Y�_Krf�9#ж�#�P���(�a�8���^�z��#�ub�K�`���(�(	 ���uL�J���-�̡2���4į�#�VY]RT|��#�'���i���:���FVW�_�5�� ;դL��xg��Ld_H
Dv*��2T=��{*��HL+&J�~�D ܗŖQ9�擓#Q)�t>��%!���	)YB��\}*���s�W���e��3J*0����g�!�z��a?��٩2M�u��}}� �b�͈�Z֓[�������rbm�y�1�_hθ\]yC�І6�7K C�І6��mhC��� ����ɔ!$�Te΁�TV+4s׃Z�1�����mJ����l��s\K�kk�)X\��T�1��6��accn޼I���:
"b����}/��5P,b���������}&�	O�+��1+��>�������:�}�-�N
�r��1��/��PĬl�j�d��	�Q �$[�E k[gT�݂ҁ�!0�ڶ�rI�(@���d5u�3�Lr@�2:
�BkWװ������تsWB��G�LdiǓ�)4L ��@��dC/@f�X���m����Y��?hl�A��EQ&�,M���@��B�Ќ3������~������d#��MNW�O	����J�U�u�g�
�wT�BAF�$�~~�fr��@ZG��rv��wiX�%�G�|VA���}�qo|�Q��Z���&�o���A�[�V]��,cZ��� �/��{�)x�������U�3�(-��IӐ�ҺLJ*J�ؗ����7�����h�z�фJ| � k�� �$��
p�>O'�G�A��	P)vLGɒt8$��ٖ�k�tܑ�U����D��9�_K�*�	���u�5��
Uۤ�-�:zI��A�A�g}�`jF���P�U���],�AJF�����~�u#�]e���ek�I yxU��������T*�}�d}��#�x��������ྙtns� �{�=���W�QbN\��9I����*��l]�RP�N�[a\����.��W���ί�e��:�+٬�O>��#���GRY�Z�:Ji�,��k�S?��HD���K���0�$��\�
_��G�����?Y��"�v�S?������l�g^��[7�[��&<���p��Ux�����IE�#�� �2���W:S�`�Ȳ�*�ķ�L�D�a
��1dT)��MPb}c�� z�IT �l8��V�W��(�&���������S/����<p��U�f~rP��F�I�)	�OOak�I {h��5��(�8c�T���'Ȩ=�:�9�}����NN��;�,�zY�����2-i6���@�٢��^z�e����b����''�:3!�9t/���W��0F"���<O;�6�Y��x�Ә!�@���S���ܷ��Eu��E��=Y_~�ĩ�SEh��Av1ƽ@�]�>��l�� �^6B#��J�Ki8����#&�!��������	�Q� ������I���S�-����U�d��?�((	��vz�k�\H��Ǌ�#E�p=F{�d�Lh�1(���ϖ��X�&ٙ�N4�\�ʯ��`o����LXuD�gN�$�=�#@Z"�EQ)��Y?����Y����R;�������-$��1^��sB����]�V��I����d���	?/DU{В k)%�jW�z^�=CUz�dF2kb���S��~�U�3.b\or�G�,�aW��)咽I��JÀ/~� UQd�q%"e����!~hC�І����І6��mhC�І�k�cK� �ꚪ^z�,�P�*�AP�q�;�'F1�?�/`#������!�@n#4�t�Ʉ�KqG���7YN�s�nݠ���b���I�Rƛ�9c����
C���Ou,�A���M"lnl�T�׮����16�J&��=���������s̘���;�/��"Iȃ�s-:}��!��Ju�{0N�S p�:@�����ކ�x�%�pzz�嚂*[�G��넼����"��$�_Ґ@��z��x!T�vN`�����z Ŭ��t�و���gKΡ=�SɀN�{�H��I,L~][WqY'�G�HK�1�gj������� �^�IQZ��$ �,q���4ߚA���5JĀ�p%�Tg�"��������lk�Ň�ϸ��H�#
�흂��� �b���W \	
 �RC�2��ͣ�uE�=�L}#r�P C8�[@��^�Z�J��Y�<k��0Ws�y�6fL`�Ll�p�H#�h�(%(���|����N��OMgS�)��)��c�uR���;R\�	����rѹ���W�z�R�Ͳע� 
�� ��V�[׆IA�L� ��9��7g��3��t��;�MbYJϰ$��ȟr�f\�og'�t켦1>F��щ�;���3t�^��Wzv@=7�� ��D���g���{!����w�T2�fWF�/�u'(��~���N�������F�A	�S$��s"�q)�Ӳ��
����Z�����6�+���nܺ����=��������9��F ���m��}��6��H��[��֌�pr������:���	�]�.���Ӳ�/O��J@@y�����y����FQ�i�F�bT�(~%�J9,�#&?0��(~�������i���f�㘳p�4 J���)`,��N	(fC��O]
�7:Z*@�X�Mh���iQ�aN�mf���X�a>�mfN�xT�󑰀F0ۘQ���h�-�&�{el�@y:?,{o��i�]����|>��?@��W4�aD̀f$~���A��%�M�OM���� ��hD4�V�D�%�����:?��A׌EM��z��.�@c�`��H�b7�Jj#?S������d��������hϣ,�`�V������G���C�����|oޑ-��������5#��T漝��9'�l:��M�a_�*b�����D6����~����|����x2������N˹�ex����~�Jk�\<�-i-� ����İL����T��QK*E@ߛ����I[歛���T<lmm½��w�q'\8����}?�?e�����A��[7n�+/�/��Rɞ��mt�����RU�,�N$��W�*����GT�+��';�峬�*�! �L�GggT�&�;͙���i�A�T��2@rt����x��-;6RbKλ8Ƭ6��{��L���z^GQ�XH�{X�!�O@C�І6�7Q C�І6��mhC��a �`AA?��\�֯c���5�F)N��+8M'p��U���	��u� 9�dKg��&� �$KB&� �`�����u
X�:��o���6L�S
�7�1�D3�@�)�ϒ�Iq�5���ku�ނ��1e��������2�]t�O�q� ?�|���@"ʁ��7��?�����=[�`kHc&s��B�GǮ?-�������$�T��Ϫ��oe+1������>��Pm�)}����2v7ʼ�J5�/_~^|�%�V�	�'�@h["hP�Ժ�04g�uR#[�K�]8�ܲ��w�E��$��|'kv�Ŭ4y����m��_x��_dp�.4�\�[�:C�w���Ld�' �d���|EcR������՛��ۅ͍m��޻)�*�Q2�g�'��
p�����/�����|�˔�Ac�.�*)
P&��IVd��/~n��G�Ei\�&QN���K�n��.&rкI�0.ē�"y���W��>�/���*�~xt��sbZ�:��?B@O]��LH�Q������	�f���.��oy ���q4�Fp�|�e�AD���J�	�k:���1���Z瀠�e�;	��� 	?����+�B�l�R���FѲ� �b�8(c�1c�k-��(`�I7��@h�U^Q�C�BP�k!�赔����"(�l�K��5��%sO,�ƽ1�r���`�X"���zKT���>N����;m��R.@\��C"C�j	�ǣ	�g�������%kU�����T�DM��e��m2P%�Ɨ�eY3��̀!��lx��=��	x��'Y�3̣|F�<��f��_T�"YyQ+Y[D�����{�Я��c�����h��R�G�˰F�A�+NN��?ʜ-{���	����T\.���e�{ʮ/>�A\��e�Y<�Ҍ�0�R	�q�&9���HYVhQ�hx^s��EO�FqS��I�1"�h?��Ϙ�ތ)㸬bL�fD+}_۔1%4A��g���(d��<�=Z�)/�� 6Fn@��}�z�7^%����y8X�¬�X�h\母Z��}?��*�7��M;a�T(3A���83󲿌�5V�g�M8]fVC��7-����gR�#!ྃ���v-����ކ��0M�tJ�d�x_��МG>2'kE�Px������Z@�F2�n&�Pֵ�c��b3 V��f��J��٣� ���aB�=O�0�؄y�1�i�'ʲfb�X��	b+���xmȦ���ц��ɝ�:Ī��j�1���Ò��A�j�7����Ӕs�v9�}������=y�T���I�b����/��W�������d�Q��)�}x�[����ុ�+�������>����#��b4�A����T��Ο� ��K��?{o�Yr����mo�W{U���޻���B��l����	f䙰���� b1v`;�4A`1�`@ZZ�$�i$Z�����������v�͜<k�W-O 3-ݔ^�W���{�f�<���~�w�<q�L��p�
��/�FKK�������p8��Y��Ιz���$�s�^G���<��k�_�ʗӹ�Ic8����Z�~�nX��<��V�ѳ�ڤl�D�t</yQqX pE-i���
��Hd�����<����	�x�����G�1ڹ����~}Q�{��-U���������󨒛���&dBR2p�{�#*�W�^�ֵ�u�k_��# t�k]�Z׺ֵ�u�k/���ȑ��)c̩ѠP��)զs �e�K��y�g+��!��ng�~
���`>�C�Z���Y渵�9K7����*����<u꫰�y&c�l�t�N@3A��-���tQc������C`>�|��Eغq�I���O�}��>8~���-�� 	f�O�ʦ�~l�؄�׮3���s����Hv��X��f$;�C���/N %g:�xRPQ4�Yq��(�K�H��U��y����o�f�ط��e����?�q��yǒ����5ԯ_�Ο'b�SO=��\&��Θ�Z�2�-�g��T�����@Ҽ�(��=�S�/�&��/ʳR 8r���������)#�d��
�H�HM[�>p�F�{�䯂d1z�3��3���ex��W�;��`6^[Y`M�jڣ<o�篽�������dL��!�F� �k3c��T`��͕e��H�ad�d
����z#X��w�}7��O�g�V������R�v6�Y���v��I��i�����`/���O���g5���iδOs$C�K~�k���Y|}�����?���=�5Cµ>V}S-XD��I��1���	�B�����Z��D�]�P�|�.%�6�_��o�q.�D����@��;�d��n�/�@rܲD�	)�����3���	�(و[�s��%NjW�O*�gu��&��*���BD�qm%�P���WpD��Ր�����kQ� �ߒh��N��UT~�e�RL+�� �PG�k-a����a`�̉�:�0A���[� �
��O�^�.�=�P�Sާ��R�9ۿ����	��($Uj�������{��Y|,IY��*ֶ�6�3��@E��"�{��=ζ���t2!��� v�Uh�/\�ښ7��)=笭@%�CT%�H�7��!_�p�@��B�sG\�]9�yWeP%�'����v+�#�Y�Ii��wO]
ˡc9f�pf6�KOk��c���ړTv�L��Q:�)8�D�z�:���ߓ�^J�K�;���-Q;�h�~�W��|�f5 ]=ȫ@��V��D��a���|�c��4׾E�t�l�g=J&�1��AXB����5���r煹W*�{L�;*��Ld��@�A�e(Ӽ��}xowm�z���p�WB�m��g�H�l���� �`��B7�:W���³M�y��Fi��4���$
a9�{��a�I�Ȟ���g	Os�� J�k�y�I�6m��*�嫆Y#�ޓ��f3H��љ�"ř������^��8�D��5M	��CeeD���������G���ŀH������?DnIvs�]w£�z{�w�W��'{������{i���o��7��_�!|D"t�~b6�����~�k`����G��ں��|��9Q����U����������Op��U��˛=����
�*iZޫ��%��'15)</RY
$�t��s�f�;�cn�ٶI�+F������ýs��|�*E�W�y��o8ЃW�
'g�b7��d�;S�}�'lS�A�"_<�r�"����pU������yu�k]�Z׾ZG �Z׺ֵ�u�k]�Z�^���4'@L��L~�g0���<�G�s&��U�s1������ae�Q�S2��P�0t��4�[��(]cHI�3]so2��M����s

�tm#�_Yz:R��H2`�3b@�������3c�_i���}{9������X~Z�9"�G�J��mj��G�#�e�gN�d��2ϋ[�>+?� ���A3PR�C�c�9��[�7f����u2�Z�Թ��+X^^���p�ĝ�������B�/��/�4�1��?Jj-h���k�j&d�<�V��)P��L`�q�@��"-��6fOv��%,�ٍ`htO��eWE���k�a �À�����$��l C�{�,ՔV���v�4���i|�i�	8�g$cH�Oן7�^c�\*'Gu90�����[;�LM�pkʀ�)��W}��8+	6�Խݝ�a<���������a�b�/�*]Pi������ b��J�o�`5��@ܥ�Fep�ڦ��N�>��	����1]X#�n��H��1(��}R�@A���2E�r!~�p;*���jW[�G02
�K�O��������/,1(`���J��,����By/6�	݊ [��7��GUR����@�7 �'��@��Ĝ����r�Fj�����2��{��u�2�y>�}*�Oe#�Q�]J�;h��@�Rd�-�2߃ߞ3��}���B�[�O�m���.��-�o�\k[�������'cˀ����"��)?�󮦣#�����\��lw��S��]&�5��@D���W�(������Z��G�l«*E�ɧ��af7�ɉ�g��2`B��S�������TQ�o�̈́E��~5J�WR^��K��B��bN���1�9K�F5�V�u�%]�Ue�D��f|��'��!�i�~��Y�4�;\�ȉZ@0cʾ&Jl��H?ӽ�;٣�륥մ�40ٛ��#GI`e� `8�� d>И�2�A!iv��<���P�e��EA�Ju�5��BigH`jH���M%$&)ۃ6���2���:���+�9��w�uܶ��4�;�#<��(��8�T.'�/�I�=����HJH�s��Q7�D=�iS_�&��ѵ��{B|��r>*@M���� x�5�+.����kۗ�?\&�(���J�R⥮Y-�Ӣj�󰔔�q�D�履��#"�c��6�[T�r���Jʫ�&��q-�����m������QJ] �A�[� ���-�x�9���x���������
��Z[���D�?_s<�·��o���/�c��y��g=�G�Y+��^Ξ}�6w���&`�R�h�x��P��޶'"
�kem�ß�	�����J����w��k��3y-�  <��=��Cu�����D�]�+ ��L��$=&��Y1�Y^��������"��=Q}>���F�tr�؉�SXEdW�霠�?@v�����׋�}��N�&/];�AW	�k]�Z׾�ZG �Z׺ֵ�u�k]�Z�^���f"��ַ,���Y��x��A/8B)lL1��Y�-��m�)&�q6_���Z�}�q1d� f�̘���N&s�뙀3,0�� �����g�`�;];0 �u�1C����U% ��`-�#H6�J;sP�eVy�\gP�px����_�<D2� ת���x�,w%�du3P�2(A}� ,ᑒe6�<��������ѣ7����~�a��Kjs��=�j��ʪ���~�'���{e��8�-��	P:f0 L!���u3��$�r+�Wj3��`5J�S}v
�s�od��szN��s+1���ߘ��T@H�D�Ķ�� *eG�϶N�Y�`�l>�`y�>��r�@5)I�>N��f�^o�4 ���ϙ��!{T�@��cj5�죁��o/���q7�c-��lF}r�J�e`%��"�Z�O�3�)��}$P�`�����F��{"w�/U@`8fy��^$�y�H��l'�x���!����X�=��Q$ȐJ}X3�#T�l7y|͞��� 5�!�k��ˁ{V	h8R��B� ��y�jLT�W2VI^J�G+r��IBN��Jj1k�ch�����W�D�3۠�
�۪�l����?�9` ��eQw�9�M�))��l��_����`�?=��FL��w�~Q6�gg�^2�U����~�s2YZ�J�2H�INf��5������t��p��@���d�G]LV�[��e��ew�DRآ���:32FAzP�?ύ .����`{�Q�P�&�u�̡͛�3�k�e���L�(=�u�1�Z�>V�W�	�T-x�r�	/�"D�l������2
�j�-��NKI�A��V���Ua- �:ʒ�B��%��D�6 b�1����\��w�����}��'{{$�?��`<�|^@��`yX�3�O���P	�&�N�b&����O�s4>+�a2�Ao��%< ���߯�>9�աK�`zo=!�DBgt3��%��{����3��χח`��gu����(����P�"�����R�z>���lE$�wGP�~�f��p)�i_l�_fr�b��;b�B �+#X�8 $/�\����i��6l_>�g���P�[t�P ��P�b��?,���q�<d�|^�Lb��\���^��	�g3ϒ�Q�^��}e?��s�������+�zK�sC�tq^t� ��H&����*�oAThx"@Dj��ĉ������I�ɇ|�����-x���II���>xѭ��ɓ'a}��+!�}�hi���o��#��#��A��g>���WI)���t�A���;?���5�C�D�<)_0!��\��'�D�D�;i����T�JQ�����_�*��t}�:���Jq��I����A�_! K�쥯�����U5ڟ�rB�ks�	@��:��A���q��ŇFY�����`��g0�Љ�y;od�݉���~��$�_�ϱ�AV�ѳ
�y��G��ê �9ݻէ3��.35� �6SC�}ƉR���O��E%{&b�V���D&_ҵ�u�k]�Fh�k]�Z׺ֵ�u�k]{��ȈQ��*3*����Uh�̓h�2����Aʵ5gZܪ4:����e���W�LV�z��ͬqx�,\�:���P5p�9�J�� }��q�ZE�C�:0���M¢狂'Y���ً����wʠ�8�l}vL�о�<g���+˯��&��:	�;�%��ڵ�p�=H�"C�-C�	�V���ϪU��:�s��8��g)Q�L��w���$�W���1I'.`�>��	���*
�)B�1�A��Pv(f�G�8����HA~EA`�@48B"�^}2��e�N'\�>2x&1f�C83xh8p�e��ס?���_o2� =e��B\a`��2/�# ���(�=��tL��M�qlo����٬���>�?�c�Ï�W?�'�~Y�Y+�{�?/]�����w�R��66Fp��!X]]�룺řS�����3g�ڕ���7����j��
ȗ��| �)/�O0��7v�Ad���1�{AO@[ș�
G��u*�a�F��1��S|	~2�$���g��ڷLs�@Xć:u_� ��F�����	`�Ѻ�`�v4`��S�c�b}��Sp��9�\�*�_^;���ǵO���Ab�و��g���� ��*��̱(l��a&�����"
�c����C�J�2����>���b����~�����6������	�F�mB6P�U����FJ��x�{�u�	uA�+��ս+��4�ZǑ7Mzc�����F��5��0�#r��>(ب{~˾T�r�G�ÙXҀ �����d&%d�MI8����w�������z�\ٞ��nͼ�,����� p"�D��b�Z���'ȺQ/�r	<Am�%r��;��D/�g?X�K��ZA3�`�����3˱�uê>��	�k�[g!�@gߤ�A��c>g��=��(�!!< Q��&�k[�'t���#�y�嫴�Nxϟ�µ�/�*�>�|��3E+��z0�.f�ٹR���CC�/r�L�N���kZ?��EV%!�H��Y�xU��u���;5����~���x^�����ՐGr�>�6|d��H����Og�����{�B:��s��}�S�~���qE����8/}ɋ��-�}R�M����x��>���u����«^�j���ޗZZ?�?�����q-#��H���?%M���_H�O&��>�3i?������~R� r����"뿼<�G}�ݷ�]^c�z�W��U���~Zβ��c>'Q=a�|Ȅ)[y�~�#=ؕ���X[�bU�Mdv kD�<~�HeF�r����L ��1��m(���i�Aq?�y�9������l�x��g$|��{G���u���k}$j�]�k]�Z׺���:@׺ֵ�u�k]�Z׺�lu];�a�	� ]#K�`�e�B�C���$�D�T�h��B����sf��P���
K����L4�p�E�Q�^��S�]v��y���5y�"��,H2�v?�p���XO���[n�V�����`i4b��� ��A��� d{�b����z�*|���K�.�^����$)%�|�'�^�M��L�@嚭�����@�h����^-f��>qƨd�CdY�^/=����x�ŏPiP���<J�7���9�~4���1�`��ك+����dN�r	fi6r�l����7��հ��f�(�	�5,]?�l�p��%��hiDD�z���HG�`ٲ��Ž[P ���6{T	Z/@I���������w��}���:D=�1n[��1@��5�m�x��u����P��}��/������%v��Ri>{J4����R��=8U^�����W0�RI��%�i�6UT_��g��+^��4�K𕯼>�����G~�HL��u��$0��駟����������0����`~�X�Q+sJ�Vדd�`����*��)�p*���|��Y�R�>c� @v%(^:F�b��cS�o5��A�;T���Y�.�9�K�
os�8��2�4��3sy>m����e��4JBP��2߱�{���dnK �=��BG^F�n=_����'��9I���+�&�"�6��j�Y�A�9li_���f��R����9��J�P�����
] ֥����$�����zy?e+K�%P(�d$��8՞TE ���o	�C��``�.R{?�J�l�DVH0�
�Dv6�:!���/^�<�<~eI%�YV�����dG{"߭Y����ʈ�c�4�6�^��o��w��7�DT�)+Y˹��݋i�L���0{5�L��/$0���!�A�^Џr��{=޷1#���@��W��+�P�R%U�^�pa��J�fh�q���U�"4[��3�+���1�{Kg4U/a��?�B� ���	8��ѳ��EM)(1��2��[���xaD��Ϥ%=W�v��J��E�k+�
��MG�C�GJNuvV��C�j�*C@/��8{p��.�FUzNQ" �	������_)���+0C����X�>� ���?�����X5�+Q�-�v�
|����җ�-?���C���󲗿���g��\Ig�g�y��r��"�k�)o��v������'�H�]��Q�����zV�L��/�k<�{Z[���g�,6k�����?�e�{O��������%/������ٱc��ܩv@J�v��SD�S?Z4�g��`_(�nv*�b�@�G�YOLx�e���Ӗ����l��Vl��z~�q?��$%_;Q�(��[��u�0f�����o/R'(2<�y�Q�qr�{Σ�j��w�k]�Z׾ZG �Z׺ֵ�u�k]�Z�^�-h�L�0�4��1��vтFE�,��*�T�>Xβw*�40��3Yg��^��Z�k	0���<`�[�y�ˁ^�������]�g�`p\ "4��7���_��k~�mo}��o���OW0��S#ف����:�w�8A�1P�k�����c�8�x�S|�a>}�i&��5f��p�`�d�I�'�9���=�X���Z� 9՞w�@�~��o�x�AX^Y%����<�B5��/�>	bsm�H�_��@�'���@�f���5(5+��U"{�R���뉜�YmH� �Gt���@��ӧ�ڵkp������`}m����u��!��Ɣ�9����ӧ�@8b��R��uEp\�������lo���'<f�}Hq�1X]Y���������`+�+0J}¾��6�7�}�--Q���Ւe���:N2�%�[c�b��M��D�h�<��?�0�L���Q��+O��~���?p�F�0���	�!�H�S�����K�%_�j���2ܼ�!{��[.@3%_$!��Sii��� c�seߩU�W��g�.r��\�$�Q<�`��MP-P�i�Y{� T��E�|E&��d�K���.c�*���3��%(�D)A)���v3`�	�V �
��"H��+�s P҅WP������5��2�˄�`�H�>��yR����ހ�x��������`�c�-|���G�W��h�V���H?���ךsљ$���1��潾G�6����5 S��9mJ�S[V��>ja�ck���7�g��`�b>s���	J���	+�����s�mG	��	A�-���HJ9	2}���Q%�}u{s��؇9��s�j�|D��5S��h��s��'Y����Wj2	��'�4\#����$�K�[%�9V10҉�����&�I��Q	�m�J�L�ǧP �'iH��8�GY��(#"g�J�H�g�lL�}�O�)�]ϒ�K�lr�`p�8��Bg�� gVC��'��d�(5�Q�ѱ#�$����Ρ'�6���yi�H��ܥ���OI!K�q̛t������$��!O�.�k������8	�8�H����{/�,��$��;T#��?�ɔ��Gͥ��X�'��Ο;��_�kx�;�	G�&B���������ե�c}�On}Q��p�g�)��-�9��?�gD@�z�L�^!����GT6	����{]:��sW:� 	���W�7��A�����Ë_�>���$���� ���/�7�FsJNB����W��,�V���}B�#7Ԃ8 >��?TS��B��X�~ܫ���\�{CAP���a�,C�$��KYq�= �y&qE9���h�6�F�eǄ	)�!�U!󨁛z]�Z׺ֵ��� �ֵ�u�k]�Z׺ֵh��#%�zp�Ye�&�-��%xL�E���~�9 K��,XI�{3I � ��,�J�D����ϝ��^e@F�q�T��cx*��-�V���)���֞v
X1`R���#hFo.�������>VFb�3��C��� 6��I�[�َZ��#��^��;O�əz�� �׀?�#F���1�{��Y�r�?v4}��;�x��Ws���Z N���Vke;ˠžcpA��z�m췌k��gAi��I\��nT��Oت���%(��L��Yn�c��hx�<��S�ޏ�7C�����:��7nQ�J�Mcy睰��E����'"�hy~����S��,`kN���W	Q��^�ۻ;D"@ ��ٳp�m����=rΟ?7�o±[n������z����{�	豢@������38-�+Պy�)�K��y�Vb��,�����֐l����n{}�~cZ��YM�,c���7��D䀆��POP mS��Vl��f�j�'�L��S]Ǽs��*0,dP�M`�u��	p]����|"@�K���p�{{t}4��H|��^���ձ��C�QD?r�t���<+Zgb�,�[�A@|���
0�~,�k�$�ԛ�U��2X��?gp�����ki�~�%��u��-�R��^A���2� �BP6ʫy��ֶ���8��Gn�7�^��5����8Y��� ��_��Hr��Lz �����L4�)3��G��u�����
�.v3Y�lR2�]�1��}��'���z�%�B�Q��x?%_�P,��4RǗc��%eև��Y�"�݆��Pfy�(õ�PW�K�A�>T$;�l{��!���d�V��+��[Ծ�&�P-)���mKR�x���-x�"?aJ����#�xe̓���#H.�#������t���(�!�Ϡ@S����"J��q�E��A,,Y��>�c:��c���߯
�qq���d�c�*�y�{UI��G@�(F�@� �&�/J\' Z;��7E��Ǌ�-�-ɒEECm�ᘧ4uk������؁�fZ��|Fׇ>�� ����m��o��FK��e���'i.�\�G���L�Z�Y���N�QQ�$|gw�q'�����s�y�qc�T-X�H�#hy�%�Fxn�4������~�����4�L~<s��G?��*8�m���Yh���O�M�����s�#��lo�/%p����"�1>1ю}_&(Y)И�bX���O<�$���AEJZ�/��d%ɒ�L�`��voE�MEH>�E#H�?!<x��
�,G��E�	/�=찯2F�W� j	K؉��R��ʖ	H�h�.-P�:#Rq	��Q9%�3AP���t.����J�ZvR�,�iO�۶i�Tu�u#~�˵��ֵ�u�k_ǭ# t�k]�Z׺ֵ�u�k/�0��2��� W����A��"���8h�R��y�@W^�XF�W� �2�D�0���
r��2L�Q4��ӛ�g	�k$���gG�nޔL�eE1��`5=��Rw3A��L�NU��~o@�k'���#p^I�z�_@�����"�O��V�xu��WH���j
&�M�������[����؟R����+A0����ɫ��\'	A�� ���!��$��<.�n��P�I$K �ϵ�=g��ܴ���%.�K�R"���=k+��L8ޣ�Ν?O$�#G*���l���e
j�X:x��v*1�
���
�:yN?s���%�d�]'d ���Ē�8W�O'p���f�H6�ڍ�4�5"-��=I}Y��[��7���5��_�2<��C�YW!�ң ��?�:�Ni6��
֊�HYS�Y�Ϝ�� *6�/��{�)<����N�]����p�\�����Q.^��� �dz��.]��ǏH�YcT�[jZ;I8��yB��+�!gi���b�� ϵН����2�9o{��`6����������8r�0���R�ٳg����>}��S�G1�|X�_*X���#��`=��H~J��0V2@P�՞�ξ�{�+6e�f�K�Kfm�=U�`d��>x��\`�bU$�hV�.Ҡ%��2�m��p�J�-�/�"��E�N�������U�U�D&l�K�_������H! 6N
�0�{Y� !X��Q)��\^D�d������y���<���� ��q��ys�s������^(�#�Dv���
жbcU�N��'��
�J���+F"!���?r�H�~K�˰��K�M���BH���0�(v�6�`��`'?��Y�
�٠Ƽ�qD~��{	U�#��\R�p/B?@{p�a�R�k�	s����9�����"Ai2�U�I�$�壈7�r�#�4��=/r�J�`R����:�xO:�eH�뼶��w�^"j�xi1p�����k	������"�+�O���Ck�����^} ��ꙤPy%+(u',�%/U X�?��@I�a@7��x�t��)�G������u	�@��g+� UTg>Z:���H��'��4N3��o`9�g�Q҉�ؒ����ҿ�H!<nD�Hcs��A����O~��/�s�L[,A����V�8w����R_�{�<���s�m�����׽�ϚX�)��%�޹��:dH�L�b^���~���y�K�zQ��N�\�|��"�q%��h>2�M���p��J���ono����t���C"��^����Й	H��� Bq����q.C6����'����)!a���Ɣ|��HT=��(��.!��j���?!ެ��~��z-���YZ��}��>��A�t a�o@�`�p�s6�6\f���PA��1ֱS �Z׺ֵo�� �ֵ�u�k]�Z׺ֵx��T��h�T$��`��Tqp���T0JB=4�,cl^R�\���@���Xb�$�%j���6 D���Qp���ף�(�����(9?�^�`�ϒ�xyQ3����A2l���9�F����ܣX�*%�/]l�p����E�:���f�	lmo����?�q}��@�s�d@�!	�|�OP�TAjV�%�]��vJ��;�05���x���&�?���sgaue��v̮F����AZ!R(8�ȇΩ��[�7K�9�����Fm�|�t6�y]3H�ھ}�����|G����.^� KKK0�#�ާ�Q�aoo
2ap�>�,0�}k�~Y�\k�!͔�	J�`0>H�I�\�|~x�9\簺o=��2Kѧ��n�R���Ϟ�o��EJ�jX��
�kC���s���}D�1+�2&[�N�0F�.��!����Y�a,�p������ny��	�9�$L}l��$�۶��(�D��U�k�鲾9�K=`��y��y�@5(	@�_�Ӄ>DD�kׯ�sO�S�җ�D$��n�>'O��}�#`\�|�~�i�nm=X�^֕i��A��w�+qƀUY��/��
x��7��Y��p�<_SK(��?g����L@�Q/�"
Ī,�*��@H .���}@�<ˌg��(��2�-s�2��D�]�(!�53��.�q�rqT\2&o��J�:^�� ���I@�Q�٧:(�@�L�X0	C��We�	(@N-�s�=e֔��� }��Z����y�
�g�M׿�vK��1�R.��pM#��*KKC�H��#�}&��/�Ե(��\4B�S��$�!8g�!p(�L3�u߼Y�=�Er���-@v�Z�wnD�}PCO�(f��!̼��*�O���;q����M
E�H}y9�f����;9�1Y���
Q� ;ȹ@��r��׉�ôVMM@l�gu�(�-��ґ㓢>s�R�c�O����6�Ǥ|���˝`�y�Q�RԦ��znS0�Ƭ���O/ϲ%+���y[y,�園`�*�����H�t,��S��62a EvzЇɸ���\ӄYZ��t݆T�,�r�+���ۀ�T��H�:��J��+We~���&���v�q�dW.o����|��/�F�P�}|2	3���yގ?����	����N�;��D�h$ T ���Y���D�}VRR\T��2?<�T6`2��t.Z]]�}
��� 74�7�.��X�σj�A�].�mZ9�>ؾNO)j_����V��׋nl��;[�y�y#M9�d[��&Ĉ���u����8Ey~VSb­�Ш�>;Ad5� vT��t}��LRQ��O�����z0Z�t�ֵ�u�k_׭# t�k]�Z׺ֵ�u�k/����
YrP,0�G/�IX�Z��&�8��[��2�S{壏���GI~{}}VV��.8�@�a809�{�M+��`9�E�L��Lؘ�|��l��Yj���ha��pݖ�\|�� ��Zg�0�L�S���\q�yy�2ܱa�r:�����-� �%�����`Ies��ï���p��S���#����~a�fFR�X+��*���%��~!Y�?��߄����@�2�د��XKh[��K &=��q��n��W��2�[Rh(��٪|����F�%XZ�3��#������*Փ}�k�n��65��D����:�Q3���9�@,{X��*��A��`D ���0)�t���d���8�k�3��ns�6\Q��@��5�^ƾ�X�	��x4k�ԍdk�#��Dzm��C$��3��VW��m8th#�o@�I��BL�p��e���h|Lh���3I��<p#�C6�"���b�Dؐ �+�a���U�dϽ�N�9/]�
{��0Z���;�{���xœ�n��{Hk�"Z^WW�\�"�g�E���bB^[��I�����k_��%�g%"�M
�`f"N�ѳ�>�Ї�w��2��7�Gk�����?��d7-<���ݙ��Z����-�w���{�������r�$� u�_f'TT����~J�K�H�'B>ϕ9\ЌM��d�yo��2'-�0�g��� �8�Zoߊ�`�v�T�$��KɃhp&[�����	�>2p�@
P�Dl.QL )-  ��
�j3�Z�t�L��
�@4�.����Z ���`����m��8pL���
��d�B02#�����߬� ��}4�3��-)��F���Y6d�Z�*�������\�AC�K�a
�o.��6S�ލ�8�wH��$c����#
� ����س�<�)�������<T5/`��'D�e�BA��L�*�Bd�]�H�V3e���E���z�Zb(��f�BԹs`�(�m�E�o���������t>����<�b7��X�b�U2_}Mζg{B�Y��G�E�:��c���?2�'�bD�@��TM�!�����\FB��⩊��G����ɾ��m��k������y�� �,Gg<�cE�?h����Ǡ�U/}-�^<
�|2�~�D�����|
�ٜ�b��n.�ϳD~�X�2�T�)=O/��Y:��p��~�=� �5Ҹl��
S^������g�^��~0�8J��y�H���9 �,���[�~��~?���Y��
rv&�\� �d���
��p80��P]K��8��b2�
0��=zT���Cg^P"�+�����'��oeQUL�QU{�f��Ϗ
�5��?��z�)|��a�dx�鬜��Љ�H%�?A�@�7G!��͜m�	�S���$���'�sD+󦾕H��H�H��}� е�u�k�h�# t�k]�Z׺ֵ�u�k/�ֶ"W�3LL�#����$���Ep{�#���>�o~��`߁uW)�X�����r�!j���E&
���l�� ��:�`@LAbт_!h�M�
�Q@S���`	��	\�~8oz�w@=��ca}�^��g?�y���_PP�$�U�@��D���$x�Ϊ�x�}a]�Y=a���ʁb��犞
L�ځ��E�Ç?�"1<���T����XYY���K ���@�]�l>�L������2�� ��@R�(�&��Yf���T��_��W���.z� 4K3��Lf>����T`(�
0r�砡Z�Cuc�|�Х�2,-�p9��Ŭu$&��77�Q��	-�z�,�W�߁<+F�	�BU�'��F���%Y�94��!�U_2�Y�q���*;4�< ׯ^������8H�!��zFkI��yEzn]Y����$������v�����
�@j��X]�p)���lom���:ll쓀�������<��v��PuˁPy
��+8ʫ��s��M��H}���UX^Y�յU����#��F8�K�!����=��Ǐ��~������ =ʗ_�x~����677i��x��p�=���>���G���42N<��K�lNa>��I~�;�5�E� P���xWB^_�����`����A%�5K6���tI�K n�O�*(X��U�p�R
Z�O�D-��fPf��2���5�^	xZ�,V���֑	Y��x��3�Q`Z�� &�o�b� f�nc�<$���+�@�'.��3�`,d�l%e�+�l�!7�r-��_/,\@�/� ��J	j�o<���|Q��d<R�����9���ҡ�O�6���TȶR�Oq�(�Bc�5s"Q �5i��F��;gcfjYC�c�Y]�)��cJV���_5^z�s.����~�P*���/��Q}d^��WA�L��\ιؕ�y�x�Y� �����­�J{�gC��}�����Z9o9�/��5�� sY}Z̙��Ca�F$�%0�����i2��%��^�ZQ��{������fI���^�S�+�m@UqD�X`�5�W���{�'�Ɔ��SRfp�3�02�������������2�E����=��3
��3\��#
��l��JL9����ᡇ�W���L'dǴ��O���z._�׮�H�vM�8�]���N�>ecVQm{&a�2��gm�VWW��Ό!���������cD��Mә1��탹̇��
�9�̒�H%�-���5暹�=���:[��\�A|8�e���29��=5j���Qdz��y|���nb�&F�lc�)�P��&�~H�H�\דrD쏂�FUʬ,����ۑ*iDd}��/�������T����0�1$9-Ȕێ-�j,�m�ۮ��׋��k]�Z׺���:@׺ֵ�u�k]�Z׺��l5�1�IaĨ�Ѥ�KI�R^�C���ȗ�8|3�V7֠7�àߧ@"��;��A\�l�D��\��w�� an*�%c5J�L���	(jVlo\���<�a	�Y*���j���_�N��]ۤ� ���$�1 ��v�v	Pl*VP8J0�C
�2A�y����z{�ɬ�����6�� 
bD�b�T�t�g+�Kp����M��m/�ӧ%�:_�8����0�<�;v<B��gN=�/^#iж�l|�VÒl+�a�g� �V��ʓO�����{�KyG���F	�b�	4#�r��gQ�g���`���&g��F�Q����V$�j2�D�Ҽ�mG���l�7����g��eTl@�AS�~-Ae�,H�=�kU7����ڷ�f�yC61���X���7���>�=�����~F˫p��U�P����s���@=o)㴟����lLA���F�+"� �����0�����P�ר��$%_��K�j8��F[��L������|Ҧ瘦�L���-� ��O3�e%f��z�x�+�K�zJ@3����2������1����5g�1��������o�k�-�}-:tX\��$`�q,���r������~���c��k^����c��}�{x)��N�y��.���R�8+��
4�ZA�Mo~M2�fI��5�J'�_���d �}Z���3�^����Hu�	���d��|��.�.��0��>eI*�0(A�I6n0��![')pU,���K��2t�y��%������'��$f��3��� ��N]z� �7� *��\��n���\H�3,�����U���E������\�-@Id��1�`���NQ�=L���Ce9o�����f���$)��	�+����u�`�����G��J��?RYIs�4�����.�=HFCG�d���хz:��',�*'*+�L�r0��x�}H����3k�ܞ$;��&_>keN� ~$������*�(��O�Di��W�	|�*3��J��b�vU'_�� @?��^��%K^��@r;pd|I��e��lQו�=UfDAt=ߘ-9���M��av��T�`p^֌^�87a��_!ٰ�s�0+[އ�P�Q�Ǿל-�b�V�#��Pf�H]v]���27�4�;�M�����!��(l����(%������7�t]��B�W!H�{�35�d뵺p�9?�kٯ�����'>��e��tn,���>�1�����^l�#xF�E�����o�v�����̱�7&bjU�0L{���
l���}���}K~Ѿ��F�S?��߁�柑4�~��Ȉ �O~~�w?Fg������S���ͯ{-|���	!0���^�!��%�~��D���x2��0���U���/c�gp%�dk�qh��l��TN��D.B�>c�e�o�})�	}���X
+U�Ot|�$0���1=_E^ۤF{��!����D�SV0	�U٧}��Bg�*�"ٷx�Ȫe\5�I�m�3�+^+$�P�9�
��y����Ƥ+�RJ��J�:=O5�%�Nӷ�P�������k]�Z׺��:@׺ֵ�u�k]�Z׺��l(��9�$`7�:CtUPY�X�j-[B���5z�ߣl�^5$^�U�?�5hM`���;�*�(�c�xS���+#g�k�YgY\h�L� �^ Z�Q��u�)3+)P�>a6�.�:s��w�2AAJDD<fJ���,��I	 �kvG��"��}%�$�:�S�v������s�����$��3+��,x�%�p����׃������sg)Seb���awgF�:r��	3�.\8O��'�|T֗k��9�.Ud;�n<#{��1��F���0�����T=��ƌ8�+/�T��@��'��HC�e:h)�|�>��M���M��`,���p���3e���cf=��~�ϡ����h�ҵ����x�����%;���dK����g6�3�	4�޼�A����?���þ}��4$9�s�>K���O��?@�3��?�޳
�|᳠}��Km6���k�����(�%�|��O�sgz�*�Ô����F�i�vj �C��ԩS���;�;�����d��zGu���5����4�[p������+v��M�@ �2xMR���p8�w��g���nM?�a4�s0����W�޽(Qp%f�թo���Zml���+��o~-��}|��O�<!0	%�>�,��@����DA-O�D����{VU����>J��`ଂm*�`�&�dE�(��_��|�~n&m9�^�DU��*�C8Z��eP�d���D�� ��r�i͠T������E�]���}v�I�o�ҏ@��ɘj-��(�_w�!#h:�>����`D�7���i�����L⌞�ş��Kl��WA���֌���4% ��LR�S�Zk����T�eF�2����&���R"�����p@�@,]R�G�}+�+��D(W!a��|k9���ex��/����,ˈ���^L�ģ�:1�7Dp�!=�����}����}��g���dO�N�O崮v�ﲜ�M�52y�0=*=I����_Q<eD��R�7�F{��bF��3r��i��}[�_�2�ݢ���z��Ԗ\�W�z� ��7��2έH����bM�2�ki_�-���}���a��: ���@�[}�7�u�H�E��RQ@Ʋ|}E�7%θb9ߤ�Q�I=o>0����;�k�*�@3�x�!��q:�����?O.��3��z��@K��JF>Ǻ�O����3�o� ����UPi}$���9��^�m�}T�&��=��������G�4�S��L�Yᣏ=�n܀��?���^�⇈$�c?�~��p���|AfE*�$�B �`�(*��$0�����-�;�2���� z/�'���J	2�Q�5�G�_x��ͩH�)+d�y�P(����P]ɴL�b�Qn�_:�3z��/ό�S�x�g�k�겖Q�!�I'�_���x���'���Ǹ\��D�*���'��-%0!�+�#�x�l� ]�Z׺���:@׺ֵ�u�k]�Z׺�k.5���9��g`^�r{P!S��h�ːXf!��D$)m��)p�A/�a�3`�B!jV��ks�-MA ���eA����%�т�1HR-�������:���"rF>��������gI�"��@��$���j��H1�	 T{آ}Eƾ�	Qn����(����Ù�:47!�ypN�-��U�G�R�eq�*�x��������/{�K����*;��ƀ#f�?��YrH�E)ӭ�=x�_��欞ҵ0��5h
d�����@��D�&��б#���γ�l����h��R�50��>�}��0ƍd��l��Ϩ< O$E]c��Q���`��y8s��M\Ć��˗/�7BH �����e��X�����s������ac���^�v�2�0�?{5݃�ԓ�>pAj�"HY���4���6�3��.�*�3�.}�&�)T=A�/R�bm}��~X^�h4�Rۻ���5�,���~կ���%/����8���B��>u:]��w�E��O|�	��?�4>tn\�Zy:D�#������(��8Џ$	�$@�}�]D"�c�*��{x�)8� �t^����w5C�GFK#XMπ������0�$]����i=�H�ڵ�D�	�%�ӵ����[P!V�.��h�zH�����4f����,}��\���g���~H�8
�;�)�<���,W�Q�}�3�s��b��^��Z#�B�Қ?Ѻ�J���N1S.kR<!=�����-3&n�����G���h��D�`g�f�-`�ȏ�*��X�Z^'
�0 ���Z��2�N��w�l6�!h�����,phHu!,��|f�}W�6�<J����r�@��*}ϙ�B��r#x(�� �>\G�~�	]d�L��� %-<��} ����k��[֒_{�ٳ��5�Υ=fUf�O{����.���[����o�C����N�~^���I�?��jv7ޗ�G�4K>�H��"u�yφؚ-+!��O�&\��=����t`���9ϋb�J�ٞ�|�Y�L�˶�`��E�cq���a�l�'��<�!���hu�t�KG��L*/}%�P�v����^8��9݋���њ�Z�!�g����k������v�T�"�4�<n����F��}C�w��%2���*0��X}qa���d��r�����lʠd	��.�@#�|>+=54���:��Ȳ�j�E�ӳ,��#p�g=���/�S_9����9oey9�}ô�Ë����<q9v�{��.�EP���E$�a9�Z�)�\gϞ��W/�rе����y<p�I:k��-��:���x/�?�<�������m{�����a�=��`��V��Dk�##]H)�:{��3ucR ׯoEAKtufs1� ��t�{OK�~�}�������d� }t2��Ӱ=��ȒQYك���'«{=&6-��p���u�XU���!zHd���Q$1%��U��%⟐�!HI#����R�y�"+Y��ۖ����i��2-�Eo�l�?���{>H1�,���]�Z��J�# t�k]�Z׺ֵ�u�k/����3gθ�i0ncȒʲj`��%����T�����L@�Y.��/g�i�i���|�l(�����.{���D�j��2�
�R�� ��$H+�079~v��`kk��������5e��u��1)hF:ʺb�tΪ�}5�G�d��nO�q�,�j(+�T�蔠�&���3^�����x��%Y��}yy�䚇K#x�+_I�Aw��|�	�FK�p⮻�F�w2�Q �\G�j�cD��20�@UȲ�*��A�(Ү��x�"���>|� M�]"NB�\�@�̶@�q���e��G�����$g��IXsvyi�����ղ�Z���]`�
��p��y&y~|O�j���!��*X�$pz�mw��C-��u'I�r]^�VG0U@� �	h��9�x��a�WQ�����Ц����\�G���m���d�:�>`��9q����D��i���/:�)��&����רڐ�o��`em�VV����o� I�cy��;;��F%p��,�Ϯ5�?�� ;j,{��;�o'�\`�}Re EQI$�0�L��R�?p׍ ��ޥ.����*<�Ѓpۭ�K�'��g�PI*A���C���@BHpxi4���kb���|J�Ue
�jL�}��U��[���ҥK0.��т�[�g�)�Z�'�+SpV���xQ��F� bAӟ&V_�M�  �`�f�:��R%	��um��h8[	��f\��Md�(?�/7g�G���ګ�vU��(������[��e�2@�FQ��2��B���ũ��M�m>� L!����v:���s��^˿��=B�h�F(@r���4�^g�޼�� �l�d��xVZ��\�K�ˤ�q�w�wޙ��'����p�ɓp��p��6���w����o~s���nt�ʍ�=��� -�G�!uHΙM簶o� ��	YKp�
q/k�4t?0�U��AJ�6��Q�辪�:�g��B��=�H?%�tO�F�d��X�������,
�����p1.�Τ��g������6B�~�+U���lL�%���8� ��K�ʩ/C��x�Q��5g>�y&(� �R� ��X~��1�s��J9/77��	��r��G�k7�W�6���������J|�QB�F��V�Y��G�{$��/R�_xN�' �
}U�I�۞��nl���W�Y��?ׯ��h:.Ñ#��%/}	����-��p|Dj�<��(�4#K��}.�?O�m,-�6p��Ӵ�Kg,|ߣ�z%��o���)���7 �?H+��������H�S�5?��V7��bB&@�eUڧ�̏����J��4�(~!(i�o6jz��5[�>��Z�-�6�(�Q|��R!�������o�}�ϭ��|��CY�{!��[�5��o�(����\z�Y��Q�t拮�1r���Z�s�����,�B�T�J�#"q�QŷI����.��m	 ��?��/򳴧�3gz������5�nji�׼��;�Y�� �qΝ��n;�;}��{����t��>���е�u��:@׺ֵ�u�k]�Z׺�k��G���e�B��,�Z�_pg��B�Hi������H.���5OA��$}��W�y>�	l�����:���D 7���ke��L6���1��E�@��r6g�Q��l�F��s�d�Ħl��P�j\+����@f�k�ZZw]
 �T� ���.=�� ��������sO����i�j��IP���En\j5kV�,},�<�)�?����#�C?��p��a
�V�e��R/YIQ�_q��91 �2��N=m���f��`M�s"�#>,��<w�l���#�����`x+@Khx~8��R�m��NcF��%Ц����G��e�ط+kw�� �o?]���8+��3��ᩯ<M��w�W��`{{3�_V� Ic�Af�$���3(�������%RO@��f���@T�V�@	m|��2̙PO�c�9}
Z�򫔍�~��2ve�!�I_�S�[-Fb}�f�o\�^�e�>s*]n��(�+��W�^��'�"[����7`)=f���ܪE�����)����gv�XOI
��?y"Ș�r�,��6h�sgٰF �����"L �]%�\��i��A��Ν;>p�7�u^����~�w�8�<1Zk�Ή;O�hy�A���d����(��{����FKd�H�gE@3�?H��g4�8���o���~�W���_���g�5m�v�}��d;���e�QK�DQ��h���\���Z% 
�ESհ�t��ی��-*���z�� ����
w�2�-UY�4 ˫�mxX��Z�\�$�%�1M.��#��E��8�T���C�ڠ�hiCe
��]�)QR��Jm�0�P��:�Y����fG�O�]�䈇z�;F�_}�)���$�i�J0��l�8�W�Y��KK���im���l���?~4������z���|	��p�'i���p0���X]Ik+���?�x�_{�)���Ӿu�\<Gd�umv�*QP��3� ہ��m^�\�yx&���������h.�e���
�۬ڡȦ؀�b)�2:
��/ �ljs
�3#E�5��X\�jQ%E�{�\ x>��DD��w�^>���y���ф�=�� ���uj����8��-��0�������%3�ݼ����X����5lċ�_P,Ȇ\�H�����7R>�D���N���]�\g��"H�S�*h����bÊK��(�,��Դ&"�c�(�u�<�ʗ�z��v���<�Ί��>�gATnB���!���������7SgV�:���;��+rvL�u$��g���ޮ�_l��2�c쏨�Og[�����>�QuV�/����fQ����RH�2%�E���3�t��HO!��������H�&T�K��㝨m d�naI�����KWt��LG�?%����xz`
J���0i�	� ��܉{�~�mڅ릿��},��wu�8�q~`/V+�Ξ�z����M9 ��������Ͻ3g���#螾{�L����=?ad����7��~n�M�{U��][�[��|�=��B��i�Um�W!8���>�E���:�:-�d�>�M4���������K�����o������CZ���|��t�ڧ�u�s�~KI#��n���s×�����N�	d�rC׺ֵ�x� ]�Z׺ֵ�u�k_��(O�к?4����O�W�-F:�D�]�P	@��1�ٶ*�2���� �w�i��c0	3���X�eaT�/�'?�)��ރ���(A,G?O(ș?��ka�v%��d��j��CK��$M_1�H���i$��͜�X�c0����8�)2`) |,�%IL̢I�}�O��}��r��Y�#f:a�7Hil4�"'�7�gQy�Y$��uA0:5�X�(t9�8�r�c������+�kD`��CД����QH
.2 �����s�Z��y� ��Z���J�^ ]�2fy"p���M��'�*���{,�v�_����A��$P�h��`0��qoL��[�[p��A������cE���ǝ]�onn�իW��m�xo��L'cz^%l�Mo�t�UpR	6�+��u�� Ê�V��1Zf0�#��dm�s�h��В�-��\w�t���{֗&r���hK��&��PF�	�G��C����,1�n�����p��Ux������D"A��[�'�TFa{���4=��K��V����U���sϐ2E����9f���B �5�kJI;��*,#"��6Ls��x&�0	�Af��h8�X���[��:Hv�>3�Z�N��i�f>R��Pؿo}��
��7�����{��Ў��ħ��qx��)��W" ��c��P�����r��� ��\�����h�w_�_�	JJbY��) aД��y��	��������,C���X��k���xP9w!�E�s�ُq�_�������	��*2����3�^[�;��V������֧��~	(�8�o0�Y�\!-��unUe/�:�7#�Q|����l`�Y�r��!o��~��N����c�J͵+��rZ�"pׅv�x ��c蠗>;a��0-�:L������������76a4X����d�}�U�T�YT��E�����>|o����=`2㵲��M�T�>g���t��:��UQ5�����@2?���:��"��M�C�CE�Tס��������l+��I��_xUq|�)� �V2 ��)�L�c�N,����x?w�en~�2�`G2��7�P���+���Aj�G���k���J�P<��쉱<�@	ǋ/��٥�K���n���ub�4'�5~o}u.�t�ԈwNO,|"����ج����bV����b��\�F�\��@P���#p#�A��;��Ig�a5��xvC�����X�'���0�oeu����t[Χ\���������x�'߲F�z�G��s�=r��<�W�j'Og�1K��kDt|�����.$./��,��f��f$ݱrK.��=�/��',ۈ)��q��_����&�cU�}J��)IVQXv^&��|>��R�<���~��y>�G��E�O��p�J��H�#��֙� ��uttn$�n���!���ma��x�'��jj����T?XF�*?�wv���87;0��_�>�!�����2޵��1��=��mzw����ݹ]��]�E�l̍'���a���7M�J���&���ޛ�ږ\�a�j�3��ݯ�nv�l��$*�$���(�"��H�Id$�� �� ?��IH���� A�4D�(��(��q�l���&�ӛ�}�;�{�ٻ*���VU��)��.�����=ԮaU��}�[q۴o��Ǩ�g���ǎ�i/=�ٴ�ϧi/<��+��<�=����8�'��g�~>ͺY���(�U���m��lb�h�}��IM�h�4���a`�s'��I��]/$�8�_��
��Ќ��5�}D�(��ic;jB��^�tn����&����=�<C�P��]�� 0��e(C�P��,�<��Ui�_�ތF#&�K
C}�N����i�񞥗ܸX,�c�=4B@�������k�u��s�qn3v�]�,�T�
q貳���h��7w9�g��YUJ�r�>;�ّ�:���y��ho� }��g��>����z��4_q�yt���$�ͽ��
���Y�˃<���t7��F�rNG�p`�fL�� #K�)����F�`,�x�0c	}~�0><:��������<���yw�j$����ڝ�Rw3�� ?(H��"2���=�GS9�C�PA�X׆��YAyn��t�������8u�8�@O��4`Q NOsv,s{�6>���/9%�>��`�������>�		�eG���������\�M���#�;�`w��ETU��a��������О�*U��f����9���b;�0^��D�z7���}���m?������s_J�6t��Kk��� ��s�F�1ф�����h|i!? �-9H�C�\vLg�k� ��[/@	�%��9CA��đ�,;����	��!U�U��q�X�2V;��s'QL�z��� ��K�O�W���}w�>��O��O<��|�I���Ϧv����!��� ���n��O��)���R����8��0 ���%���s��i�z�s�s�r,"�ֆRa(	�gERR�yͣ�� \�v����.�9I�A ���A�`�	���IgϞ������i2�f ���}�K�����J{�{��SO�J����6Oc�Ͼ�^z���;c5�0�![��'���<�K�"��R@ZA�`ഓ�G�oi�$��ۃ�"�ȐYl9�Iv�φ��E�D҇P��),���w!i.�Fs�Î��L�sJg��3��ǀ���j��3���ކ�V����E#	��m�㆐���48�J1��i�I�'(�dl�Ȳ�m�~-𥁌��3a|�����[P�y�%ڸ����j���:ڛ�zc��2��`��M>����+L���OsjJ�>������������_�.|�~� ��}�S�_�I���_�O���\����=�&q_p�&���d����	��	_��.�:�OV �ͅ���l�d>K�!�,r�XS�!��p&#_Q&�Y��*�0��j��%ѷq�Q�m=^����ݐ�%�9߶q���
 
��rJ��Է���9r=.�;��r���8��P����u�״��;!�0A!��RK��U��`|R���T>Y����}e��>7ޮ`�WY��zF���R��$��וS�Z�ے]��y@W#M�"�� ��d�Hz�!��9!� �S���$�sW/_��f^U��)�����=�����&�1�J�x�5�JFG����(�� }�6��큓��^�lK����19pk�6}���������}��a���/鐉�A�n����E殨��^��o��	��̲���6�H�����M�5�m�!L��u��se�����sȐ՟�7��,�sK}��7��0)�����2�
�ܠ��Y��S�)Xj2�b�m�VV���x4��Pی��L����&+� �Pڇp�~�a�$�!�b������d��=5�'Rw�Mz/bu �6󦞠v�hi����H�����k7��e��x����i��3%�վ�>�'�>H�9Ǟ#
�,x{��X|e���c��TgV���n����}7��]����=�
iޤ����g/��;ױ`�]iW����w]@� ޖ�!ɺ����5����"�y��t���a�i<�`g8�"1�i��i[�t5޲��=JO�ɽڞ's���l��M��``�3�>rԿЙ���5.��������~���s��8�MǤ���zd�O\�:$H���K������4��0� z5����s(C�P��2 �2��e(C�P�`�_>���/6�=�����x�^���0��I����_-��y:v�ކ&��ē��tʀ�8�m���ڟk'�l�ҭ���.]�<tб�n� !a��.��P�Sɮ���onn�|������E�8��Z�F��N
l�q�#�����X��D
z�_)`)�+9�97 *>��g�>�I�r��o����cv�A*��S�9���Jϳ�o2]KwZ��(x`�����;"�/R�^ABxl�	�[$���*�ʟO&��x�Ə��PvZ28Ź4Y��ٷ}��Fi'��i~H�a2���Y�Mp�E�G��C0]2j(�ID�}/�Y�Z�e�gg�@����\�O|�����}�uH���P��]������s�^������x2���h��.��W�� j+�<�φ6Ϟ���9�e���qz�&���\��x�������dF��1��l���B�������l�v��Йt���Te)H!�1����`2����ޏ�x��sݾs��t:��$nY4r��"�9E'i(�H �w����!�z�)͞�V��l����l�lpD�;�l��=��LV�t0? E��O��ӽS[5'�ى���2倣�#���g�m��8��9������t&�������mz�{Q��=�5(L�x��#�o���cg;y��z*O<�����ãH��'Q]�L&�=��Sŏ�ã�p
8d\�%���kV8`p8���K,�x����������ܦ�΁���њ^U'\��dg�s&�px����+�FRe���pm����DEd��[��ʜTyu���9b u��,&�D�KZ�Z�d�M��)x%�

��2�e�A��L�����qeoy��)K�\���<����wb_r$$	0�� � Vnq~�6^�|o�8b_�?̰ex��$��G�f��B�(�Um��g�l4*�'�=��u�Wx�I��>�KQ�]X]���-�_#
h���>j�`3RYa��`�����h���p��J&_(ѬܕQ���WV�`�F�u�ٽF��?�t顇)�h<������q��(�������O�4=��7���v����-oNsB�Nލ���9z��oIk�c���twg�^y��#�w�M��^��������8�1�k+�R^������\>�]�����5����x�l"v�U �������K��#�%��gPH	���ThBE�U���5��Z�އ�6��px\�B�<�bt�\�����%+G�s�BX1�B��2������h"�!B��iԿաRA;���ݗb�3)��M]]�˭so�J_�~	W���T��S�\�%��=/"5� ۈ(�_V5l�1�a6����i��45GT`�_�z�����W������������L�{�檼�N1��U��g���3�<�� 1�����H-�}3O�b0Z��&[�R��LV�ؿ��Ŀ�t��Yؑ'�|�>����;��,�>jǰ�ث��ui?�j�y^7� x�%V���t���}̓\�������ނB����S*�0B�ѵ��˺edi`b�*��}��xR�"��Nh|>���9�d>+��������76�imm5ٴt�����
��l�����OV��~�/����+�|y%���aԈ�X�l�q�O1Q�S�a=涜uF�*�aPb��e�cT8�J�@ڶ�N�ྎ��������q�ᑴ�yW:� ��QM����u�R�=3x4�݌M�R%8�#��y��b��_ ؟���,��{`��N�\���=�*���:q�Q�(�,t3���I��� �N�D._I��[y>sUI��~'
��1q��>]����� +T���v)����a*ݯs�?o�Z����E��>��r(R�i��^O]z/J�%mw׷��� ���Fꆡe(�?-`(C�P�2���T����/n���<z�ڵw���y��;�]׭t]h��i��ę���^4C)�N"��[ا|�MpM�7������W�?���|!��z�w7�u��H 
���ׯO�}�g��z�4��|�	a�o������%+��ؘO.��s�|oQw�Uf/2ܐ����+�f�p������yI�fɞ7�1_�)�i��U��]��̡�4��R��X?%+/�!x.�>,677��e�X�����۽�g'�)",���� v��Y�N(����ͣ�����j���[t���$d�M�mn��. �
 56���G>G� �7����$�=|�B���z���&��F0�';%�dgG��hHvJ�(�b����v��G.�c�!��!��sfšU�5R�WTڛ���Ý�֭[��g�8�SΜ�M���k�%p�"y!���F ���w �̎% ćD��U���5u�Nƨ��V�1��$���M�� ��O� ����;[4]Y�յu�N%Z����G�"ĭ۷���$�icmJ/\H6f��1;el6���~���Ϡ�67�qݳg���ۨx{�� �W�]C�N F����]��1����#���^�#u��[;d�}��$ �l8Uy,�>S]Cꇓ0C���@����h?��
�r���x�s,�
4��h����9�{��tA���͠0���I_��M�ɳ�6c�^��d��i�OQ���ulK:�3�瑲c1�0o�IO��m��d��ݻ�p���N_�k�#EH%�~��z��aL��$���/NhD�A�=����Aƭ��1��mЂs?�裢ʐ��d�D/
)i$~�����A����P��ʑ���UB�Զ�%_Q�p�M�B%��}��R� �A�3%
-��H�#.��m.�e�>�( �w9���
RS�~�|��NH>���=he^���`�C!Q�),�u��8ƶ4�N$�M� 2�\'��6��SpZ�"�ljܸ�7'<��)��DG��`�U��[!pb��łf2VNts
X��^5n�h"�|�|US���3ذ�D����6R��}4� �����������D!X i-���+�gΜMv�"�=4؎��N��E��R�z$��1ݼu�V&kt��t����k|����Q��vd2�3<��k�E!�8���ܹ۸�{�m:�޿��M�gRO��6�NZ��4K}n��u��d�+��K����+��ǉ����^�e��+��Y�/�r_��j�.֖��4X\U�拍�� c��Jv  ��IDAT��{���h!U�=���}`����ԯ$�m�c�)+� �N���1�����Zn�N�#���՘�"ﳍ�Z�i%��u�nS�a��~Z~�B���w��c�ĺ��.����V�kK�A�"-��b��]Qa�4 �$I��ɽm�f����R9�ܼy���������Q�/��_�E�'��
�����^�m=��|�w~�;����/���'Hc�i �k3�Cۘ�
W����]����]���������~/}����c<��c���y��`H���3דI���C�rL�^��>]kAoy�[Ȕ<X��� �9`B��59���ൡ��h��v�P@��]'!�%����bӖ$�RhT�MY`:�A����M
iO3�h�k��xg�6X]Y�M�td^zI�"�A����G��7�Q��ʪ�� )��kL��:�_Q�V܇B*Q�I�}�1(��B�sʀ�X�!�iD��������'� g���\�����^d���P 04�}�)��M� �]��E����m �su,�y�P�ҿ�7���5���x��k���[��eo�i�L�I	�7��JH¤i�B��ZR%���PV	A��&(�{������N�v���e<;������|�oJMp�4)����},�P�2��|�2 �2��e(C�P�@ekkk|ew���/���;[[���}<�]L/����q�a ٱ�E@��_�c����A��M�C��}:�d<���x���?��#�����ڌ�j~w��KX3�?��Ϝy�ƝK��ѥ��ك��g;V\t�t,� �8��*ԃ��@q~�8%�Y1��yɎ!;�4&@�ر /����%Z<��G%���4��}q���?-M�+
�
t4��=����N��i�č%�K0�P���`"�r�t�<=�I��I����|����v���R_>5O6�v�;����\��H����*R��;D�4@S���r ]��Q�:�z����m���/�}9xe�D@G����^b6�9�$�:*�/��Q��:O4OqP =�\�����s������ώR�-����:؝ѭ�R���/�8T��1I���oK�l�3o}�Ν�H��/�FO*@�/�O�}�����E�	�p~{�^|�+���)�ϡ��	'�`z�#x�\�Q�aw�
4��9��6��L ̌@��8�m����K �8�ŧ� ���8�\���ކD�z�5�����i\��15P�QQ�z��C<��<9>���]~�5Z@^�'�W�n���-D��\���[��4������'�z�;�E>� ]�z�nߺKG' ��9�uvBC�!�c��ɟޤO����l����F��H�B��S�$2�����=�o�a9U�B]:?��n7üa'�h2�@[+ ���՝�/��������uBӑ�[tE���9Z]݀�#�ډD��p�.R���7^��������'������_�#��)|2���'Uy���^"m1%Zi�Q}�������@+�B��_y�~���U���767���+�����NI"K��;^8�-��{����A�3��2�� �&9�	ˍ����_}��������W^�����襗^�����Z��\_���h|��W��� ����;  r��HрHH���c�q�^�2�#�8��{ccu���	qG p�1B�i38)�U��>d�~�A�g��IK�"��e���d�"��+���^`���覫rW`���@R��J��(
^�Iv|��&&6$*��@Y�O�𝓔��@��Hf��,��8��6�_�5!Sr�sTҔF{kx����b�tfޢ�c1�4�ٖ�� �>s%�����Z{��tg�&�d���ڮ��#���@��g�Ѹ �"mY̓�!�4H��osf����f^O��ez≧�6���1���v��/͓͍U�����d���_G{���З��U:sf�v����}�����^{��y�3��:(x|4�����4;L����ig�6�%�t����༩\4$]g�u���5��P0%j8�Q1R�����g��"ky��l�A�2�e�g��h�e�c�ރ&b�.���%׸ikv�.�<�ȕ���J������
.O/˷��פ��@-1.%�E�dB)�c�ymW}�f	U?�U�U+���9�R1?K��9U�X��U���"�Ň�v�s�앬��
�+B-��a&v�g��Iu@���3N��<����B���V^B�� :����o��ʯ�Od$�������ݿK������8��.�5���A���?��q ��~����L�a5�ɤ��ms
��_B�������?����K�<D�������_h=� �<f"%�P����0�����؏���{��}4��N��� ���Bo�M����s����K_��}��i��&�y�Ԓi�#�=��D�>#�FT�AT����N@E��qT�A;؉�N7wt�	����e"�ͭ-�����.� �����4����&�y���k���48�{��^t�����{�V�J����*���R"x!xyWr���=K���e�Y����z��Z����.h&��i%�![�b�Svڹ/�q��?	{@�I|FF�������^�&�������^	��N��}o ���L0A�,��H��H#&z�Al{�rT��'j-�WB:_����TE�:!���
�Im�<��r
�녎�X���IB
��cϦJw��+�8m����T!��s�F��p%�EC�P��]�� 0��e(C�P��)nߺuk��_|�k���żb��}\M/�#��9 ��S �W�z�Й��������F��֍ڦI/�O]�~���/���n�q���t��n�oR�}~{�X,.���7]�s��;��|pt�H��Fz�_�ޥ[ �E �|�Пf|P7��`�h~ˈ|���n������
҅�IN�����NoTס8���Ke'
�~v�p�(d�S5<$�ũ�x��u�sXt0@}f+X^N��������/�����k|�D�"-��'ݢ�8>9yp��v���hmmա7S�\�v��\�yQE
:jT�q��i5A��P��}A�C�Q~.fys~&�gG�g�De��x�|��36���sG��+�9���ap�� ͥ��s� ���7�;�k5�"���5�c��������W_}������~�����ЫCUz},s�����BT;�R����E�T���`q�� 	9:/X��"'�#U��T���&@9A"��;N1;��^���*%�x����,����3�L��g����X��Gk��wM��#jnoߥ���52�s��m~L'G���u�ED�[��Ϟ9K^�$�#��Z[[�@� ';�G�Οߤ3�k ����D�>����D���H��Gu(���W�#��ЋT�S�3@?��P����4�s�NX��}襯�X�^sZ
���4�-���k%� ڋ���)��K���ٳt���ݼs���g��ߥ��8�8#����y7�K�
#������I�!�X�4�U���4l�c�����}���v8>:�H%����_��>�"�h+�kń��t�U���EW�^��$�a;���u�LG�:D�3	�#M�����,uA"D�z߸y���ޡ����B1��HBB���5��=�2ܗz�ډ����|��Fx��z���V�d��eŊ�]а�<�d����q[�2�38��C�~���N�
�j�u�f�O�=���00�)Pc׵�2h�M��v��<N���}]�M@X[{����'#��;�c�!9���T���9ãzL,_J�t,���)H�8a�_�E����J[�ҽE�9o5Lbݞ� �@� .%%DTI�p�uc�����^S�)��r=�J���d��� UxQ�p�=��ء4'fi�����ᕫ��O}ġ��������I�m�g�_���.��<GO��t���o���u�!�+����j:wJ��\��P'�Q��f@����>��衠"�?!7�W�e)(d�`�gy�k;g�E�LUK9��z'���2�V�_6��c���:'V�?�mG�nd�D��3�|��l��!d���|�����±�a܇eǡ�� ��a���9�SZ��R+Tc����������Υ�Ӳ�e������?* �}�ɮ#&����4%*m�*�X�z��y4n��Q��,V��Y�"��K/�'?�iz��x��ϩ/~�?E�x�;���0]�|`�8�w}�Q��?@O?�T�Z�����'�~${a��ں}�V�ְ��Z`�F������������~���7�~�?"�Hg�0�-���BAs�Y�=�����G��7=���t��5��:w�\ڧ����s��o�-� �fZ"�����5����d֣Ne��XM�`��c��ǒ��T��<vI����>(c���5L��A�d11����{��g����6�Ux-�}�J�_2���IF�ڪ`k���µ�Whww7���Ǽ��Y4�^���8� ���1��7���X�(-�����v�@�����I��t�/��e��}Em���NՌ� b�� ��:]'��<M�c� ��J� Q�C�8Yϑ��Q��5^_ZXa!�*������q*9��,C]���-�����"�f6^�x?�HT^S�ȃ�Y̏�1����A�bS�eNW����F�~Q�~�������^�y���hD��x_�6��e(߮��e(C�P�2�7@ш{��vtp�����[f��һ�E~�N/�N�q� Oz���S ��F�t$����mӴm;���Vf'��_~�Vy����g�F���x�ܽ{��O7af:������p��M��̧�^��t��/�Gc#�[(���U>�Tj�ʥ0�b���}���3؋��Ֆ ��eG��)W-�Q��\�uo��ՙh�8�,��'9�u b�W�3ҾF,�����Ez�V��:C!-��QOsv�G�fX]]���v���!��.�N �L�9����8ZЕ˯��s�i1�!��h�9��F��Q�$�Iuu�k�Qs���� Wז��SΔbv�zK�9������i�xV:��{�!u Gt��9�썦p6Ҽ�Ӎ7���p��l2�=�ŉ�+�Ƞ���.ڀkȀ�/� D��A�0O����&�:����9�!N���J��G企&E�Z�A��5�6�� �<䭿+�^oc����xs��U��k�y9b��4,a9K�\���pW�O�D1I���š�O�i�d������W����.^8Gѹ��2;��~+��t� ��4�vӘ?wfS�zQX��?E��D<Xox�<F�X��B�2�Z����Ur�����mZ_S҉IwF����&L�����R�]��s:�;��{���У�����(ى݃C���� >+��#�AL�$纀�"U�`�4 l�{�3�IJLJ�t*iJ�4bW J�	Om�!R�����cD�S�Df�c�Dj��V&c��Yն�-��ǯ����_�o��w2�te��t�^�s��ʜK�-o~�>�g�R�����'ҸX����2��#8��h������?F]8",�X����<��m����L@a�u���H Q�e�����M2��╩_@] +�pRI!�����E&�����~*�h��9�Mu�@���ϑ�ߩT�*$���%�1���d{&�& ��'�uh�˦OPpO�t
�����0��k���� �X;��W��� �r���ٳ,��:~*�:]�n���C���i�H��GXJ��O���sp�&XCY����l��"GՋ�6�Lm���<?�oi���EG'�ɮM�'l���\�J�bN���6Z�'ۄ�7�k�v��ˍ�v������7�kQ%J6Z �f+�!�y����ڂI��o��������7�2��m�}|,��j�5���}G�}F���Vx��P��|�nV�c�5۞=)mZ�Aru�P���zbi�5��"-%�pb�1�]��3Xhv�Qua���/y���n����H�e���Q�$�V�i�l\e���q��{����v�S��̀=9S�Ym��`�<���Tr?�<k�� [単��o�Ư�{��.Z��K:��ٓO=A����4G�m�����n��k�׾�U����8�y�jP��~��ң���{/���ܧ�{=~��}�ߢ���~�>�����&�>|@�������q��C�����A�[�GI�M��[m)a��Z:��H4u��������/�1����>���=�����4�3C�ߺ'�j!.C��,�5��UkLy'��0|�NS�@�,�AD*��?��,�|�E��-hg�.�ܺI�ǒ��U�B�I�y�ml���鞁t[\�;'�a!��"Q��{�2R�J�� {�GB�M��;���3�k{�:I���c8D%��
����w�����wYIK5_���%j_��ntm�y�6\��E炀*�ɝk�<+M1q�Kl�����S���F:�dĆ�s��(M��u6fmӿ-} ��)���7��HHb�]��ޕi:w/�j(C�P��2 �2��e(C�P�8���v�p}wo=�D��7� ��; #�vDn�@��s�K�s�� D�y��wx��'���'g?��?}�񧞌/^x�O>�ugkk�����q�Fs�������յ����_�օ���f��ËEw��:��::q!���ڻő#V��8�-ZS�-q0��Du�D�M���I���,#�x�g���([�/���͠ZӈL�ܤ�0)�+�Ů�R�v��� ^�:���.�QA�P��ȣ�d�FHgC�R"tnܼ!r��#�����9^s��� Ҏ��'����k��`�p<n!.�����;Q��\���7����&�����e}D��� ��P̱��R�G�--*�DdEq�I��t�N�X��G�vn5��&=#Gg�3�۱ɼ#��������<6ٹ��<�#2�/�p���!o��k�0 ��^U��02+�1h�u��IN�U�t���~�Y�:#!:�����w|�/��(��E97ԃ����P8���賴h-y-�U� [�';I'�'�Z�6w$�{�`�9���R7����!�g=]�~��޽��f �|�4e�&��Sg^���+m��m������܇�9�Y_C�ZȆ�_�r�:�d��i�K?��4�a�[IT�;�Yj��t͇z���Ʒ@jL�J��%��IQe��=r?�
�GG�o)��H񑾟N'xζ��%4��j;�O�� �E��î���cLWD�B%�qԽ�U-�(X4�.=x��~�i�x�|�LRbg?�:q�,d�ı�
��7���X�3��s��yI���i~�$���Rp�vnCQ �9"Xq����V+�>��<ǩ8��-��@Z(�x�����<s�5�\��*)��2�d ee�r�j�E
��� +�ey��Ej���E��X��o����[lH�!y�R�O="-�rDgv��@�+��FP�ib ���{)��"��^"�j�Yf�
`h`*Q[�M�pyl�s��ڣ �=x,����٥�� P��@�Cɍ<��I
P� Xں�0@ ]�H���"�ISG���u�N�H!2M�@�y��k��2���ɺ/{�y�v"�(gRaD�C�c.vw1�Mf%������
%j>�z�=K�s� *:'�j\B%@%�m�C$)�8����g*��^�Ƿ/����3�]�+���)(��]�]�׌�;�Y�򇲟�b����P�`Ėe%����ꓥ}����#{�{����+���<������Y�S�.��8:}O�Օ�����r�b_����GhA2;)�*���@��-�@�i<x�c������D������gWҊ �~A��HS���}�`���/�~��~M�>G��c�Ti����@?�����<pdD
uƦv��d��$������K/�@�����lq���9�џ����`�O�ϛ֑Dd�!{]��G�+`o�&�����o{�EN-��!�?ɠ�3;*�oN�4O{�l_s�5�f/1���G�і��Y�
Q��zU��PMa�w����O����Q�Yzx��驧���3Q������w��U�>�����˗a��) :UJ	�{x-�y���}�~�sȺ#�Z����9B�񶺴��Ur������4z^�FE�ھ��<��=)�@�4^%��� �
��~J2.�$�Ȳ���B֜.+@h��H*�Z7R�|��X��p��k���^�֛�w��B����X[��`?a=��e�g�U	�Nz��+y��=���P	D��!9=^ީ@#y���4n�J�@ �P�򽗁 0��e(C�P���),?���];9>^g���*�'�hq$d�< �N_��DG�ͬ�}��K��p�G�QzQ?s�ڍ��w��F���w�K�~:�;::n�D�7�n�Z:q:��Mz��7`' �D��N��  %�8��/�y^��Ϋ@���k�*�i��8��m��	�l"\"�4��8���#\�<�Ү��1�i���,��Q�d@�k�I�o��B.�rv�?������ɈAS���<���s��sE�!\�`�C�y5�QN��9�һ��,�����B%"xq�"��%Ku�u�hNC��:<���.�G���r>"e,����/��� D�����ky��A.���&��.��J���Lf��Vd�^�U]7Y�,B�F}��z%Q(PŤ�7!�Y��,����b0�rf�l�����
\�g,��"EЪ�V��As�A�>#���ќ�.wa�R"Z����ڼ�'��Ҷ�$�C�2م4�Ȳzu�X�s���D�=��b�k��ѭ[[tw{9�(�H���r�#D�!���F��ն�9��,N�������%�PӢ"��X"|x<Y�A����{�K�أO'A������*��Y.�H<@-�j�� #y%<9�v����x2�
ܞ<gǐY�z!j3 �� N��p�w9�ι}�6�k�l���k�[�v�LR)���F"��\O۷o���۰��8�Q����G,��$��x��Mq>םS,8�Ο;G��
�-��|䜍B�a`c� _GH7qL��ǐ���1���}�~��f�>�<ǯ��:���۷��ܾ�%m��T�E�6�UP�~�B=gk�6��K��Ñ-�e�ҵN�Bj����_Pr_�CfcKJ#׹ʾ���и�Ge'b�M6�#��t�ج�E�?��^!G� T I%Ve'�j�xi7g�E�[��E��i��v����l�[}F&YO��t
�/�q�3�[ol�a�ћ��������삜�D ׉mb�R��>=������ַE/i1@\ ����AL6��յ5���D��)�YD��ԳB���&��I qJZc��7Z��k��Z�d���/�c]�(��}!Бb���}��F4o��R!�YUz�.��k=)�r���_�RN�S��$OL�f�xc9��#�������ɍ�*���]�,/�"<[ս�5�g*.�0	v=��3�n��r�|l�_��E��ߎP�f����Wu%\��P�ʙuS�����Bt���3���P�k��._�|��+{�^	�����G���������3�x����U!I��i��'t��m���}�/>�TC�c!�r�_<Go^�N_����;�����-��
�[ey� Rm��x�������
��gG�}g�r*�����C���z�g�K���G���i�x�� 3�%�!�oc���7n���E��g?M�{���o�x�����*ظ
�$�0�����ǟ���WF��#�#�
�6$v���{~�x�����o;�={�8<8��}߳PE`izT�{M�`y_q���Y�����
���K�;H~G
����f���U�)1w��Y����H{$d~��)�����,�M��U���I�虜���XVﺏ�ȞL�1�&���Q�=�_�Z���(P����U4��4B�m��}0+ H�8!�{�+��S�����HQ�*+fA���(���+6!�{^NUG��F#��[���jG}�d�c$���b��D�ZA�X���A\�v���e�����e(C�_[�P�2��e(C��03���q��F�~�ޡ[��v��E�Op�Yelz�@JO�dї�F�++�xf�w�n�^h�f�9pf���y�=3�Ř��k��>�@;����.^��k�<"󉲌v\҈gˍX!	���.j�EI�&��^^�#3��KT�#�����fg������9�vU���J�I[AZ!H�i�y(5Wgc .
�8i�N�L��*_� `�6\htG��s4�u���H��t~zNHv* k j&�*��"�HA 8f�ώ!d3T01�|?/��5I�xoNoG�E~���@�hH�㚞Ö����9{�T7�I�o��Hy�ؽ�ه�7�.8*ҷ:G���+�.J�.*�����%����bTiB��%�<�E$O,�1�㸾ƺ�CZ:��� ��w�q&cSP�Y� A�;���H����k0�j��[��@���A���1ox5]�ٹ]��^���X�I��䤣/`,p�������cܛ�1��c���˸ǚ�AlG�l�E����2��ui��lUɣa<#�(�����/8X��>�ez��5���ќ	<�'�n&�l ��uN�["�=�I�?����e�M�1��|��x�I�������WhmmM�?�kv2����蹯|���O�$�ߟ��Giw_�PB�;bg̩+�g�/�C��2G��- $A�mPj?O��gh������8�| �d4l_�:LI��^��lc��d�\H�"�A��G襯��Hf�� �3V��y�moo��3���<~���]�r����A>�qj۠��8�˸1��\J4��Ȕ2\�� J*�8.@��ݶ�ť��rJ�]��Ü�Rg"��,^�������+@L>�h�⡂�L޼�|���U~ju��Ĕ�YQƀ�� `r�9UO��7���&�歩TxK��qd(}<o�U�3��m+��=t����Nq�ie@`sF��3����d�(�l���lc�u�羒�^{'�}��(���K��
��e���n��9pD�a%����+��HJ��.i�@oi2zYE��+.���+ �iNq�NN�1�����Ks�2 B�_��:ԣ(��J ���d�d;�c�"������3�pUu�.��Z��wj�d;��߫&�{ ��5���@P��z3Pow�J��y��^K)�T��cE�)����8]t��.�èK\��h��gT}��)��=�Z�=�(m1W���Q_s�������ty<d�ݺ���NKv���sA�pze����9�i,Y�B�F y^����ȇ?B��?���#�<,*4�@u�G\�z�nݺ�T �bHsZ:T#M���������&���nf�����Ru���۷o�.������$f�����_aouu-]{���N��=�9O�<�SH �1YO���l�~UwtM��9�w"#�:�P�w�i)�w�l���φl���``d���>�۷��k������:�����.���D	�@����޿�~��/�C�<B{;�鼣d�g pJ�9R�Iꔠ�s�{���d���T�aݷD���e&Ȼ��Z%oW;b������`��.����OJ ��T�����!�?���U{p�#}�6�<�r:9���^@ǅG$?�1*��J0n	ي�L��0)OljZ��������2��ab���l�.��v����>�c4ꛠ�7�c���Fƛ�xe���G��jv���^z����l�P�2��|e  e(C�P�2�����b����ۣ��l���M���,+_�"�HF@�9]"�iR I~��pG}�]��6�1��W�0�c�=ͽ����*>ǜA�%�Ǝe�d��yي?V3�E˔H�
�Tஸ��ɓe߫((y��� �����Q��X�-�^U]C�It01��<GȎok";�8�s:��
\�D��ߞ?f� ;,ѩN$��Im9u~@jP#L����F�M�`06Gshd�S0�s2U	gd	r��6�JWn��o+P����X����|���
&�ȇ��X��!:�vv,N'��.���P��,�/D�h2�:ޢ9�JzgajXc�J�H�v��U�J��������o�<�Ϳf;#Ԏj�� pQ���=}&�D��4�TV\�U�!�@b>G$e�S<��U���) �@�4Q@�jK���рuu�[��R���8�Fc�Z-�&�<�YݢC��C��$�3K��;Q葷Z���02��"�� 
qy,R��s���R�l(5��\V��o�{p(7*�� +|�g����g>�eZ�E=�xv���,ھ���c#��6��q����g�����}��+/�7��M�<s�6'+t��z��'hmm������R������s�|�r�;���گhd��dMh���e\�(H�Sg(��)h���Inxom.����G:�����IZg��Y��֢/m��3pd��?�s��g>�D�/�ՠ�Q�+�����h+& p#;b�|Y'6��7ms��jn�X�x��,vЩc���Wl-���)i��KQO5HV�2���t��E�(D���t�[�⨪h
8�C�[�a"��}�̓>��f�?���,��)�%���n�'f��ٚ�؏:6��U�Xk��\��U��FF.��[���?߼۶vaO`c��=J^�w!u؞p�??�(��흭4��Z�������p���3 ��97n^���-�v��-t�r�Ƕ�����1���J4�ݔ���0R��Ӻ6j�6^HQ��9ݵU�,�A���l�.cϾ�q��g���{m !&PV�q'k#���5G��/kr7������Qݍ�V���z�-ߗ���L��J��S����s�-g�_Ĺڶ潲|ƻ"�?���S��y��mu��x�(�\l�Ps��B�͓��-�T��kwe�N��퓗��KTm[�ҕH��s�j�m�2�lߣ�=T\������uՉ�T*����c��4�����t4ׯ]��t�i8�^�����s���E��uΟ�5;��v����PvJ���)� nt���$���(Q�i����͎5�Z�f\��1��]��_�_�g[!�q5Å̎m"Vc��<(�������8��`��r������W5�v^Obx��͛�hooQ�w�܁�ҙ�M�8;R�*txg �X�Ν;�t����v3����d���ur|"���$���2I4�9_�G�����(��H� ^pD�G{nSO�� {C�_i�?mAȔ�b�w~7��\k_۫���̕���iFĀB黧�H�>KC0=M[T�l�%=��P�ʄ~D�*r�Jg�|�˻��q-�]��(f��g��%B�_�R��D�����0wl��62�p��m����{O��:�m�Ý���˗�>5w+k�_X�2���;�� 0��e(C�P��*����~��>x�@`�i��#Wt�%��Z��0�c%:��LbAp�@��� �]l�f��N�9"΂�@����Ya/��3��� �v�|���[�c�d�I4��	�~�i����.Pp��MR��:4�]�����?�C��1P� �<a�?���іٱ�r�*�n��z+�f���grwo�r.xR`��b�]dN?q:j$|�*����R�D^�S����%���z��%�ƙcY�k@OMU��Q� ��4:F l	��[�A>p��ȩ�䅽�2NT�gm8���iN7�$z*����59Fhm<#����B"�:`��9E�i)�f�Ng��|
�G�������4Y���zN��ZW��^��H3a w5�EbT�9���g�y�!'jNlu�#2�FL�K�uu��ZS��!�\��/Ѓ�$<GG��N�g����(v�̙3��2���U���ujG��}cc��� �z2�
�s�d�j���i͜��G�lp�;B:9���q " �)j�V/ ՜��\�ce�r��q�P��F���.ϣFe�͹�ux�����~���ҥ�ǭJ�OƓ�>������#
�4W8op>K��6G���Q�e|Q �(+s��<�u���þנ[G��Tec��{꘵h����Z��7N�m�˓��&�m>v�09l�l�:�YI2�]��6`L�3�m�h� 
���%5ج �Й`�x�\��^#���fF�B�E�gژ���vvՙ���|EJ���!3e�zms�����y�1Q���� ]Q��9.Zi�"���J��xiTF�椑&��]�$#�iV�v���"�-�7l����c�6f���kkJ��M��,�?�t�u� �:^��X��a��#�����V3[�������\��|��a��\9*/ }�J�L�������HCi���&P�F���ې9/PJ�\h�d�e�[���H���Bޛ
��<J�Ȫ:���SSƣ�f�@�;�fX�پ+�3l��y��~I_�xظ<��{���nS{i���b�F�+c�"��{��t�\_�;7'r�����m_�M=�mlUY.ݛ�冦��&�'���ߦ��^�#fUo'��ytKU�v�Y����E�w3=��Y˥&S3��˗BԵ����N�Ql?hm$���x>��ږȠۻ��H�F�j������a�)��Q/��]T-� �fm�㞱�'�V�l<�۸��4Kk�Fd{LKꖷ|y� ���4+��N��
�Z���`�-�KcJ���R�h��FF|�e��lȗ
�9��,f۟A\���- �-�t���n.���,���[�}�I�R��8�~i��F����vv�d/��K㜶�#�ǣ��HY�clO.��x��6�� ���<���=�D�W�p��_T�`�[G,g�z�YG��P�kzi�J��~S��QU d�鼭�M!G��^�{x/�>U��7�KJCC�O��9�ҽC����n�b�0{�܃�s�(-ޥ��}�^�A%v� ��>+��}���}B�R�혟!MIZФsӻ ~���@oR���o�qH{��է:�Զ}ڳ�S�k��K�9�����=��o���oFm��N'󕵵ٸiw�;��������;�;#:WuC�P��]�� 0��e(C�P��*]��+u+���L٪�O^����1�}�cT4:�e�F=aN.U��#����y��f�%�0�]M��v���_�� ��K�sI���>��5`����|uJ��@d�k�;	��D(��p�W�HPK$�82�1@���T��V�U`U��H�˒��%�Re�ފ�p4�/�|Zjv$�' �H�g������#�h���5	iξ�%�~=��3�6�����}5��9��H'��K�9�,R�b
>�r���R"���Aږ���LMcj���xҊ�K�{ى5
�-G(Y��r�������{2���:�;�T;xԳ:�#�s,S�{
�ht��*�cU�[�����dMsr�
d�3,�!��ScT�DNPB����8C����7|N��4#4���y�ܔ�щ#���ΐ�����:/,r�IѻMU.��3_�聋����6|��7�A�ԯ�=�H�#��w������1$q�x�q::��{_�v%=�����CA���1�{����m\�#���%���q�:�Ba\(;s|F���p���t��e�N��NftN���|�N��\l`�@1�q��Z��{& ��vv�B��S�����L�j�"��ҋ�]/����<�~�a�z�*���`Ip�E�,OѮ��FU(?��_��� e��m�;�w����|�I@�����*�Y�W5#�����C �`���Xl�^�\-������|����>�~���ZC�3���;�6b�E�u}�X�s���(����&�{P`�N�����A>�!=�+i�-2ʚJ
��}̼��qF���
����� ���K��������1�r��~�E���^�� J��IV�Q��r"�=%���6i��D��m)�n�E�`$��G��1����w����z��#�����_�qR/�&�,�P9I㶟�u%B$�XI+ �Z'
���R���@V9
��)1FMk���w
6-�}��	[�\�9��,s�2�6(����JK̟	)DZ*Q*���Sf������D}��s�T7����$�N}@e*-]�6(��|�{��*��\�@��%�r��\D�����mSۈHy��.��iĿ�ಝ��y	_n�eZ�|���CY�>��Z���mFd�� *�so�pߦ����I��~�d�`m���x�j�E3KKf��\�5
�����k[��{�L����}ʶ���L�nX((i�k:.g
)B��
��&b�["��B6+������齪b	�ۤ5����fc�o�O	hr!)��ry/���$��RŦV����sߖ�`ĭ%�߾õݿD5qBJ�NRz18mv�m�g����˜b�%�G9-כ�}�Ӿ���[�*�=6Ϟ�g��4���C����b&� ��59������w2�o5Y�I�s����M�Ac�ċZ��`Z+"�h�H��cow�Ҿ�a�a�jN1��AHm}�U�_��Y �6MD
-?@Z������]��G�;��"��+�Wُ�v<��h��F�`�p�|lGM�ο��j'#i!�����֏��#L��8�L��#1�xe%���Dn��d�D0N���ޡc�s��p���~�{J�|����ɘ�}�c����x'ܥ�;�#�����e���('�	I��������̧�R�,�s�����wǁ�fne�̙3��Q�:��2���{(`(C�P�2���U����f��zǠ���[,�U�H#���V�?GL�ݢ������S���x]t��2�)!�%s�@¯��b��"J9�Ԝ@A�2�{'Q`s���.�����|�\�Q�@�g�)Os~�� ���s�9��H�r�E0�37mr�@�
`1g�z��PEyQ��HJY0[��cS�@d芄=�2�ų�-�ho����S�b��VcB�rT}7/Na���ݭ�L]�$�6���c�}�eG����!��P���T�[��J�`��H�ϩ���{�jd��D�Q�CY�:���YY�����㘕���r��@ �q��2Km-m�N���wU~R�$ĖZ*\@]��'* v����;���쀴up�S�&V����D3�EIG�(���s3˃j~h�Ǒ5|� �D�&�8�M��`w���qEH��0�b>v:�"*�����/�*�\�v:wfĎv4& �.����Wl{w���4]_G�rގ������^�Dt�� ~i���oD]:g��{�,�ՃLd���s�P&[	�GZWU[ ��sNB�J�q4VlSڽ���(� ��f�{����S�pH�
	�4�'�	�������7o�h����]�|������ߺq$�Gz�._}]�$H��Ev�u=��UI�t��{�e�R���aSb��:*��4CP�
�yS1�ՈHh#3��S���WL�"�/��[&�`\[�(hnY�zk�$�FU�y݌(��r���@�k&���IڃL�V�E&�c8C�v��j О�]�� ��!�z�=]Nk�uv�޴�m/D)�L�1l�(*��Q���3B ��{�����<�j?U͆2@қd��#:�O�!�a���r������5\~�L�LV��XG�:��鼿����v@��b�vX�����A?��l���ɾ��!�ok���}�ζ6��������N�Gư��:�M��a��uJ"�ؼ�vi�Y[[:�屉��]�K���a�K;�
�8E��y
hKE�sI��Ċ&� .uNI�MK�5���.=���<'�}b�.]���8>�z�'�U���U_��K<�8G}W�p���T]�� �����j��p�5�|��q5=�I+}�I�T:�ED9��2�\�:����s���!	gu9��I�<�SY��g�\�֩8��_�艏3-��s��wd������?&k�<_�-��s�"Y���62��b�o1���tL������90�2ɂ�IMA���'%�A9˷j<�*�|T{���y�{.�>�{�N�E��I�-f=eAxW�RV��jL$n���ɔ������NԤ�h��~��0d�tQ�i��H*b��L���;�G���!�	b�^�$l��I<�z%Y��BsM���)䀬��Ą�\:b�Lĭ�Q|%��U�k/�5W��k�����cZ[ߠg�y���ڢ��M���=Y�3���{���LSX��7�L&��$
`�g#6�	���D�1@�&Ux!�k��X[���/� p���[`�r�"���4�B���b�鴟z�h��"���̘%�^E�-�y�,�t����6z�kp����Ґa }4��a�鄶a�}�ީOs ���WU���'a:]I?G���tԏG�~<Iu����x,Q��F÷��`�5�o\h�u�bm�v�g�0�ڐ�8�?Ք'��è���pB�g״~&`9n�&U95��M��y��m �"!b_���<�=�.~o"׿k`��>6xYe� ���盅Ԫ����Ԙ'���hz�̌lC8��e(�c C�P�2��e(o��u]z>��[���C�c�8�����&2�^x�H�e��f�}*�7�_T�T�xs�!�8�G8��t2	Su��A�\t�:҈7��_��+ΦZ�Ԣcq$��\u��mu�����Ѫ���W����)v�\��C}m*�1p��bBm!�Z�L�9r:G|kr߲3��HF��3����vw����T9�S��l#���ɑq�a��T΢P���'��e��\�#~|���Q���O>��J�"\C�>o�c��d)z��|q����<�Q���^���[��~P�,���p�ƭ���	1�*5�!�ɔ����\c�nO�
�����r��H�}XG�G�&ek��1U$���>�֣!�b���E���E��mMP���g$����	W؟ƃ|Ą��4���~e(�%��BK��o�nӴ��͍�ˎٕ:88���c���!�'d@Q*�j�AA��UՊ�]����y�M����u�*lO[\��w|2���bv"�P&sX_9����%�+Nȳ�-�o~�m3Fۏ'�L8��.i�m��߆��'t��!�MZ���Ϥ)u�$Ww<�d2	Z�{���QUƗ���l���������, ���c����:gx��*cQ"I��� �������Rc{N#���Q�Ag�N籪I(XdR�"$�tޑ�f+l���+R�����eb_��O�+����z��Ŏ�_�b�������poT�@���v��c�&�n���J��Xr�R��*k�W��� �>�+v�&_�=sَx�ٻ�&s����ҶTl�ߕ>2���W���ԭ�x�W(i�䀨:�h�E�9�T����ֳJ��Z�%�7_�pTǤ�m%��F*�:^�X_�0��e�����^ٜ�10��fi;뾆�q���>(Q�C�6�"e��_	#����خI����J��;R��x��	ŶĪ�]��.��a�-*��p�˖Q?�f`9�_W������շ�#�)��Z����a«�4���[ ���PZ��8YOr%�Ʃ�kP�=�;Cf�N�qɶ� ��ן��i9�����	��H��+��2Ȁc����[s��N�L�C��9���˸�:��G���5��e�z�ہP.�H�J%��Ƈ��H��Jf�e<��y�yއUk��=�/�7+7v�Hdd�X�r�V%��=�R��3�.�Y��Σ<��ڳnp]���zK���S~��DmK�aJuu�/��T{`]V�H��W��z��N�v��3bMR�ے��c(1loߥ�W�@r��c��]������ p�z��;�t󭨖 ���ލ+0�M�{(����s��: ك5N�)���i`�m��O�⤋6׻�O>u�v������d}t�6�����O��;6%���Yg"���!�Ud@z'	�����q�7#�9/Z�?�3u�5�Lm���!���o��q���?��.��1�t�<}>�>�}��d��s>/4�b� �(�s�}*�4�'M��W��LJ��.r�?<K��T1�����ǿ�c"�2������e(C�P�2�7PA
 ��C��#*�`	��U�z��>9~oR��6�I���.�hNQ;V��Μ3�X�܁z(����:
͑�4�FH�!u� �S�� ���=T�-�Iԑc��T9X���������s[U�`�3(��,9����,����]�\��ה�Ga���5���V��R��*aι�g3:<:"8�C���`���V�2�G�Hs71d�{D6y��Lr?#3 ���8�fv�$PG ��<�6�Hrp��1 �To�N@`��p���ȝF���Mpl'9��)|����|��9��5����Q{�N뱷�	���އ{:��R�j<ʸ��,v��RC<����:3����H u�*�Õ(2.�:���Y�
��.�D^�e������P�\2�ev#���N�P%Dp�Qιz����^j�/-�}����8��i��d�����'����� 	a ��/�a �S���[��!P�p�j�A�ދSD��u�Y�T��F�0'G�.�QK'�Ԇ#ͫ�w�~&o]Y;�-����M��iX��V�iYIe��o���d�BϾ��P_����i2�:-@ ���62����h ��ݪ�xD ����-�0�����_��,X��:[�{���y&��)S�$[���NT)K�PI%���~H9o��Y~��R��*UJ�Uq9��D"CI�M��!pI� �^�����wwz���?����ݨ�{���w���k�o�o�O�ry}Eu�g=���m����Q���G�&�b%}T�(�� �7)QeyQ ���#H 3vXzWdH
ۆ�/u����2X�SИ��m��D{��Gd9�Q��!:FA�Gּ�4��m>b^�y�E�l��K��Hk}*�(�Ӡ�Q�����*a`A��0%s@1͊��N�@Փ��{.#7��*�r��ʱ��;y����|�Ӡ(l���#�=C����z��S��S���D���9D$Lt<u��&Z,��/	qѽQ�i%ZցX��"x���bXj3c%6�>Z(�?��Mۏ\�-�P �t"���FT[Q�E�J*A�%�.*����(s�s �>m�t[�}ܮ候r�.dG��kk:�AƂ�l����1w���t#p2~T�� �,G���g��I���b@�֞�*����]�:�vA����!���1J}_=���a�Q�"�M�0�y;N�8�D���M��(��"`���d��l՝6�L��>�
�3dC� Ӻ>����\���~�*�DY�A�`$�x|c�2�7&֔ξ��,`:���z	D_��\1�9��T�xA
����Q��r C�9c�ֽ�i-����I���N m�Ni�;eh
V��T��A`�9���?���A7�3Y�9��Xy��Һ���S`Z�H@]���
��d�zP�[�_8�R�-!�K�m�#�e�hy 3ѻ�����]ř�W�Ԇ�c6�8p`{sLA��Ϟ����_ݼ��/U�|]ߨ<L����spڽ	u�G/+j�?��������6 �!R�UD�_�HQ�j�w�����<m�H@���3$J�4J�M������<ha��u��_�k�����������[���W�� }�[��ַ���owX#j@q	P(�����3�"x�^����9�o,3. ��:^rH{s1q�����accv�i��㉏�?y���
4��T� �h'�RnKt���.��:���A��#t�vqu6�S���9��̉�)�}
Jj_�Mm�<��iκD�~�,�WC��r>'ώ+�M����,�����8e3� �M?TB�sP ���lQ�����c�ϙ}�"�3-4ִLo�Bv�5Q���}Wqeٻ12�DlC1��ݓ����2��Y��FZ��ln�t,h��8{�������}v�6�ʕ�a:=��k�� �T��܎m��׺f$��@]��?�s��q+�<�{����L�����#_�D��e��u��f^��>ZV;g�5��N���Ɯ���=Z�΋�8�߬(KS��F��v�n��>�Ų�Z���(O�����V�����E�s ��b��W���$!gp����:��n�&- ��Э���@����% JafrL�5�9cG��:w�ߺK��[��v}
�6eM��]%�Yev�`tzޛ7o���g	d�{��p�6���>���:�f� z��[{dӝ�(���6�c�[�]��WN;�m%�f��{F<}^�0 �4��Ŝէ�
u7�tLհ��9��>�`k䔿W ����!p�GE�*Nօ�M�!�S�5�!����ns��|K`2+K�F[5�Ρ3G�U�PI�UԪ���P9W`pY�Ө�����q��LtM��/Ε��f��d�I����6�]}�x�5�)0K|PIy6ʦ������s���=��te�����~����_g<�8����
���wm�w��&���58�<7良4TfE4���V���EZ/�.AQK��5�5�EK�<(�Wf[w1@�P�ld��`f{H�:��}(e�����`�=О��C�e�6U�X�E'w��꽵G�5`�E�\g�L���ϲe��A$X&и�"����7`�<�{��N8�?N�c��Ӟ�JS�Z ��]��I6�o�oʘ���!�?^ �"���.Q�P��2��	�E��Nԛ�K,�s|�G.\����6pr�Mp��fX�&���tPs_��������'�.���ֱ~_�o��1^S�j{�=T�)3�� }	�5B6�nc��tV��9��l%�1AK��*'�;�!2�����֓���@3�=ך؄�`�"����{J7�T��~��s�o�&Jz1OŜ��s�����\v���.1��(�m�V�O硣�Lw��%�tT2:�H�E��Gw�����@f��J6�2�R^�l��Km�J�C�vq2���2�+�j���!�ے"�I&Y#Fc!"���۠��B��5�6�el���ho��ݏ�1���g0q/œ˗/.A�
������o}�+�� ����o}�[��ַ;�aT|�";���^?s�ٌ��B�Jn� T��i��2 hMq��LΒ���a�3(� g{���厀9T��
uHk3g�˙)���뙣�Y�FyHԲ����P��7��x>K��R2���@r��@k���O�O�M�u��g$Y�0�3q�?KF1�C��q%PI�⌤�Ɯ����sKc�S��kd�P�;Q��۟Kjoɶ%Ѕ�S"����-0#_�2��97�i��W�|͖��c��\/U齵��:n�)����)PҶ
��(��j���À2j�1�S�3x�\�����2α�'e`S� �|�֨�sV����ey]�\�<;���_��!Nj��Bfdm��`�|u��9m��%����X�PiVa���yl����PT��@H�����e�.Q\!�iiL1k
�(����NN����38��H�\2{����4�%P��tQ���vBI�>~~F���^�e.��cZܵ��t�����2�G� 3��!����<��*j��z����{DE$ ���YO�ŜƊ\�m0�i�_���ia��h�g''0H�"G0�a����+��(�jU��̠Ar�����汼M3 �sdZ}�9,�+d�)B�:�Z��I�������f.�U$;�=���>�İ����\J��M�΀v+<�`��<�����f0G� '@�1)�`�S��6@��@���C��S�Z�ksU��ݽ�-D� �BK����gWV����$H�ʗ�(�e��#e4���y�	E� H(��O��9��w�o36��Y� Eh�-�09ЖA!�[�:����-꾏sY���Z�@+�9�򙎳�7g�����b�h��L��~(�#��h45�̂��f�,�.Q�$`(���%�nA��o��d<sG���l����;�=�.��u�Ʒ�%� ��*�g
�a���q4TN���8�.eVDi��9e�M�0��u?��Y7��R��HS�c�m���/|^�y�<w�<����Oa�TF'�����Ʋ���4�爚9�re�����/�~fb,6�Sud�� �F��h�>����߄���߁ٍ�����~����;�~��8�
��YE�|Ad�z[[�),��]R|����Lv?P}�N-���s���(%�4 ��^˙�XB�l&eUX`���כ\�5����t��`k��IX,;�\�l���ʋ��e-زR{"�\�C;�v�;��ե�k���v�d����������@�c��eż1��+��x�	W�7�j^�e��tόL��'�.����z��D��b'#O��'��#�#�d0[�-���8P�ڑ��[ٷ�=߭����`8.����4p#R9L����`c��\Z��lX��~X�l��l����0`��ZB}�[��ַ��� �[��ַ���o}��' ��;S��s�Ď"���JyȓK ��R�ĘIL�8��S�AmM���RG;Rל��U0B3�Z�u<���+2(���Dӣɿh.ghW�m�QL�/\N��~��	2�6�`T�g��.;�ؙ]�㲇:�יz!�!�W� Tg5RM"�+>������|}{�J HX*��l�RF���\��\
�I���*��s �L�Ԃ8T��r�>������͙��|�����Z�e+��޹f15+2�la����ի���Q
XA]�x�hބ����"��u��*A�}ԕ�(����f�˄�������B��c;`O��nw9��;�"���Ut�h#/#��S��j=Wp�pvʒ�" MFc���&��<@���ջ��	GG�p2=��r+�����,�<N際
F0���_3��G�� ep��՚�"�(�^2��;���9��f+ȕiFdA��ٹ&�$K��5��
*c<�\� ��9Ve�	w̐��a��|�~�ڜ�k������|vwwaoo^��p����1����Z��)���f��ܹsp��5rH�d|K�;��%��r-��+��w}����/�ㄦ�P��A���@�������"�?J`9�%M�o��,��:�>���佩5�B�� &�	�q������ ����3N9<Ǫ��|տ�����\��@�������Lï用Qٗb��;�M��mht����h�`*����>�s;���vE�9�[.�Lk�Ԗ�k�k)sJgO��%�f��ۘE�v����Q�|�L,Pn)��l�u
���`�F/3t5(�4��c ���ו���Zv*�J����G�_�w6�x����s�S�k!��N*�LU���*X��>�2h�P�<�hD��|��D���$��������q%,',5�i4	��TCܦ}������EW�Y�^�,Y�f�h�yn~w=�^����
'Cx�{~|�:ll��pX�Ԧ�jZ*�\�^��m&ԎE�I��P%����8'�4x���:j�ƒ��ষ�/~	�x�����h���7�IWc�����:��Dyc{�E\L�ڼ�sq�9)?�ړ`kU[� #ol0Nm;;�!5R29�� �J�"Au������ b�e�4 ���z:^[���_�ڡm��|\;{/����u�_�o,���+�:wmt��c�s:5):}i�LO�'Xk�E���6��*�\��Cג��`{[�婌Y����=�l,b�K�Cj�iɡ"�OX�TFTcU#��c��4h$�H�'���	�4"'5���oOz�W1���f��S�GS��=Ǒ�����o}��[ з���o}�[��v6�؅�D�d�ys��@i�� J�*��8�8L�CG�Fy�#Յf�B0'I�ɦ`Q�a���9kрg��u�X:���aeǲ:ƨ�۟2�$��Qr���^;g�KW\�M+�t�����,�]�αp�i������-�s 7l`*�@�Y�ʷ�3�������@W��e���f�������B�$%9���h��B��dJK��@��6�]�kΣӴ��Ŝ�n@��S�T#tE���`T�1f���Y@�������T���:պ�Ē!��A����s�{�4,���SG��ug�1�x����Zn�9>�����\
Б3�y ?�P˲#ڂ������]���J=��L�:<<�ãC��fiA���d���l6���c�������7��ʀ�a_-�,PɓÔ�L�ѡ� G�-�kn�a=L�4��e<�`< y�$���LE��=�^AZ�1!����D�q�A�NgU&���Ꙣ��p��|��>>�0���\���_����8��<�����9$����*��+�{^��9P`��RE0������q3�z`��J[X�BW)��R+�|.a!o�|���gϝ������h�[["k̨��:s���p�'��c���>��[J�6�@�h\P�ЉO���
�˂�J@�(z�GщXIkVu� fQ��xlL�˞G���I�#Xђ/k�%lf�,p�	��A=��`�D� �u�&� �͟�>d�Z��>�ͦ�m���������y�;��Wt,`�d���,^�l[��r�A	y:TB�bAv=W<���T
�ؼ;`X	��;���^P����c�CEƻ�n��'�i�3}��;�@ʖ�{��ߑN�^�w���x����k����a��D 5s�9�X�&��J���8�hЄ��m���)��%ؖ/�AC���ˋ��&�ʖ������<���l�)8��c����J�gk��#��*¥G���7��ξ`wg�KJq�2'َP��%���e���J~��l>'����ſ.���/:�M]�a��=ޅso{|�_��b��> ������F�� Ԁ1�u���0��"k^ǰ�1���tWl��JvkP]��/[TY�8enQ=��-�a,`E������$B>�~X��1����C�[TƝ�Le��akc�[t��K�|_�W�Z�u�2�1�2 :�$?!� �H�4��,���Q��T�`ly+eP�V�	�M�)�N�rO��%e�����l8�ihpMת<��H t��
����^u�0�a�5Ջf���ҡ�o$@Ee�5 W'K��O��0��`��ﺵ��o}�[����> �o}�[��ַ���k����*f'�:�J�Bu(�G�d)�oG���7&Y�t� ( �~�"}�_@�#N;��Y���(����iv*���Bޑ�j��x��}����c�si��Fm�;W8�c���o�;dr��=l$:NM��,��(�q�J��Ҙ�u0�Ư���Opĉ�J����D��9�h�	���S����L?H19��,�/d
y8kmm`z��.N}uq^	��}"4;Ͻ9�8���H:0�-
�Dc��@�A��ں1��2kI��P X��2d�n����͆T��9Ǵ�]���yS�̀DƭQPQ)�����Q����ˀ�rڠ��*x�'L����pS�@��*+Q�j�\S�I!b^7���qC*���}^�a<���lp||���Lj���5�bm�f�������tF���/�DY������kW�JІ'p�x(g��>H���c�� ��ZW�^# |sk�뎓�Xdz������4��:x�Y��P��` Aå����l ��P���4�����;� �7^�&��¥�/���m����7�XL%�@���_8G�@�����=Y��/���}PL�xP �!pItFK�֡nV�����)`�DJ~p��qN�໤�c�1�<�0ln�g��Jù\��N��:�az���C�Z�@�����P�w�$E�D���f��� �X�E	��ǫ�R���fb*|S� �Z.k��ӊ�(Z���5�#�4�����y,�� -мX�\�7y�R����V`�<=h����Q%�Bd��*g:�281�$����@)>_���Xj��\p�nB�%����pW����7 (Ƥ�e��xp���,�NX�9�m�e��y]�>b6��� Z����ȸh������4�K��A���4���J�'_/H?<r�=Xxo���ըACk}-KEɧ����d�:�H �Ӟ,sg��MR�<zP��4���h�Q�.�-���FS�љN�Se~֦'Z��.�\�ųB��Ӓ������Ӑ��A��4��{��,|����w�����_��~� 撚���]h�5��;@'��yS�5M�jR�ީ6�A������I�#�S�d��?9��]��E8�I:vĊ�:O��.[�B����$[�kc��X�Ʋ\'k��-�f��H3I	 �K��� 2��(@�u̠�j0��B�ۚT��t��u�����mS&0+.��P����&k��	*��_t������ �kH�f3�5�_omc]�/�~��P�-��%�$��� m+��\�(�oO��NͿ�����T%��,�4=9�@B�g�("�Ɩ��MW�rຕ�*��:���\Р��/ 
�u ,���$ �JW�}M�D�+��@p
�F�3�f���^����۷���o}��[ з���o}�[��v���G�L[%]���Ù��ڑ��f�B��sfq�N�8K r&W�)�}Ɏo� �e3��["� 0�>P���m�C.��q@�i��)z���s�}30k�Nǳ3�()7j��Z_r�t�O����A+�G�Q��@��^�Yg �)�L+�.�|����@	���ɜ��Cr���Mc�E �1;�v��%�?���Ub(s%sR+��tQ2 ���!dw�<79�bїbzܡ�������"�� �� P6=�b��� �X�q�~\���^1u�:x�¿� ���vB�<F�iv�wJ���)�E�D�t������1�k���t�K�2��b�����v�@�8֚�Z:D��<�G>�x���h,�����]~"��l�����{��'K㾄7�|��q^y�5X.�ppp ��M�MOh^���S]w�+_�X���G��F����z��gΝ���]���ؘ����J�=�d�5DS�٦���hcG�p4]��� ���5��`8�M�nO}�\�,}���%�i�+OǱ�ۻu+=�1��|:Oc�of���������y��uʐ�z�*����x~� �.�s]���ٳ�`�L$�nݺI���
`;f�p�+pAf��2��:Ԟ�;��N����'ao���4t���4��T�$��Bߋ�H%>�TαP�#H�BA_pM1 Q�H�ԬV��o�H�F�R����
�h0�U)�O����ܱX�tfT���%C j̺Iײ�(�D�]P=�
�K@�w��E���|�3�c�9(�6B�׀į겔I�2�R���� �,�������,����#}�X⼗L
<6fF�F��{�	˼��M�
���e;��K�N+�Z� *��]��e��]`?Yٖ����h�6Fw����X��]%X� �
��J�ˌ�t��`���l�_͒�!�ل8���{�Y�+֬����(�
�m�W>����@�u�lD��;W�P:��lT2����� t鲭zWȰ�C��撵]��&���,��L���aKTR [-�;�/�8e;S	d�H��>������������]�r ��n���Z��������!�=�ձ]��" ����AH�����fV$*˒l0���¹8<؄{��y8���6�D-酠ϥk����cC�mdd�̀s�[ձ�T�_Ν>7����`ikI`��q�����5(�B�X�#���A|���I������>�2�P���6j~&	�M_��i��'��v�=s1>�[eݤR)�(+�+���Q���;é�T��\>��(g}� \�m8����p��Aj�A����d��^��@���֭L��h�`p[]��S�Fv���{=�Oł�N���H��ί0��J���b���Gye���r��t}���_D��8l�)*�!H0��`�d���U ��� �ַ���'�� }�[��ַ���owV�m�E���3s�xbWS#�;sJ��824�ɉ㟓b��Q� X��
�b��ԥ�@���f)E���z0����
x��Cw*��QG�;��^��<�d��-�h���{l���Ӿ�o�J� k� ��2g͙�=�S6Du�3�g�,tPa���1 F]D.6�<�M�:�؉Ԑ�_�V^*�=řDd�Z��˚���(�J�����N)�]�UiqL��Z��Z+S�*4b̝���A�>��l�Gv����cP�4�"�B��Dհ�<+89�$�Ǭ�����T`/�L�P<����7�����B���b#��fM�Í�|1Q��A%[���"r�Y��09C� uHz�S�P^�r����(#��`��c����<��������vp�-��?s��	�i��$�+���LC;���)<��C�\����'GS�ƣQ:oI�h���N�^�ŏ�s}rrL�֎��7�����'ny����]��~�cp��{�z�#�u�%�@�+�A�V�h��1o\}�|���,����p�};��~$�~�7~}�1�jr>c��t6�7�݀��#����=88ܗ�HwK�����\�x�!��'~�_}���Ȱ����H��]���U���~�}��E��G,��Q5��gw���8˜G��>��O���������5�AE�;
��{��2��<��8b  ����"���.��st��z��l�Œ��J� ta��� ��_���{/�X"�dn�S\���|2�1��<��͝�Gק��Lo�Ak���'(`��8��j(d]	�'֧�]�ҟ���qy|-���W|�`���yc����4ݤt}�k��� `u�i��y	��c��1�˱���>5���u�7�v4-���|e<���0k��Ŭ�5ostմ��j��Ub��n���Jͯ��М�����b��~��DaP��NU�Xjtl�MM�Q�6י`L���f����SW�P��')��ZZ'd�;����8��Ps�i�˺F}S��C:�ưJc0��� =H�ttE{낃���֔b����̕�",�xi�)�h�eH' ��6�:�B�/%t��l�*�ט�b�߸��+�(Z)�Ș�/�v�j	�h Ue,9�pxZ�Iw���|�C'�==�0���W��_�Z���]��0h�9o^l�I h�M�d��ZX� Y;hhӬ����iY���gr2�L1,��8���+��~�;��}���F.�#�W�TFb��
�a̠w�֕�)3�R�G�W�]�b��.1�e��С� �̘Bc�a�y�z�������Nr���s&}�7D��7	�ˁ!ˣ}���#�6�.��<f�R<yɺ�y����O)�e��u��hg�o�;3��M-���p 	�O-r_SpdM6�&��/��3���a�Y6"����-�ˢe�=;pttl�c�UJQ馸��
�%c AO$8w��ֽ��l��	���V6�6?�����Bl�6�f�h�YYY�9-�� J���i!wH;t�]�Nz����ַ���owx� �ַ���o}�[����%��e���	��i�\��"K�(��%U�)�WFr @��A�`f̧������s|������#�XfWv�ܟ�Ǩo�|q����A�޺�ٹ-��:s� 
uB�ik����%�;��lg`OX��8��%��!�lL�����r�L$Ў_
t��T�0K�x���"ǭ*o�'ԧ�Ҁ ��#���NS�]X�q�.m`�q0�cП�5�3@��h��
���;ם��dB�	��t<#}x�XP@>g����[ߡ�@��α�E�%$� �a�'�:�]���j���M�z���h�Wen@�$[ZW�p���	���u۲�=���F�I ��F�`�ch��{���_�U��l:���O�'bKh\kB0(��k����Å�`��1��/�J#�Y�_�tΝ;C��~xxH4�D������`8�-�'�w��Ex��?M5�IV$+�!���ߗ��%q��'�s��x�)��� ]�r��2}�Ԧm��Dh9�,��#��^{�u`��&p�@��n�O^��=��c�c��?�C��ށ��C��!9� ?>�`��P(8�+j8@ǻԌ��ܔ��b�f#z�!a.��\�omo{=�x~����M���e�WDI�	������{�3in�S@G-A2
��>S���X4������c������Ȣ �z�ʚ`������b1#}��#S}sPR�^�{�Q
jI�v�gu�V�$�-���|��I���tlT�AY�|��������M¶��Q��=�	uU�.�۝��Z�C>b�
]`��z�̽��.!�
��<��]\�d*_C�N�X`�3�=��&��v3�#0]p�d��!�5N(S��*�#�[�p.z{�R yx��`�|�۳�"o2J%c�\��-��n[�I_���(��#��������.Y�4�����)��+ȃ@?��5�6�P/��VX^9LV4�<���1Щ� l��M�$=y2;I:iDt�C?�,�YZ��Gi';�>�D�]�Q 1�oft�qt��~�m���#���`�@�(�D"���J:�\td7[w&�k�D��WXoN�6�R�K)�'h!
�0p����:'=����`������ux������������G��Ɵ65�	��X���+^�ߖK��9Os�D�EZS��)ĝ��:�! [�3�W��� �{�L[�]՗�B���1쎨���uc��y�Y:��X��O��*l�B�@tQ���8r�xy��p����s/�G��߂����2��I�vtY�K�0er��T�YW�B��������ֶĤ%Y�܁y��Pj_(�G�$���51�N�\�o��4�`�^^�a�����܀�l1O �`R�������|�;����prrHA�X��#fx�tߡ b\;-���Xx<1h���-��%�|�}� ����xL���6qKe��ųWƶ��#��	 �9�u��>B�Z�����SRγ!�A:�������Y��o}�[�~BZ з���o}�[��v�5�Ew�_j�Fau�lEE��k���H(� :	2ء���8��$�+�^R���qP�3Vѱp^�{,�^�����^S�����c0@�����9t�A�u�u�������Z>�KA��e삓��ȮV�9N��aF1��Z4�u�;eB�L�F�nZ�p��9vu"�G��jgR�}��au��8���[Tp��+�,Ǡ�B�����.�E�ȴ���NAtL߸~��>��4�x��z�9+�{��2��TN� A�X%̌�צ��T��@���Z��P���|m����������U�"sF����D���E�J��lU ?=�k�s��X��2J_�L�E�k �30I35+��m�et!���2pʙ����zqPQ
Ҋ����)S�q�Z��3E`e
e���ށcjV�4�GGG�,�s� �sH^,gjS�i�� .f�������AM�Ә!=5޿�B�y8`��#2p�ɘ2�uM#;�
b�`�c[��ֱN��PY�g��12$���p,��'�3��w��=,X.V�Z�`4�P��
�O23J�$ʤ*w�R�1c}|��
ؓ<K69��� Kk���N�<L��\[0���}��q(P���1�� 
@CB*��ۆ_��_J�ؤ>UBM?����+x�z�=��w��I��ߣy��͔��`���VS:2�$���ZnRZ��U1�" ����Q����'g{���0׻�ļu}:UY'��)�1`�ĂM���8�B�S�,�b����y�Mu���9� z^�	݈�r��#�w�A�9��l��~i�M��i?��
0�R�罯5�#��F�R�Z�����!ˆ��;�D����?���̶��_u�g��Y�����]����F�BQ�Bm o�R�7�5����s�����Q��>�	���Һ���%ꙍ����g+�'!����3���.���ٻ��~�o����'�Sx���a�8AG�����pϽ�����(�y�
�����Z�����V`*kȦ�,3T��ڍQ�I��gG��e[Sב�)YT���y̶�}*��d���b�K	�_��s1��E1�E�����|E�ujS�\&]��ԉۀ���8���?���08?��*�%��� dl%�_�k�����!��G��l����;�]1:�=�fD�Y�-S����Pn1�*]kr�A8lp��H�&P����<SG��/��S��o���Ԋ>ͯ>9hG������I��]q�hsB�'�"��B���.L�.����;�Կ����~���t}f 7Z'�+�b{33L����9��M��S~�̎˺I���Փ��[�T��`:'ʳ[))���zP��~�%n*�ǃ�tN�w�_X���~g� #��(�<m���Ւʾ�=�r�b,k*��Mv����M��:�����ֈyh@�%	��b�h�P����%�=����k�E��{�;��(v#��D��;s&{�[	_3��oh'r�\��%Y������o}��OR� �ַ���o}�[��6`@/z�9��/`D�:���F����Mi�ŋ�Y�~��|A�0�\Y��BV�8� �k�*�C�%��O��KG�P^�V�����:W�ߝ9��w�wv�U
G�w�^����Az5�Ikԣ�3YF�||���S_�Z-9�d3䤢l����j5C*f�.���l�7�)�@=��HO^Qf��Uϙ�<N:��M�f�W0��_�}o�>�2���ܦ����M���_s�����	�>���S'i���N9�(e�G���8qdF] �ii��ػ�(�,]���L>^�^��U)�8�S�[\��T�.r�U���=�k���r�2	9����#�<��RT�]�:]1���3E.H�w  �{�ZV]7��d�������m� {��g�G���|Aw�Z�H�z|�~Nfp��-�߿G�'p3��ry|tȠ��G�A'1e\Iv:! ��	�E�
�ض�EJ�H�/`�!��T�Y�ZaSȠz����s��i�w�6	��n)��fq�<G�#9ĘO4�J�ފ�x	
a�K|TIN�vۧ�$��A%O�\�A)~��7�I���2o�%�k������6��-SP���������kTs��:pd���a��<eSMq�bg�����P�#�Ի���x�'`ww��	��7��P���[{p��U��� ?x�0.� ,���:���^p.��)h�=���yDQk`M�}D�I���N�&��`�(��ٚ.p�����e�
4�-���\����,��S�����k�w#轺�t�X�t�C������*cO+z�T�ֈG5�+:O �M�Yղ���V� H/�\��:g�A�3���cfv��(���l.�m�2@@���n�PK̠�|l*�\����czo-7��p�jzV�Um����x��}4����ԃll��3��4<�䓔A��'�N���?N�?'=p���'��K_�2̒�/�p�=����X��?�X,=|�k_�+;����Νۂ���p��Mx��0J�ӵ^-y�Ř�h�<��X�ZM�WC�7y�T���R��lL���z���g)�<n���\��C]��f��zrp��
����F ,�<��zr����4��6a��g��[��o>���.�v�m�������$�>����;9�х�L0aI�i�j��O�>�8�g��P��xs������ڈ�Qc�ڗi�!�8��L�g�$�f���(�\1b:�NeA �(i�AI�֑��kK��Z�fi��|~!��o�'��u��d^ima�ڧ�E�`c�k��WWހfz�����H�T�1�Q�]A�/�Sť��.f�	"i�׵�����nc�؁N
��%��oc˺��� `�y��ה:���\��I܃`����������d���6\-g4gdي>D{��ߌ�g��b��g�6���^�2�@�x��T
>@�)���j,;�$�N�C�Y8���e)`ى4��]��Xmd���"�N*�����D�w��g�jx��(����o}�۝�� ����o}�[��ַ;�Q&K��1�Ī�f0�.�"{�p�s��`�DQzw��e�߳�q�f���� �w���=+3#�Z���o`R0R?.i2OSfv���H���1��D�X��ԛ���siF���o	=�����%U/߯36�����>�&�S�,�m�?���j�� ���j�zQƮ `����1�nq�4H���7xy��K�WL׉@ah�1���ł�tΦK�Jfyb �!����_<�k���";��4�6ąXAq�.�9�@u�x����Oe��a_˱�+o�pB��:b_���#�A�~X�g�4ƍ��9��	N��v48Lp�e R3f�\���xei�P� ����u̲� '��a�T^"{�%S�f0��Ft�O 9]9�[�oё� S�r6��e������.�}	���n��dB4�^��1�=$Y	�b��jِ�\�z��g_�/���)�%������������3�#"T;3s�����*�,Ҽ-��o�iۈ7<��4%1cp� �Yȑ�խ�,�"�T�� N��u|)C�����?8V����ӊ�>����c�>[[[Px���PW���&pͷ� ��]�u�}��g?���TS��'���A��a:�(z$0 ������l$#Rk~ss"%�\�w��j
2PА��J�+?������x<���L��"t���c��w��?�qz>��2#^�a HpM�A���ϋ}^�Z�1���r@�W8��u��Њ  
���˿���ٷb^�F�4����]�s	��q�Ew7�ߣ(Dt��N7`)B��Q�4�+
H�����#�� *��6|�h��7ԃ|i	�qҷ�s�.V;Fh�5� >�X*��|�������6��k�(`s�<rd��m:pXe��o�1h8̮a=��E�Nj��CkY?�_��6��!�[U����1�W��.�}<�����{���o.�u.\�n�݂Ãcx�;�	�M������y���ÿ>� |��W^;B����TC���w`{s�ο�߸��G��4��:�[�)��e��IZFD�or��� ��E23��Ahe��<��kG�,]��)�ap�b��Me�ŉ�-�u�\�M���.�Lxej�g�q�Λ���DW�3����Eظ�q8wt_��'�ُ~�g����r�V�=jr�I"�G9� R����'�IG6�V��W�
�8��,�ڋ�@���!2�lm����Qٱ����h9��ͤ�w�P+7��m�&�W�q&��+	X�®�hC/��B���ǔ%fMnnӜ^S�I
Yǥ�����]�5^�
6�w�f�5�L���C�=�}�+IUM�5�vbW��Ƣ�"�ٕ_:ϰ��2�YG��G!�tj�n���Jl�弈��w^Wb3��� �����9�v��!�H��6 ����G��w�f�L���0�8�|h�`����qz����Ɂ��l$@�4hiI���~�r^)Ì��9	 V�]��,w��ӗ����@'�����+��yf,����e�V��vհ�j���cgn��;���|��L~gaa�M�B��h����o}�۝�� ����o}�[��ַ;�yh�V�h%��Q x�H츈�9*�����	�u8��,��e��?���ó3�T׀V�=Ҏ)�92J�����qȠ=�1��Iv�����z�f����>����yq�g�>�������迍_���@��p��Y8����ƣ!�S��ܠzۻ�g4S4�����,\�NF�2eӠS�h���⨢,Jt^U�4�Ģ��ā�"��3�W� �yo^�	�n�b�"P�xZߙ�]��q0 
xQRj��#�C��S�V��:�J��T�y�`q�e[�y!}�U�-�+$�����e�f`C�l�P�sQ���*	��&�\C, E�&��\��~�N@�,��D�2h´̒UU^3�K���>1�
���϶�+j?��C@iJ��1S�����$�͒�0�B��px4K�8! yH�' T�Ӕ@0Ǚ�,�u�.���e�� 

6���ZV#ژF
���L9��Ǩ,�#�D�/����� Y`��,#��^S�t��T�����ڎ��xM��AE�eKuE�{��U�/���]�z<���0�)A0�#^����n A
MÀ�R1(��ՠ��Ɛ�rD���<���T^e������]xr�8Í1�פ��@ ��(�;�@�L���'٫Q�O-p����gV�����pa�1�c�X��S�Q��W�@
TH���m��5&㍴&YWZ�TuG^���(��na�)uv
���ft�;��c� ��X`  ��}�_�$�3@���S���;$��͸ST����>��-�z J`��@^��Ry�	�>��5X���(3��eC�EbU�s�>0���z�e.א�L�i�P�$�씽 }qt�$���~�~9������򙲬�Й�+`�٢�N	8g{^1�1g>H-9�����m���5�Y�X���5H�;�5���}���J������v�Yr A�l����{�}�Ի����1�-�@y��G�ڍ=x�wQ��8�;�� �����#�q�:���� ����?������x7��6��&ϩ���Hu���zqP���A�E[rm�tv<؞�� Tg2F�y�[��������)Q�f
������bE�E�vc� �e\ɞ�2T�D���<d�qpR����Ux��~�����O}��d�XR�/��&��e�F-��2"�y'u�q�p}�χ�!���~�{�$���$3ˣ)�n�	�j�yҫ�$O���t��~�[0�о./��f���`�փ�5����&8S��:3l��R��:=>�X�)	*?fKf[N4�SߝJU�MP�!S���ds����4��'���T>A���O�@��1��1��ߙ�N�ZH��1��&���K8�����
v[սv_	�q :���X��v7��A��@[�#�������%��>�ߢ̓�1J��� �rG��3(��Z.�Sp�'�A�Ɍ�UX�� ֭UVko���ȲFs4P�����K�3�ֱR�)X�^g*~k�6�: B�7�R�����	:�̗��Qy �x�h����o}���� ����o}�[��ַ;���bW�XVz�\�RY�@'j,��F �9ɜ}��ۚ��}��ţB��G郃��R�����o��p���N8�HT�?�.e�n(��[ �% ����� �8K��8�ם�|��7N	(0�凊3��3q-W���z�w_�~��>�cX�氽�I� �Fc�������L�M�t!̤�/f!�:��3T�9=``��Whٙ�`�2����Œ���UHןí[�p��&���`�ΫVu�UB�π(e1"m�8��ФZ��:���5BE�ÄR��NV�L���|qMxu�9�����W�m沔̎l���A�2]sRB��9�5 ANtliy����KY@�`�Dp���[v���Gr����:�r���γȿ�KW:C��},Ɩ��6����NRB4�x�X�����%#Zs�r����lsxhZ��ڽ4��Ŋ3��5�� ����2H u���
5�y/l(��Lxd�X5^�|��n�؃���%��w_��������1K�K7 x���1 �g-e�`�|����c�����bc��Y�Q`�,���f�k��hz折=�P
^qtG� H�{%�|
�0 �����W��o$}��#@Q �!�@��k�BO 	�@xmX"�V��=��D�]SQN��@f^�K��˥G8�%0�v����D~�mo���߻�����L��,H����%�I�<��M�Ǥ��3�7WIV^x���O~��h�
���	���;v�s`�7ݛG��.��R
��r��U0 ksc��D�b,�0�\�l�|���z�N�[����3��F�,J�XƦ Ԫ�uo�
��@3�A9̘�]E��oA��#��8֋tDq�VԸ�1�D� �֬�%=>?��qph�(_{>��/��rB�`��d�1��wv����v
�q�xl��g M�;���>>�s�xQFr���POT���QY*���߱���(�C�'.�}7�����ڂ{﹛��8J:����C�����"1��A�������\���3i]L��G�K�^"�zX���']�`��K[<�=]>ђ0
H��+h�
e���(y�Xms*�͙-ܱac^����wڿ�ܕ<�A��X/��$��	�Lc�j�l#x��<��(�l%��w�a7�k�K�=��h�����~����O}��������	/�)Ï�I�T�������h",����O��~��`]���st�,ԗ/��L$��	l��p��e�a*X������S���6��s�m����M-����J�]�S��5v����t�b�砌h��̊4ܒ0�l�O �Z�U�'��,b-����{���;}�a/D*m"��(�{س��u��T�(���f#�f ���;�<n�61]�bw�����f����&Q�,v�A	�f����=.p�'7S�P�B�lS� ;f Lg&}G�b�^�Ђ/�u�������D�qI�$��5��쒽�1� ƕW��X
����6��F�ل��E��n�_rPp����G5a%�}�[��ַ��� ��o}�[��ַ��a�q�Y�L�L���3��(�&�zv$	@����ZƵf�Xv�|��{���=�@]s��[���<k�;���%|H�J�Kq�n&X�{���>�.�h9��Z���ĩSxΜ9��~����[�ϝ��Y����}�2<��3���	�G'V/xH���uo� ݢ  d�f�)e�O���A��f�;�^��6DC�5eo�>a}��ZA=��ι��ڏ^!�[d�l�X?vq�( &*6�#�K���׌^�5_o�P4c
t���q�/X���c�Vl�Ѱ��X�(�q
��)��p�[�C����)�$Ōj'�:���C5���Lg-k�X�Z	w�RD|MK�k$cA4~L��2���Z-����	D<O_�N%���a�Қ���dR�w��Мʘ5��#��w?�O��j�����qV|�"׳�Lo�LK5ǱF�Q�%O��2�&��s-Xt/+�U}ttL}iV;�gR���Y^�e�ZQ0���\y��46e�b�0��x:�������6�k���v)}	���Y�Y]N�'1ZD������^|�{�1V 3j0�!��@ƙ�nT��`���p��;TR��S�"ɜ���:�N�uP�	��u���<���8)0*r�<��4cF/�[��6���~0��p�n�r=dY�6�:�$S�u���~��i�d�������(�B\���˭�M�uk�����3H���CZg��A$����;�$�Œ�����g�s�:�M3�U�()�:o@Xф�̂a[��YFt��1xӀ4a���|- ��o�^t�J�dpL�V`�à`�ޫ̨�Ͻ1��F��s�@9��N����'`��Q���$�� [d.��b�fi���0�M����'b=\��tM�8�Q�0R{����н��^䦀�1��F=p��Y���{�r��Q�m$��_�z��9��YŴf�����$>����S ~$}�p ?��'�}���N��AdH��@��kL&5P�FHk�{�{	y�>x��0N��0�d	��8<���3hPi� �*���p90����ȇ� �ny�����/B�L���+����!;���mղ�˧� <&:�O�%�$;#�JI�/�]4o�mDL3LNo����0%��k�J���uç54;Y�巽�ݵ_�׿=t�yv��C&���?�5P���^T�����q�CMkA>�(��4��Rn(�+djI�.�J�ϓ�܈ x@��,�_<Ua�lwټ�=�n��?�'��\�dÒ����۔ (�A�_�n�?��*���jW������A5��9�{��4�wZY��
|����zY�"��(v�ɂ�	hP��V:�����Z9,���G�q�nQ�GU]�E�u6�Y8�s��PV�r��Ρ�Y����0H_�F�م\ҧ�}휴�kh�������A��t �c�},F������m�}"�s|�Eܢwf��~�m�������Q=�3g���w�E}���|��������e��@�B�L�0f{�&^����������?}�[��ַ;�� }�[��ַ���owP� ��Ǌ�ڣf�F%�CP5�c,�����
��T���%�Ԃً"Φ*���-�@
Q�9�J�X�Y,|� �:}��Q>q��l#P�Y�s�)�u�ݾ��4#R1�Õ./��R3�9&X(�R9SP���j-���<�r�:�������u��w_�l]��,�7yF�8� �����Z ���&�?{��p��e�|�}0�l��\��X+X��f�8:<���XL�px<)�.nq���:�-�A2�)c%2��BK*@k	���"u:
���ZSY�k 0�::�@�s�:�U+��\�!����j^s8ǲ��s�Ŏ��#̺$�O�k�Yq{G�-gUT.��=����i�f�������Jπ�<��{��ļ6�/�O�>����7o���]6+8�s�(��i~0Y,�{�Q�x�\z�!����$ ��18�?��o�3�l�x'c�G���~��t>3����d�NON��^#g.vz�����b��-S�#��l�>[.	l8I�v|t��"�{B����iW�t�koL�s]�j���p!(��T�;gϐ\_�v5��8t1S,=c��ik{']c������vՀ�7�ʳ�����=q^�@K�����3t��g��+:�tf���H�5�&�c��\#���𧰷�'kQ���i�)�+��3�`���
���J�!@��#����9�?�3�q�߱� 1�"��S&2�
S�=/��2��FӸ+�/ {�`S�`���<I�>�3�Tr���#g���RА|�Ge��p���:P�|�=r�� �t�Xۡ� h���H�^WF���E�t��,7��]�.��B��

V<j�e.��'K��>~>��Vx���@�G��+M���P��  �BQ�M��)7��*.��r��B��vomN��+�A�Od�4��˹�ȟ���%}.��� ]��߅�S�MԠG��3���),�۶H��K��1:\���|�/�B�;P>[gנlRόT���Χ���W�/S��a���O�w�)��B�h�7�_��O�Gb	��@��������p��=�ܚ��, u��W����p�V���&���k��~�lno��6�������;66�t흴O����_i�����>3�/��aks��id�ay���eY;P�!���<�9�%�[]PT�h����a�I���Yk�DZj������z���zĮt�D��r(� x����������y^{�%��V��SOCL�c��)�.20�,�A��>w��Q�U:u�o����΃��G�c�֟}����@�������i�?�#����&݆{S8�
����)ߺF�%��׉8H��f��&*1�_�9*
N��
K�T8�b@��k�sy/��6d~�2�Q7`cw7���=`�]ZfL�<�!�&r��Nv:k�X��Iӵ-�(�B���kjpE���2��';�	V"��"*u�ЎP9TR���,jVw~�q*kN�-+$�ҷҖ,��/�0�'��Mt,X�kѧr����7*�@V�Y�j�2���G-qR��D'�ĎpdGA)�l4�~fDj�ڡcb,���uf�aQM_�})s>�=����&��i/�Ē�t��/D)�S����kB9;�3��}����3��~~�	
RĀ�a�ߙ���/1��ɑ�6Ft{-+u>Y�y�M�Q��|S5'eW!�JQh�zD{��ַ���o} @��ַ���o}�۝�Xü�L�*�ɀRP}`\�Q����(������R�8��%�x�:W`��-�tu��_(]H
�}r����t4Y���2#�<��Ĝ(S|�����5u��� ����~�т�;h��V A]xݺ�y,�CN��  ,[ΈEz�!��%Cw�,��$9ь�������
A�ݝm��܀�d��1�	��?[g�����^hz�bLG�u�O�O�\��|Z.6�GpP3���Vj�s-n��րe���4�y�9f��aͳ*N|�[���
��9(��loY�u�T�����c��?<��*�� �h4��w]���666�<9�Rf4�P_�x��,�)f9mnn����-x��פ\�G8��.Wd{ѝ�<3D��`�2&�yCZ��3g�	��#���~�g`0��Kw�$�;e��!����=���3?�!ؘ���� 
�	��\,���$0���1���[��ǯ� �F�px|���'`8�$c
�bV����ֹ�֦�����sXe����:�`J⪭���L�s��2�pᮋ����R � K�f����1	���
���Gd&@�� 3��in��_J}Ō�%�Q���(A��Q%�YZ�ǃ���瞃_�.��� m�״3P�t�'�:��8�H��H�C�ӌ���g �m��_����1�J���"�#��|���x�%� ;�y�A�'@��%nXJ�Ͼ���{��&��� (�dc���O���{���?N�qـa�;d7��!��J׶�D��E:�h�*��4�^G����1�eq��� ���op�;�]���������+ݖA��>��<� ݊�2ǋA����V���tOW��N�#P�h�;�;'�ҌY��
,E�&zpS�W�������=a})KN��P�i?��&��H�a�/l.�b�j��8FA(~L��<�"P"�0�iX��T��@r���g? �.]b�j%�o
x�D�[X����^5\" pݥ�` �ի����'8����R�zsk����u��|~�T�
���cf�I���d��^@�|�Qһ�s���*���t�k��._�D�b>=�r�1J1��:��rʢX�-�Y0"8�Ud�W&����� �P�J�Q��A9�]�`� ��3y;����v��9x��'a����+�A8އ�|�m�Oa$vhv�SCx]�m�,,�bg+0�`�D��>�~L��E
��]ғ{7����p��o�p�l잁�LΟ���/�V}��璮�Lכ����a0�Mv\M%U��`��-��1�`��m��b6�틻p �)p E�)-F?��u�0L#0^���|���*��I���w���5�P���6�'��]��B1/�����mp�lֻ��4�ʌKQ"1f�^�K�f*����G����//N"�[2F{���n��w���'9�j��b%�E�6��nm�
JY�y?�^��4���^YZ������Qu(�{��L;�����_[�#�E)c��>��IjccK�����!ϗ�+��o���hyN��}��g��iɜ�|��8H��(��`����t��ǂ��iݡ�A��,+Ʈ�ǅLمԖ��N�o{-?ۛA�w��ɕ�}�[��ַ��� ��o}�[��ַ��q�^����P瑀1�<��=� 0?�:��Ѯ��^�J Y �,}�Be��L���p�*]v��s�-i��f{��z6��~I�>�����c�ѵ���d�]'ll\�݃:W3Ǥ��@�x��LZ��_�"���}�CzඕL^<9p��C�Q���;;* X��~��ނ��m���,��������D�K�����������1ghv������u�D�0� �����r���LU֙
[3d�:�ɳ2� FE]��r?��&9ūZj�W������)�я~��}p�=������g`��Yx晧�=?�^�� c���hLuA ��S�Vf�оh����J��T����4�Ho��}{�}��/����2<���p񮻈�7�����
Bx�����5ߝi��9<: ���h��_g,10�ىV���e���3�(3���Y�
�����>���x����O�ƺ�N@3��`�9L�r�K���:�řJ�0gΤ�'�S�c�/'���<��R� ��%� �N-��?��L���k׉u�,/��@ 7�_�Lݚ��`y���\��!]���|Q0K��L�[o�:����V�& ��
H�k*�V�1����54�����4�������H7>�����w�������^C�
h�uE~��T�s��?������k*�y�@���f��/8#`2f�]eB�mK��D�Hs���c�<�e܄��C�C�BZ�����0��*;:D��ّ��^4'?�T(���w��*$���S�E��m��a˝�u������~v�L��=��R�43Q��NN�L�6�h��6�.�0��ݍ��B��Eb��m��^�<��8G85����~�`wOp2:���D�᪫������e#����>S�Z���S�#@�Kx,ʧ��7��;�xhMn�"���	��xF�I�*ۂ��OfS�%�񐂃b����Q	f��i�>�X"�%��U��x>����4�*�y;p���p�ҥS�]a��F	�T���Z��M׵9]7=t*��1�Na^[9��4�-˓k�J��T��@�G�:N�v�����X��?}�S�D�Zd})K����7����V���;���	3 �$�Dq�,���%[NdYr,'9����*��ʏ�b+��X��(�[vYrE�$��D&H� �bx����ϸwwz��羧���ɇ{�9{�ݽz���[�[9�D���R�U2K ���c��)o߄�+0;z ��D8��kK�ψ��ޅz6��Ͻ�մ��,��0�~���ᨁ�˰q�!�Isz��kT%�(S:J�q%rH�@=���H�I�+y��5����O<[�ؒ�ux�Mo^�6�݆ۚ;�${/�m�=8��I�w��߀P/��f�j^��ƻ�k�
�湔9 ٭Ė�C���
��`Ʊ,+��T�*��p�5���2.����R3�k��ܜ^1���>�6��d���U%���=���>̽�eSԑ\1#��v�8;�W�e]��E�y���]B�x��?:E[Oe7��z'Y�T�k ���E)PZ��ل��T��(������6V^IK��}4c�Q
�+vww�����ϒ=y�}����׾7�]Ց�;S}:�`�+s�2��|��ra�"sU�u�k]�ڷK� �ֵ�u�k]�Z��f��Nf�rNjAb��� Ǌ��'841�S�r�>�JAO���ΐ2�A.�p����_�'�P��}~
���V?V]m��\�G��NWǕe�̹3�rG7�w�����0w7�A���A�}׶�:�z����, ıD�L3�)��av� j��Y��uA�5XXX��!�/f�9v�������<d4��ұ��^��հeGapٓ��>��,�����(�O
u���?��8q�a�L"���0-�"㜼(5wWǙ�>����N�<	�ߧS8z�8;z>�t�+
��f�oo�9�C��
��c��鋽@h����s�	O��Ї���KD���/}����/!L����(|���ݽ]8u��p�LS���,�y� K��#���n9���hl�� ŉkU�������S�����5q1s��ݣ�x�GCz˓���cǑj��ׯ^�����$���rX�qq�j03xv�WR���ZXQ��e6C�yX��e�)eCT&E�D����r�� r-���hD�_�Qs&-S�3}>�v�ic���=:�A�	�a_���1
(�1@��d2eǹL�h8���-gޣ3z<S����6�S`y�`!,��8gs�X�bn9�@�E8��QBD�>o��_��4n4O�,X9$YjZ���@kG�tK���	��4?䡁�uѼ;e�a>c`���Y�=ҁQqt�Db���@��c���,c^���H���zPP�Bt�Q5O��A��`��I��|~�_��׏WNd� 3�( ��:�2)��2håM
 L(���or��Cݫ���n����/xr��( �%��lJ2X�G(�X����{R��gA��t,�A?azY�[�$RlK:�
��<��rळ�ʶ�R�Z��P��Q�7J��a��/}��I��p��8y�����_�3o������E@��w�,x��z�����q4S��&��'��V�o��<������I��u�ܺu��;	�àX\�/�i��&=��>@k���}<��sf�&��y��	�Ɋ�rE�Ѷ�|fu���l/�ѣ3iH�t�`���[b&rĎ�l�+y�@�3J���<���(�e���i�����H��j(K{q�0L�F������k��{��I���l�b�d6X��f�Oc�@}>H��Qp���x|ڟn_�GO�Ť'�������to���,&�8Ϩ̎O��{�Yp{W b�[�ؾفe���y���t���y�����qpXZ�5?����k��^�~���$�BF^����dB�W����ˉ�'���W`����[�|�M*-��d���b�� ��H�5>D�+��P
E��3�b��d��AT�|w�X����߀�g�w)š�4I�e.��H�elqb����<��
�731�C�em�bxIi�k�Ӂ� �n�&�Z폎K~)���A4���V�"��V�&�C���`�,�N,�4R��/��1j�+M�)���3[If���xޫ�)����{���'�5�'��I���͛��oӳ^<6-ㆋ��M���e�b��_��\y/�[-��@jV�B��b�š65]�Z׺ֵ�}� �ֵ�u�k]�Z��f3@^왂�tv�{+2}��l4�e��8�x���%�3����S�o?�?X�I������v����+�� vq��O����&W��h ��fdr�'漗>���o�c��\RZx�;��d�u^<T~ �ʔ���Ϙea�Ѧ�ڗ��^Er�./q���{��ߣ��Hx&Ri�#Ѕ5�1���*;��Y�S��^�뮬�Ã���xu��e0F���@#�cv�$l3�?e2�L�ʹ�� �:
 ��d5�m%���w��<y�u�;b@p��F}:��f��0VؼE/��"�Ts�eK�g��w�l��ځC��S�Vp��Q8r�<3�3�6������t"ˬ:����^Ȓz3��z���ç���̙��k���)3�_�*�������&�Ko؀�]:種�IP�k��ǬBoN�h�ӪbP3�1����㚀^��F`��Kcs�d3����7��[o�%��揆�4��qp#=���3��w��}�~k�-X]]��䣒@")@����Q�}�1N��6>l�l��P>t���pA��&Pn���LOt(�g����t��Lq��lJ�8�,s�B��#bkh�!��RX��+��0��g���©{�!�����ھv�1(����k���M
����8��ԇ/}陴�{�K��K��@)�|O�z[���g�k9��='���^��A�7�k��?�3�5?~�����$�0�3c�2:�yx
�\ց�BF�=ؼynoކ�7n��!`�z�A0�'��#��#D�ں�V��!��tͤݨv4ǉ9���9�1�r���,�XcXk���.��A��w���'.���|�F�دxA� �\�R`8�tl��#��fwa��u�a�h�������%Р�M@؞"��=W@���Nm��l\ e"@��H&�W�x���/*ѹ$�t\-��|噙�Av"�M�Yc�=&d�`��:Tu���Ʀc��tk�����4�7�
�Ӟ� ���jy�)ұ� ?X��W��?'�pI�:��{�я�]�0'p�"띐tPy�i�/;�=�>��ԧi���_�����ӏ>ˋ��CÍ�7��߂뫔=����Ξ;Oϳ=����~<�[����{�)������i-���O��Ko�W����
�v����0ĂN�6�J[,l.�#H���r���w'XW ���m������s�;�L��j ���z+�~o/���奫p�ŗ��{�F�ݴ�B�u�����	���ڔn?J2�t2�0�݁GO��܀{:
~��+�ɮ� �L��i�v����h�a`���8�z�X2��t}!}�Ai��C,Q�dc�� �[߀��Y����I�I���)�O%�֖`���m#��2,.�#uoGd6s��s��p�qr�Ɨa�7�I���'�����$J���G�fo�a���M�3�q̰��H׊���d�"2`��z�ԍW�>���>N$We�Cn���8�	P � z�q��.�k:��L��V'�k���&�m�^�&�Pok�XWD�K۾�wfP���� �����{�(ayV�g��3��"�L����~y�o#�qB���T��2���Y3��E}��L6�ۏ7+c\�{N��R���f��ޣ�E��� �9PXنh?C{�(]�u)!���d�S�Qq�+yψ�.��@��ɻ,9����-�Mf��wN��Hg6]@׺ֵ�}�. �k]�Z׺ֵ�u���\oP9~ɏ�k2 �N�e��ޛ���=;���ggO�t�� s+8 �Z�$�);d�If���QZ*D�A�YV:^�1�_����[����
N�?�e���O�5�E��lq
��9�>P�@(�F��+)�A�+���CK/� !W�cjP{8u��T�uks��3p�9�L��и�M��Y9�Y���� �O�p��	��X�lq�a��NY�Q��J?(����-�}@z`@g��-f�ϐb)��{�Sق�XJ�^�U���Np���D�����(Pg���#@��c��@ק,u� �N��RV;�p,������l(c�{�9M����$�v���HY�-15�s���Y�Vz0���(TpR��hKჼv8H��օ�E�F0�i��bvx�GI�l���$#8th.]�D2���R��{�߃�dB�#�<��	���:{��q�q���u���Q�����>|�0e(^C*��ex���{�E�p��=b���X��b�3��O��cM{d* z~�z��=�.穱�:����8���N����x!+�
J���Abai�9;�JȜ�zßKVG9J0�Hy��gc	Խhy	�bE�<}��݁Ci͢��L��u�\�r>���7���μ'�������?�<��s���x���A��z|7�% �Gg<et�Y�Ƥ���%F�%�$&���_�+ǮH��
�{�d�;P�
'��(�pН���di��8Ec���i�ƴ����b�k�~+�������?�1A&R���HV6^�脁�����?��HkO��N�7?�� s{�R���g]�e�K�H�1�Os`�Sh�Ǿ����`�)0�te[���I]��sp9c�t�f�h h �M���ǂ@��"�4��h� �~���9�sA��L D�Bζ�=U�&ơB�Sf�jw�ر����`�R9OyRM����� 2:�ϥ��s`��=��_�Z�^j( L a�U�	6�`a)�6�?�AI���4�v`�Ɉ�5C{gI�M�C8y�}�օ+�湷������s8�t�מ�|�駓~]�,�CI_<���gI�PG?��;᳟�<<�Ѓp��ͤG�
/^�&��_z����~/L�.�"eG�1Dl��(#bsl[��Fs`���L�$�L<��IK��}��M
�1������b!:���"`�L2蝕��O��c�NN��go� `@�ҩ�����{p������>|ey�d�e�6|�A���p._:�}�4^���<�4x�5�\!���s1�K5��4��ǳ1��&p��*�f�.훸�am��o��=�`<&��d���{���#���8Is���o«o\�[���wC d?=����	í-���xw������U8p�(�$kd�}j�l����m�G8|�	����Y���7F3x�'�~͖������{|�J�*� �����u4�;�T_�7H�lya�Q�PN���	�A���&,�Z���s�N��v�w�lEc�.P�w'���(����84倽�Ne����95(�K�1Dk��	��`�<����]�H�%)�KFٽbQ����Z��DG	Fv`�l8H��}�6�x2eۄ�u������� >�SU��I�m�`���r��s��1���V�G�ق�B�� �Z��߅���ȥrX��0�`8*���L�W�TԠ~��]	��v=�;]�Z׺ֵ�� �ֵ�u�k]�Z��f��z�2uK�Y���ya�O�p2��Qj
:�<0>Aj���g5'H�9s�X ��?�|> ��w%@�}%BORd]��B��}���v��P���_�-���<�B��pPȷ#`-�׋��)ffTǳ��F��bW;r��a<�@a���dx2�M�LgP�^���DM���o�9�SC@?L���Z��	�SS"p�ٛ��$��R���(���a�Yt
#7RyO�Bg��_��P|�F@��#Yd��iA �6{"%WW�P1)𑮊�R)�O�T�wʟ��( ����!�����iJWӼ��0���7t��RG=���6D�q9a�]-���Sf�(���Zg,+������yj�S���tݥ��:u���g��K�.�G?�A�z�*�ƻ��+���`	����aeu���ik{��"HZ��z[�dSp>g�d«h�X?�{���$���W���ӧ����0�:�n
D)O}N��5C�y�&;ߑ.�� ��g?���p��40���I8S�,�9p�Pv���@4l�d��u0'5�� �7��q�$��G����K��9��yL�YWD�^�5�� ���
�dFz��"�1`6��a��&Ѡ�g�kk�:0����~�~��4����8�Ar��` 5(������;����:�uͪU�4F��������fA�lN�ͽ|����>���?��t8.���c&��T�t��,;$�m���s�t"�1�������(Ha���K�P?���|�
l!s��=�D"S���	�?�,��8ݛ5Z״:�	 ЌSrt���O0e0����1h��f��fX
��V)�%� ��jS	 �A�]����f�A	e`Q���l,dZE��@�A����S�ڕ���?j�h���>�n�O��܉e�7�=�-��.�-�D;T��؃��/�}a r��S4P̮-�l?�9פ�ę�\ub
ד^���P��g��AH��>�����VZ�I>˫�ՠ�Orӯ��AD���W.�0���h�x�4��v�{p(���vړ��������R���{N�8
g_�V���_�H2��2���o�����H��j�#?IY$5Y�9�Zǧ�8eG��B�������/#4tPi��u9���	��Q��ȁ1*��o�����[J�p#��=�! ���M�^<p6N.����׾
�z����&3j�,�)�N�������߄�3��0�v���O $}��`��E��_q��P42 H�G
�M����I�����3�֡�D��kBk�/�i���֖q?Js�:��z��w��(���=x��5�����	,�����l ]	1R��օ�T.�N{b���R��G�\�ށY�gf��W6��F��4���dQBK��C��[2}��u-FD]W������� �̬"�i;�s���]a/iL�ć�����ky�zg�R�*�2���Ȏ@v��-�k:�*|=��qa�����k�6�w��Ɣ�8�7�]_E��m�A/��L��g+�R� �Q�눮�}����UP~$�A\=hk	&Hz�I}�b���d_,Q`)3fa�#���2E�f��3<,--���5́M���K�ͥj%j����=XӠ �\�_�Ke�jc(�E\� V2#��ͽ��:�k���ʾ�_9E�=�1��n�]׺ֵ�u��ܺ ��u�k]�Z׺ֵ�Qs��zWi:�� p���+� �_���f���c`4;=�{�Z!���U���F��x\�Z�ti��R���Cɜ�Q�\v�B��](��١���@#(��s�V�(3�wߟ� ��_P+��:�ü��I�
��Ubv�V���^@F ��Mx��o��cG`mm�j�s��,�+��:�6�QmdOԘ9}��A8|�������8�L�A`ee����ll(�̉��"@�����٥L�ݽ�k[;;��d��1�  ���T2�k�\����1�yԥ̠�r�a����
��Q��iZ)�3ЖAu��Czdv��gW�;rF6p��%�?��8@T�����2�=9N�\��~.�2%O$�ωF^����Pyz[ȶ����RS$+=��BZ3 ���^��۷�C�8x� |�O�����.�uV���駟�'���[4��W��*�������G����Dێ(u�lI�_��ހ�ﷷ�ags��?��OG�D��=�|J��v�
1J >2КAP��%2���85GiT�Pv;;�/^�7oܢ��g��OءLL��Y���A2����TԼ��G0)�q��l7.	�Q6���:\�{�??��?���e�ͽ ���6f[b`������#�ǠׇY��7/�cY������{�Y����m�*����C��eM��z�^�bd}��u��(ˋ�xO���$�Q_P̈T�=Ҹm�v�_����� �$O���x�=Fl8~�Ν#ݨ�56�rG�!�2 ���\���8��&"��B2Ю2a���1�c��t�$��N�SY\o,Ӵ̺Bz\;" �b��c�`	�$�{	��ڐU��}E�_�`���(2�m��"�)�3W��h �fӗ`�R"-zk/ы^���/�_�Y�1Scg`/���{��)wCT���ʫ..�(�|o-�@����A�<���0�u��{����[CXX�S@��!�Û�;p��9�ݾ�d;$�8� �)ܺq���W�>��
W�.�#v�QM�7���Ef�`<ʎ��7��J}z�e��!
6A��̆����kX�c
���n�\,����̍��
 ��ⷒA\m�"}?J*6H9�}sy���lY>f�4�~�T���";o��� ���4�5��k�t����K}�y��Y��p��E|z�u�؋�����w�*�vnA/�-�]���NA�!#R�4{�_������G�l!��K{�,�i^0r�Ah���T��!�`4��}oee�XjP�sX���^2P�����/����M�g��%l �pt}����ɆH2��w��i��4.U� ��'��U4Q��t��Ձ��[��J�N�݃�.몼�J;^�P$��L;۲J;��ô�>��7T����21�N��c�`�Ɛ���l�JJ�E��@ʪ�,J-���~P��V˕Q�^%�v"��'����A"�K��@�q��6771=�Y�/�H�{���u�vs.�TY@2����v4���P0C��%�AƁ�7_�ָoY�T~�x��Ʀ�1�	�9b��d��fX�(�3	��]��^�A�͌�^-τG�lc�~�咔9
�����1�iFބ@�ۙ.+6*�3y��������� T���x�;E����4��gNl�J�����J�z��@iQ���u�k]�ڷU� �ֵ�u�k]�Z��F��1.Pmך!rNe��(��c2H�)A����[%2�ֲ��U�Ȯ��j'�)耨�dӈ��;�����o� F����/�IF�8C4��ྀe������o^2�5���Ҍ���YG��$ ��x��:����ݎ�u�a8j��7/P������kp�����"Q^b49���2ϑ:����p��q:faa��S�*,�d��׮_c�o��I�����-����vw�`k{�7w`8��g��po�)�	A�:6�]�y��A�X����ќ�^�\��3ZkF_H�BZ�Q+�F��\\K��DˮrUN� [��5l��$�~�_����"G1�%`�46��%셁��U��loot���0{0��d.;�L�W����L��|��a8xp�2Ա�*��i�_�[�ȣ��O<	��~6��������p��-8{�M�u�&��� �!�}@o��*:X���]�����?��$9|������_}� �tꮬ��×�jQ~b-�-��������$ڣ|a�/k.��V���~�I�6�J��:�����0|�%��9�(�z�Y*$�/}�������Y~*goeS�ǆ�����P6�F��+/���7(�L[ ��7��s���m'�~��ɖ� ���t-����� �$�A�9�g������B��n�xI��h�,�<A}����yp�;��L��R���]F�L��$+؟�����(�\�3�&���p,��Є��XNđ�,%�n`�P�=ewP������A�VД�oe��a�%[Z��o�����$#���������Fi��Z�+�LDfsA{��)Y�R^��\u�WH��xh ��i�ĊY'GWfYKf8͑3(��.�E�
Pۂ꽸V~�Xl�1���%w�������L�y�!W�� ��k��`�Y[�,"���I��2<��y߄�7�����K/+Ho����]�y�\O�n޼���f0�
����˔Y��X��MY��I��Y��7b��1��hT�x�����˶���K���Y!|�h��'�+�
E�t>>�)e���v)�*�,K�m� ߎ�c�$����4�$��p�Գ@d��1K���n	f��͉�p=S����i{Y9r�z1us!=��Ǝ�dV!��#��fWބ8|�n\�(+X=pv7w��I:�d3�=_Q�f�oh��R(m3��W/@���=%ig���iD�#�8� ���&�d��O�*�9=�ݸF���B/�1��بHV'�#�}��:�N���$SA{5U&w�i�Wsp,�)��B�J�ίb�g��O�]a�ހ��1H�m�U׍դ���Wd9�Q���.��l�ZD�+�Tg���喼f��%/�@����I�g��^ž�Y4��5�w߽����������<ȼ@�E:����G�W���'�")�1O��ŋ��}^|�ds�-��
�;��9�����>q�P_0X�2I�lmÍ��a;�m{{�l��G��Y��i@�	Μ>3e��~x?$[�f����[{{��S�Ƥ��	p ��Y281@K��{
Q����]�`!�~hC6��Z.�$�H.j�������@K���D)1�e��lA� �r='2B���qhD��[��.���ۮS��w�@��,�#wٽ�ֵ�u�ko�� t�k]�Z׺ֵ���Z����3׶3LҢ�һ~]�ه���\��l3q �qm���)F���s�+T�(P��U+-3esG��f�������dGOk5[��[��!K��P�s�3PA N���.�@ג���^�ˎ�9:g@�z�����0@R�+Р�����Nr���(��|s�:v��Q�:��<���1x�����3���Lf������؀�ۻ4�|��cB5�%�.F�ʙ=���P�a����E�M��o�Jt}ʸVvk��A��� ��,c������2�� D��ݞ,��%�T�Ln���l+ύ���W7����.R����l�3.�^�xN\^�Z��8-��G����;�n���Wa�2�[�&���O�	�0��'�Dv6����P�:����\Kφ�\tƢsg}eu{�4�Mǹ�/���G�֭Mx�o��K��/���w~�S���}�$�퍉f3F���f�ܡ��!'����x�~M�\���"Ae`_K�Z�M&<ͦc����.@5��:�@dR�~Kz�X�!�J��I?�WeNk�qL��ξ[�~]�����D��^��~����9�ж�,g
��%�@�
<Ė���>��������R:!�9�Y��~��p]��,B/}>kY���Obq��xrK�a*D����X^��rfrE�����&��@��ޠ�L=t���Ī��7ᬿ�n�꼒.�r�켥(x����F%N�@{��D�6E��5��7"3�> R�$
��8#4	�\����b9�{��"z� ���H1��M�AK����w��ˢm1���9P�Z�����m
;�Fv8't⚍X�D	�iC����'��AX��ಸ�@� ��K�`0�(�=^nC9�$���|7�큶��	�}�Z�"B���s)��9c4�U�3QNQAjGs��;�
�6��4B��*�hM����4��"�<ȿ��Agv�h��y�/"ļ����};*0����f�*�HÞ��G^M���<8��=���x��O���1� �)�P��������JJ�w���_��S���(PF[x��^2nf�eʲ�*xY���=[�Y�`6�\v��ֆb�$H����&���>��Vb�o� �|[��m��y�S�ֺ��}��hr#,A��1�$��^<=WE��-��X�-�A�d��մi;�	T��d�c6�`.]~!}6%և���{�9D��&����/(�\(�gĶÁ W�\���(�d�++�2J���\j��wue9}���� V�V�����QO��t:�w��?��{�t|�Ir@}����cE	3Z�.��
�z�T� �f+oh�mʬ�=���)�!�)��i�2�В`
��<��5��W<D�s){���x�����~���2Rp`��Q%&^�Q��T����?Hz��p��p���S%H��J3�b ����]�?�c�{�.�����Ϝ���� L��}�#�����H���퍐5�� ���4??��?�?����~�Í��l�&��d�"p<�8�K?���O�X][�{�ߵz��J� ���/��ux�����3g�~<��a�~��w\&���S���{��?��kP�H�[zi�����'ɿGr����(�}Jp����=���^$٠�0c�lav������;��Wy�D���u¦@��`�vT�z��o��J3�߭�I����h� r�vg~}G��������:���~� �ֵ�u�۠u ]�Z׺ֵ�u�ko�V��=p`c���=J��S�]�&E�n�x��D�����lFXg Ԓ�ԩ�Z��^�纊=rZ`m_�H>y �a׆`�!��y ԓ"ٸt��EV9j$�j��N�ĴsI3,~t(rf�X���N����'5�:�imHq���ˈ~�n����=��E�h�#��)0�Є�*�l��U��p�-���c4�B�N��\y/v���Z�6�O4؁�F��� T�, t��ABu����0�Jm��{;���c�ǂ2�̠	���9cI��s-��K���y�oR�^g9��{���	$1����M�9���?D�!����$�@c.+�k	��N't�6��S����a[S<F�,ٜ%�E/2@٤����[p��ex��������SǓ̜���M
@�أ�NP��ŋ����K0�1����3	��Y��!Huft���W��eS���r��y�����̶3��R�?e0gp��RЄ�^�_:HNh_��"\������n��B/�k�檒��$�Ӗ���/��2#�79L[ = t�	�	K�#TK0S�d4�C��(��QpS�b����ť$9i�{�^�=i>���J^;�!�m��Ȇfm�z�+����P-hG%B*? d���)��F��&��U��q��h�0@ܧ�t�p���E~Bq�R�;Z5VYW�=���Gy= ��<��'�̬��(�B�H�账�@�`��e���;�}t4�P�ǜ1�V�[3 ���a��U��30P��F�%�쀞�/F٘͌��F�����L$f�(���5S�3X֍y��L?msX�O�@=�z��jEAIЁe2�&s�}��l@�e��}��fF]�I	�1¬�b�l��0����~����F߀�|\93�!�8�l�3'���}"����/Hy��7nȹ^t�����.�C�Ī��k�>pj� �X|n.����,���� �HZ_2��ѽ(TȚv�9���p+A����2��DQ���<�G�\?z�0S8-E |W��n=-���\/b1�P؏����K�����Z��l�,�'p)[�8x�Si�Qj��# r٧�7( f�=���B |�c���u  5�>��;�6j�VB�ƍkRj@�a4�S����Q���u�TʙY�"`���3@����/nA�[�a�n2��c�A�?=g���#���qv,c44�����E`I	�nބ.��F8�Q��@)��_��z�(B��닎@F�[vt�t���C?����c��t��OB?��Ͽ ����]mG>Vn�x�<S�c��p���}��g>��������i�?������ɶ�@�,5��q��r�Ճ��������W~���K/�x����?�S?	x�)b�Lg���3�4o�^2�>8	�|�]�w>�N�v�����|���А���F�eLA�">+�y|�D� ���\�яr�qK�bg��qh:XOE
Z�3b>�e��Hl� �?"L��TV2
����4y�,��@�C�`v}�	*^,��1���z�*�)���u�{}ߡ�$�_�й�u�k]�ڷS� �ֵ�u�k]�Z��>-�������'�I�򽱯��o]��{�B��Y�yO=���d<�j�Mm Bv�;�^�����������vP��Q�u�|3k0�ʡ3$;�
m����s���8g��{��7P=���W}*ڜ����A����D#�A� ��o΂sc5wL��>?������Ҳ�����GHMi�U#50A�/��X���k��:��F��Ռb'����y���J��ݛD
�@��(�/�aNu**�K�N?py���[iQ���2�F�+;�C1��݌�8	�`p�/���d��ak�^�7:���͙o
�KFn��ɧ�\8�#wp�����3�©S��T�����1`@koO�3���f@O�W��&t}���s��3J):��L��d��q�}{�����^z�;
'Ng�����s_{���a{{>��S�ճo�	;�{2,3�`���Mu��IJY��j��#`,ӗW6�L=�2��I��-?��ϩ��(��0[-����eR����Z����*v�2��R�DeY�
&D	f	Pc�~��*���|��B@d��R��/(�^ ���%vJWZ׳�7��>���<���H�ƅ ���+PO*�s%PE���ZQ�b�����<�ܱ���2w���ʛ\�C��HM]^<Q��R�e�)�ey%cz��Oә�q�` -J S�lq���^��]׵�e��g+,��+ P�.����P8����:7:n����2��oQe :����r(`���@�
H�Υ��L����Gc�>�B�7�x
a&9�eX��^@�>OJl`k��e l=�ǋKK4�x_ʆL�S�HR:e*��3*3�O\�T��j�0�������܅��ґ)r�
]>7)y��e[���@/�|���g y��<��b%�ICϡ�"�4T{:2hN�M�:�s�b���Q�9�໕`@�%%+U���\hy��젨���x��; �`������n`
�i���o��H)�v,g0[2���D�=Z��b���������ջ(�}�}�lc��2�T�<p}d�#���>F˶��Q���i�UQ�����f�1�g7��?	��,/,yXZ����x�	�W��.s�A�(�jo�5gi�ݸq��O�Lُ�Sf��	�m)x8�i?ZZ$F�@c�J�2�P�g��g_��_|���= Cd��}�5d�I?k��~��Ju.�Q�L�<в���j�d&���B?E{�2PG���3���_��$�"��)I�?3ӨL����z��A��0�o:��N��3+��"s��"+j�"�������0h���f�:�#ɖ��'?�ɔ�>�������x��o�p8�����/|��>
˫hg\�������k����ܸ�t)��$y@��x����)�ތ��H�D����g�$c3����tL�}��O������?�#b CY'Ʀ��7��1�;X��
f�����?u5��vr�3��f�	6=]'���0R�	�l}�*�Ak�mV꼒=k��.�Q�^�f���+K��	J5��|�е�u�k]�vi] @׺ֵ�u�k]��ۧE������_8?�6faV���]�`<�8\�ǐ�i�X9�۶�G�Ѣ����~�k�[�+!�~�#�A�L�j0-�����u�n?��������ݾ}��t�b}����A���U>����j�4�V9���'!ԌB����N=%�Q66��@һX8\ ;I��/0�j���Ns �iu�*pT:�As���]v�� �'��K(�N9�!�Â�gt�W�W��W�4Hv�k��c7f��2Q|o30�B%�U�ɝ5��! vh9(��J�!�O�����@�g�k`�kz�9_u�+�A�Vs�Ѕ�
H ;��o��r�\�<qvx��E��RD�Ҝ�%�H]��Ex���w}�w�>f���[��J"�1���嬝�5�y<���P�8(�2�Yc�c0ֳ?u�$|����|�Cp��%)�T������ �|�[�����i~nܺ���
�4�2-��@�+�k��{�u��TG� k.@r-s�ّ!j���E��AF��3�7^�P#S�������s�@5*��UM*(Ç�����4o-�VS����:W����%v	���I<���s�����:��i�1����<<���;y�$1E�![e�JM�2n�8��l%�(���ig��b?�&�z�t��bfZ��G���  ���{Vт=l>d��Xݡ��ގa��� A׫b;���i��y�ϣ䲖���8+:�^B�(�4;������e��E��v܇D�AG��x,� ����6�N ��?�{�<��r�{��e!��9�z^�dE�NwH� D�ק�|
|H�������W�&{ �'J}b�lQA��L�1�H��iA�(����
�w9�"`�u �`P��8��f��GLu��88)qa ���{�	�I�f�k8�A����8����.��k��8w_�-�$��pa´cAb ��A���X�U�^t�`GW<�Zj#(]��9;��x��׋�Z+���ޓ�s�s���.�5P��8��U ����oݣ- Po����V���Z���dQw�l:*�y%f[U:K{��8вz,?�W�{0���Ȯa����(��[#�jdJ�<������7����}�QI�0��$� ��+nIf��n%h���)�f;��~�����$�b6 �ڦ'��G�'`��S�./��s��z�v�98Ц�}���)�ǩ������@�����.�7jk����y��gy_P�3{�鎽O�����|��k;<O(Lo
X�ӣ2`		d�9 �f�����>"��dk��ګ@)k�Ί9 �v�4��#S�l��<���������TXRB�A�����w��o�j�5��y�������������t>v�g�������F������g���Pi��dG����;��w�/�{����C0M2��%�ٔ��'��v�v(�B���>��6�1�b}��>�[���-�D�A:��Z����v����R;��+�ʩ�s1����D��$^�U#Qօ����JG�t  ��IDAT�ӇYl��Z	��J���[��е�u�k]�vk] @׺ֵ�u�k]��۠!�/���w����x���R���h�Gz,~�5(Ʌf-��Uh��Y�޾v�����ǣ���� Ot��0��/T��W���k����;�--�}���2��^8n���r��^>���}r<kO����_/��:�Z�<��C'-=�K���}�>��Y�.{nā�Y����~7��F���c_s��
N`��Jp����oqܔ���u�����C���r�5`#�,Ea�WEs'c���\]�f�|�c'��/h�_<;��E1�s���=���QK5�i����~�zPH�N,"�9b<�fGlv���ʦ��Sw�M:�^j#�I`�,,�K���ǋ*u��&7ţ2��Lb�)|�N[����|Ξ=��CG��#�aqq1}�P���_x����N62�_6=�Y��٭�;ƥ�� q�#��C>�C� x�!��@�#z��z��~��¹�o�o��p��u�F���=;�3�u�k*x����՟�f6���3�2�HYe���b��
3�+/Y�<o�V`5�c���?s��@�"�=�'O���o@R4?����y������Nl(�~<�Ҍ*�՞M2�.�b
X�:�4;L��&��2{�1a+���DXfM��w��{NQ�\l(C-�m�	|�Q��AS�[�gփ�i��M.k��_���A`����|?~zi|0��Ǌ�3�ۼFh*�ѹ��1"�Yw�z��q��DHP`]�Ja�I�9��l9�:P�.q�:�u}ʊ-����V�k@�sH�#�&<���` �fij�=`.8��+�����]�u�1����E���^A#ä�D�_d1V��`0�G0d܌������B�_�5e�F	6�s�3]޴�r9��ƚ�i({x^(`M�]Y�Id0(�a`u}��0J4���* ���t�b�	)ck�=�>��/憏���>��Oߒ��b��L��E���J݈�6�YVtHy{�"����Vm~T�����,��5t���Gy��܂b�)�WF�% �<X�WD�z���`�/:A�d�M��4X`�͉�� �V��r��sY�=��<e+�8�Y�t-9`=�D������#	�%{��g� ��tVg���:��U��w��G��hg� 獵%X�Wp߽���U2��p�iҾ���*f�:�@@�(P�f6J�`�w-k�%��q����.�0���q��ĀK{��v`ewn��E8��������������J�0�cV0"��ҩ���bV�¾+�#S$2g�� ���Ӹ��i�#A&3 r� >�N��̼4L͎Ā[-w����,@Ї+W�p�b�O��EA�������%f(h88hyyN?�(�&�K���/�_���N�`��hw����|����O|�|�{����e����sgi��9
��"�iK6�����3�z�HJ���׮��/���;�����;��x���yP�]݇G}���3iM�yL��-�;l��Xx�Ә�#JPX��T;ۯ��h��Ȑ������~U�� �=��o.�E���u�o��w��fcfq�[G;Sü�Fb������(X�m�
������ֵ�u�ko�� t�k]�Z׺ֵ��M�c>���z���|�8�n/�^~�_\__�������wC۞���q����E�Ze@��ˢ�-:d�=?������`��[P�8�ǟ~��?�ȃ�d�ȳ�~��������6�vc�ľC�U�\Z�=g�eM�wRS��L��C>��lS�hـ Ns�)�S���[fw,ρ�Ѥ�  @�w�[�8$�#?g��r-G��b~nK��{8q3*UpK���� �,�Xc�	J��2�}�u��N8��K'��[�LK(�69/S;�]v�@�l��n�iʙ�*A��]u\�)�PF)���ε���VJ3�5�lq�׏<9�Q\��x>�����;�TY*B��Is��P7�߀��[p����q���gΞe �@.�Tr��{�o-X�[[۔���u8w�<����/�������xHA���X?=='����t#G��B)�uf�0z`	D'v��4�>� ���>vjG��U�	g�"��h0G~�BlΨv���l�-�@��7/PH���`N�~�j���m�4Q�G����0����Ԓ0�� �q_��.��*Y/��nz$���<��c�����DznJ!�P�l���r(���T|-�9
�ޤ���:���=��L�t�d"ࠣ�<����A4��C?/�-���齝�%�W�Q�'�e�h�c�yߨ�@N�fZ�B_ȽH��LM��(�%@0(��y�黀~qN"�aA�@{��Tzj$#������@c�񭠕ʑ~gl*8~XA�$�5�p��9fC���;D	���鞎�&�D�4G�^#�H@�ԙ�`9�F���\`�W���sf���)]��9�u���f<�{	�,����r1J7OA��U�a�t�26 �}"�o���M��\�(4��N�כ;U%:*H�'5�$�L��2akxnq��e��Y�B�G���e@*곺�)Z�:�Nd��HC���YT���ǜ�!]������A+&��n��r�r��P�C�a��}8
(g r��vz��
#�8RW�b\�ԗ��ਃd�o�ud0ٓm!��T�gG�7���d����S�g�;pd0��}�Q��Up�'�
#��~Z���-v�Z����qh(���_��Z�O۶ƺ�5ᑂg���0�dW�U*s@�]�/--gWy/'��7d�*�K6@�Ma���~r#���'��=�v�A��IπA>�6�Cگ#��^晙`�,su�}g4$�(� �CXt�u6��s����-��f�SI-�/������Q��?J�!�� `L'�f�AĘ��y�
f��������x� #�!3�>��;e��uzI��VVaiq	�v�%p/���)�w4�Y�U� �~;��?��_�'��N���I���'>�C����?�^����H��X ��g��.�=�
� �� >���k��+��cX]_����c'O���<�ē��瞧 H� ��X�b� YN��Zs�.��Eh6�b�)k�"�5m_�������K���� ��I�W%��!s��{��РiaRiY�i0gRRM%���1?�L.R��8���R�!Y]�Z׺ֵ�s� �ֵ�u�k]�Z�ޞ-����wm�x"�˗G�^����µA��jf0�U��؍��&h������s���o�^o��_@=�S��ߝ���?�ї���8��~��_��sze����ht�׋��=�&9C�1�i��{h28m�q�(�Y��W[�X�9���4�Ĝ~n�<�y�5x78-�m�%��i9���'�s�x('`p:n��Tp!s(U���Z����1���
�s�eqS	��.q-� `��7J�)L"A�O� ;����Κ���� أ �cw8�u�d��G�}�Hut%[�c��=�.e����R�d���̕:/餣9Qٹ�AHQ6����f�o�@��H��z�[���xD`�|V���ss�|)�1�y�1�>��D��`woLk����M8����A��
�`G�3��p�U��2Gz�u.��c�@���
��hV 3�����?����'Je�dU�D��g�4�6o#u����YtU�*��<j��dR+}�uI:Qzx炐�XY�H#R�Nޠl(�eȢU30U�CY�=rt��)�.3�ρ�P��N1eFu��jG4QΠ�Q�
]#��p\!69;Ms��E�`��̓+FCwYx��8��0�4�^r ɚ>-Մ�6�+�>�!��x|+:�h�U���h���fA����u�������`���	`��b��2c	�:�ԯ��e�K���%U_�b�c+Xh\���A����y�&a�h��Ce\!� ���%hJ!
����f���X�DǄuq�]��*a@v2{�� ��ͭ�YM�=����V���Ds@�a�� 6V��r�����@>/�q�w*��ڕU��+���O�Z�Y���jI�Qޗ�"_��  �p���l�E:~x\��	d��s��G!�*ŵ�G(�AR҂�(��w:���6����� S��̓��t&�8"�"xm"̶���x�#l�o�T��X��}�l.Wɾ�0��cݪ�5�d\A,�Sa@�~c��S���Ë��nry�)�;�`!�\?U�t(K���,s�镲����}~7�h��$a� �]�1��yiq��;t� ��#�ӱE�����IO��>�qx�W�K`{�	�Wn�+�}�{��`��;`����vC:�F��
&[.��Z��F�p�<v��Zk� �=�����<�&3w�O������v�B��L�%0 ��Ը1��A-��x8� _�牒�D�{x��,�^�P��d��% �rY�w�dk�������]����$W�ԷY~Ǒ.����Ĥs���o�?������*<��㰸��
��Z����� R�&��0 �˔�h�MG���5l޾��~)]�1�̏�쌧��� T���E(�,�=۷��O4`3�{��%�a��Q�A��r��J�-�5��K��A�=Ü��~��._��C��A
]����v4�^���(Z�K0� ���Z׺ֵ�};�. �k]�Z׺ֵ�u�m֜���zcWT��.���{7{uǁ�KM� �0ĳ�G�C?9��7��`���z�z{}}}�;��J���Wׯ_?������O������_���g�!O����
b�B6 ����1��ٖ�8��C�9��,sK�1%��ot�6�q�2�֜Iwq�ѳ�V6d�߼�ʴ�s�ϻ�3���UvvBsv�#'H�5O��%�oQ���@#�.�z`s���3Ѐ���Eơ�㜁w�ۗ��9X���@�SȊ�|�� 
�hT��p�s�f0�����5R�Gc������3l��J�ǴE9?�3|	P-N.���qF#�/0���m�[ɤ�9�L�0���& Zn����2$n'��N��| �y����p��M�ۛ$�B3�`H�!��A�Ʒ���s��z�tmO��3u$H���q�4��d�:	8���Ү��M�'�$ ��|>I��f�M���A��T��+Y�2�JA��!��r�:;����6g4���3AvhK��.������}$h�Pƨ���g6
v�c[����6-�w�@F<�t0e�f�bґ��d��ŷ��o�S��S����Ev�aUh��!�
^�VK&&���E8p`"3E��r���C`pJ(#c2j����իW�������$v�޶�+�S�2�'�JK#D�eA����۞pǾ28P �s��ʨ3(hA��I��&C^Aъ�m#m��";l�dQ����g�{[�ߥLdjv����䙈���������_--�����})���_���� �|@�B(x
l�'���\�����0�K�M�������z|n<���s�`N�k����I *H�s���?xm��`����`���٪f��M�d���M�q>��n�!����Q�u��[�`��q x˥+h��<��Eg��W��'T���O����xg|fg���X<�2^�A��tΊ�Չ�`�I2x��������qiу�=/��2���V+{:�i��/т�� ��F܅w߀�f�j������:�:�"�*�R�!�X�x߈s�{'�Vp��MbL�Iz�>.��tO�2 \�ﰺ�V����:��Bo�L@�w������>
������G�����J^��<c��"�}��%h�!�� z^��4�lg������6�uU@�����+��ԟl|���蜕�ҹ�e�:ƛ|�w ��� 3ILE?G���
�*�9�R�EK����:��J(�I���X����(+It��,,,Q�8����gϓ��LoR��z�k�d�{
I�_>��?�'�w~���� B3���%�NWl�)�ʵk ��!�B����[
��_N^��+���?�w��I*14��5�D��t���_��V�����(om���|*Z���ԃ�bN�f�i9=�23�Uv�8޿�8���){��E�R̢1��B�_1J��uT�7*Xw��,{v��c
��@̔]�Z׺ֵo�� t�k]�Z׺ֵ�u[l�&���PU>�Xź�b��d���18$���D�]���tF�n�Qt4�S�Π��9z��o��_����������z�G�������,
<5s.� T�
�@Ig�(�5v���N�!�J^G�:�	p����ϗ���+=Գ��z�}���:*N�'��$'�h�s�nV>[\�d^�֔�L;�7;�%C7�SP�ɾ����<Ѷ�N�J�q�=Z��@\�k�ko�/W��s�}CG$vj0``�NV��{=�L�����o�Ѡ�˟���y�����0��ayu��g�b �2Y���c�]�B���@��i	��Lǩ�=t����r&f��� �
�%ˍ�)�2x$ҳ2�T���������Ƙ3�
��b�g���Y]۠���CXZ^fp�UĆP#}�����n�i�y`�U�7R#���7��S�~�\�~���-U��8�k˺�rxPy�,6J,��)E�<��:�U��+�m��#F�V���V�ʺ�P�o	�0@���*�&8&`Djhbř���2w
#��R��� ��L�S0[Gԁ��I����B�L�5�%j]��>���by��xL����'�ф����h��"L'-ܺ���;,]x�}NlǺb~Vu{+���Ю��'H��=��/|�ӟ���EX[[�a��"��X�r;�.������oe<nbT�G�%���L3Up.{�1@��Q���Z-�aY�}d_P���K�W��ب��dj��l98�א�?�{�Gz_S�鍂�� ]G�[0�gTx�` y�X��i��,J�ɩ�����U�m�)��`���u��3Q�M҆ ϡeo���������Ҙ�2�JE�{$�O��- �=�Iyf��4;SKU�<��w4�D4����B~�>Ꟛ�L8f�����]��v�R�zPJk�¾�i��u���?+���}%H�qрc�2o��Mk��ʗʛ�Ujc�/�.�Ej�G��*��W4N���Hׇ!hі_]��͍�Dg����rO}���x���M�H�r���)�E=�����J��máu�-X��B����a�F��̆�v�
�(
�[.C�I�u�"}M6��6�]E�o�_z/ ��(�lCvĊ̹�W��>�9j��<���l]��Ϟ��y|d6U�g���l�� F�J:u	&�KvX`;��� <�݅W^�:|�{>�t�@��qYo�Lc�����Ag�u�^$� ����If��T������2R{�ȁT�8ݗі���"�@��Ep�� Z�@�F��@����T�#Ȼ�$��O�1�
-..��ǅ�Df�9+�X@����/ԫ�g-%��_����ϓ�~�r����4La!,���.�چd���}a��%S`�������?����%��]Ao.�S�]�U=UyG�of� ��R k��:p\%�5�k�֪�KٔG[�Ĩ��YUD/�o�_�� x�$���hA����R徏=��ϣ�k�=��(����`�^43�k]�Z׺��Ӻ ��u�k]�Z׺ֵ�Q{�i���!�˃9%͑�r#U�:���ܬm�A���rsa�{���7�|���z�̧>��o�z������Ao4���L �m&*�(�`Q��h@��B��1��P�$���D��w�����{�-?�*�G��)�l.�E� h&��-.�ю�K6�9}��sf��&�������͎�HN���S-e*�Ju���>���O�QzXX�C�_���Tڱ�Ղ)�1<��7���4�!pƟ�� ��D��A�剞�<u�a}�vз����&�ns��R����W�(tii����B�h�}��^@�� ����(�-ey�CN٭�|3P���H���wc@@@�"�{�M�䗮�!�Y ��Mz+�(��H�WQ�>u4�.��A�H����K����%#�Զ��9(��m���q�M�X�["�6g�8����1&�!�ڐ÷��ct$��C��ڄ��1�&��/|��$������c�����K�h�����{�`ے�Lle�}�=��o��jR�TR	�����m��m�t��m���f0����;�GӦ�nO�耆V�5$AKH�U��zÝޝ�9{�L�3�y��a���ҫ{����re��}�[vN�L��J��8ٿ�CP�1n��U�X3�ɞ#��K��Jj�G.c��\�����>9�Z�N�ĵ��Q:�Y�_K#5�;!?Hme� 0y ����U�<���	 �1K�#��N��F�`��D�_�=N��>�@sl8���AY��$t�;����=���9 b�?ξK�vU6�UT�D	ET���b���p���%`do676��{��VF�F$�s���iGT��������$�[a�s�>�	�R�ͱ�z"����j)��EQ�t��9H?��t��('����;�6���F3��� �7�����̣�3�}�	 ��E�(�_�^����YĈFz��ؠ��7��l����@��b�P8�\����ת`�^/�c�L�����B`�w���:��	4Dp�uDJ��1�G��Y)������T��@������mk���10Y�2G�v��&�?c%Cbq�zL%O��:�4�
���hd{�)M�Tw#78���e��}��� ��w�9�0@�$��9ӱ����/�+]��VB*��U���9�_$��_��,����{v#k���A�(�o�x!@�	�N�
�#]���,���1�Q�G�ռ�����wS���w��*�r���"ڼ�\�2�x����MB��kd�����4N�vGso��L�����X"���Ga����T��5(��ּw)z%��<�Ϥ�n���I�q���8Ҷ�J,xY��$;^�pm�L�6bt�TF��O�5�9R	�۾�;�'������63���kpߙN�����9L��&��i� s�tcX�a�R h�.[i�ώ��?�!8N�����Ԉ�4vx�Nk͌"+���S/�Ԛe�T=*K��r:��3����^C�7r��N2�y�����l9R9��7n�3��P	 ���"O&c���P�����s��C�:�ʤN{��쮪F���G�D�	�W'E��L0�~v��8-к���[8��J���4��R���6���8����7B{#�O'�8T�U|��G�=�J%��[��SZ�?�v�<���9�#�r=�z�H��d#���N�l�A=�����L%>�Jx�c�5<��ؼ_�\��+��aY%Vz��C>�&{8M��\�םi
[Q�x^�q?_���>�sy��'֡mhC�_�6 �6��mhC�Іf�|��*z�:VU ��,=�����"$ޢo~Tl/_�|4�������?��ٛ�_��q��Y1�5�%��H)j�N�E8�f~��1˙{˗�e����ˏ�14>$$p�gs��-[�T�2���ò���h���ޙ��� p�\0��A����T�9�D��)G���lxcvp���L�r6�!$����!��"K���z�3l�^L@�|�}�P�#0$� �[�������f�wVVV`<Q0���w��^��x�#��� 0��o�s�EW����E�����1d�D(��&�!(��%g߹��H�/����U�/���N-�6�mF)SS� ����2�����&� s�U��-Y��9�?�2�x���Y�a$u����G��t�c���HL��YZ5�q0�f���'��Yج��iG:�#��(H��G	R2@�eF4;N�K�}����Ʈ͡N����jp^���=�����ߍ�=
� ��L�*Aj����@飀�0S
2��MU!��B�x��k;�֚Tm��y�j�mM�Ͻ _x��>�#{�L�J��s �qLU �$������z�<����H��
�uIAjXw���ܑ맚�ɏ�������]o��Q?��y������0.lWA��MA[&��V�i�n�ޓEח���b�7���Թ�9;߲�����;��`*ۑ̕(c[)�*�nДl��ٲգ�����듮�E�-U"u��R@>�o�>��f��	���p�+6:O�,2)(()%�.�u��ʙ�ϱ=��ҭ���4J}o;�D1��כ����ZA��~EIP|���W� [��XH�{��� ���*�/�����&=��'�����I�<#��h"(u�s(�Q;�ς S���O	����Z�#�yH_E��j�ñ#xg���׌�rg��,eq�L��~$6.D#/ 0�	�[�2GB��iK�{ZK�qVҹ��,l�&�A哮bRe�wD�i���%Xv�r���� ��p.�4?��+�J���D������ Y�cT��F$ǿ��J %���t)��*��>t2�����[�]�3X���]��&�;8��_}�{�%X랄3��+g���֓RHD�x�ܽh9#쌴�gc���tsSIm�S�?�ɕs�X�t��<��Jjq��ҽ�zh�Q�j���6Vf�v�
Nț�����!�F�?U�RU=!�l�柀�����1��0;<6�1<5����;��x:������s@�c;���T@m*������a}:&���թ���8�jǮ��N��q?e��[��.�qt�h��Y�9O�����/�M_P_�_Oߴщ�<E�t"���<��t_�d$�������s����r��h߃�9��OOjh�WBn��]���}fR'پ+�QW")�c����l�����І6���/m C�І6��mhC�6s��c�ة����)3���8��2�	̡��&:�5[:�1ڗ^z���tz�C�>�x����r���BF����.�w�(��@�xb�� &e�'�H���Q�~�e9�ޭ����K�[A�%`ߢ�q�\�>X�ʱ4�$����!cT�lb
�S��4����ũ�p7ږ����N�^\�Ep�-b�
�z���o���ßQ���^@�W���X*X�~R���O��g38Mہ�_۰��AY�E��M�*2(���1��qe����~"bB]�lc��縦��z��n9���� 1ތj	�cHۉ�)8�Pp�̷0s�W���ڇٕ�U���^�C�g'�
�%�K�6�pBt-r�-R֝^K��al_��A�J�g֣�A;'ӣ����Z-��R~�2}%PNW'��Ւ��}����H��S�M�f�+a!��FFs*��,��x�CXg\An��A	�r'yf]Q����m���3\ c�K R����`��%&B�����{:^^2�y	i�2��6�7YJ]� �1�|&P�gs��j���MY�ܯؚ�)�MXY��!�C*�M5�琔�kЩ(q`	"HH4��ءt�;�<�
xl��Ws��1$��x�խp��{�Nz�2��j���"��J��P�cK�I*K-��.�����w�%��Ι�;�a����m�N�k��L�:f2��;TB�a����[�2�g��J��5�8*ȃ�G~���J��o3��D@%�Y�x�D����e�@�z2Y�>W�U]3��� a间ohҩW_��Vl��v���sɒ5�1p���9tAc�u�	(���6�������ɇ5��}A�׵(�H$9�W�x;�w�⼥���D����b�� "[�	h��
��A�ڤP� �;��Yw���*8@IP�����sH;��}V�C�c�c�>B�u�����(t����)�9Q��N2��w0΍�NǟW\ϛ�1lL�0;ށ����47�������}#)�ȵ�X�:��tKʒ�B�M״� ,uBD��W�̢�&�$@���򕑷���x����	*��NH���H�',���,8#��3g����}��pz� ^�2��0�E�ʥ5���H<�|���C�?�E�%J'�J{��t�ṳF�;}����?%j�/�R��.���a8[��N�]���6����be��3َ��ҿ�#Zw�dc<9�r� ٍ�|Cu.T��s����
Dͥ�:�Sy^(�Xx��� �'�Q���[��.��ri�׭���m����O3�[���d��k��Q��\齊s҆Dh��� JM���_5׭Ļb�S󍬔A��(���^��2V�B��f6�gY��'��y�3��Ә�FT��������R#RR�*����IG�%$Z��T��
8�]�[�{��І6���h`hC�І6��mh��źv�<� ` ��!?늃�NA��Aϩ�e<�k��������!\�����������G�Ѥ��Z��UfU��*.Ǆ@��b{9���Y{���|���e.��L�(r���=��F�A�"�l�Z���s�W��>K�kƟ���ON@M����}�$͵��~,�	��.��饕ј�J�@�U�;j>^\�-q�_�^�)5�6FZˠ0X�����m��B^��`��P�8��=��S��S��`_[0���������Կ�ؿEf�ȓ:��lY�AЃ�&$�,9�����%U�"�TvE���#N�T�D�5i9 ,vӈ2��rFt6�
�א�A �~���*M�H���
���R�A4�N�l���!���(�Qay������0�i5�{��\$��r6�Z�ւ��8�s��60v1�Kj�vrL�ͧ��@/�W���(� D�Eʅ��:�Clsy�M��V�E�E͟2N��P �t ��ǥ�
0���X�o$�����1��G~�G�۾�C���Q�#�)aA$8��}���9::&`����x�+_!5���}Pt��Ԕ��|���G!Gh�]��=���T3�ћ��e�{5U�|oԙ�~K�`�\�c
���ޅQ��J��L��B�6��#�S�SI6�$�,f���e�]�R�Ź��G˫z?�]�)]��s�u�Sv�|�� �����%_��J�ٱm���6�Yj�z����d������߹��Ѳov����V
"g�G];�k1�G���㮸6N�er�ʖ�P���g�|H-�!���A�Ey�Q��5�Jܤ���=8��V�`m}Ο;��p.�� ^���o܀���A��'>O>�8��X!E2ecq?���fN	%ZZ����hF�����|������`��������&�~�އ"�$A��
%Ó���-�bv��ƆF�Ϫ�xo-es�<�Wm��d���/�����9k��Q�y��J0C8��+� ��NE�N����	��s��g�9L��q�Rc�0N��ԑ���UΞ;�#�( ��F*�5�)�#�[�Qx��Jܷ��k[kpW���/�B#�	�TC
JQ�c!���[����F<�qN����7��/��tg�};����Q�c�'�N.1>b�7Q:��ρ��IH�P�I���s�31�;aϟ��Iن�����LWW�`o�f?y����������i�QM �Z�2W1k|P=y%�f�,�������]�{"�?K���(�ɋ�9Ȥ@�	�h�){�h[y� %Y�LJ}�u�/X�؜���{--���Q�����KC�Z�{&�xZ�}�<`�XGKҖ����r3
��l�L �'�pr|��Z�u�T��w�3%2/�L��TTJ��ў**��*��c��]I߼�6��mh��@ �І6��mhC�	 �X�"�s��%�E�|��-��(��n%�P�џ�u�ϟ?NǾ�N�Ļ����'�m����Pi�J��IG��˅Įv2�����d�3��5	�;=D�)��M�*S���˄��T��l�-��(2���P�����
�B�}�լR�6� 7�m����*��I������ǧ'2E�ڙ��q� n�2��~rNs��r�\���i�>��Z�٤��Hg}"�ш�v*�˘Q�<|�Hc@�d�Lv^��k��- ��o��)�L���u�%CL��%�:g�e�e2H�*2�%g=��@�Y!�!����@��R˕O��N%@_z����!���W�rt����u�Q�I(#Ta�[�Z�>k���5�5�7�f�� ��{�=㝌��t�	E�X,�NK���/Kͼg�cQԐ�!x
� )Ȩ�^�ff+p�W�#��TdaY��f���ن�X�ǚ��#_6g�gѫ9:�OQ���X�c^US
P��Y2u�9�G d�C��\�b4��ʆ�X�8�K%~AB�ʘ�Ev�����&]�G>�x�ŗ�{��{�w������ )���Nao^�u�Կ���=�l-6�u� 0�IcӲ��o��Y�*���1?��%�s�~��17�/���FŷA3%K�wv��_�LE&rUZ�#�:��P��P�G��)z$��W���|������)�k�2�;+%dV�3y���x�q��1ɪ��:Ț.�l���O��8cY�&Z�B�� `����^+;W,Lj��c~p���h�D.]�A֯��`����X�er0�+?�eױ� ����2zO�V�JO����S��%�_E` �y�s��hxo`�K~���m�ѿ�ci�O��իp�}������acs��I��5]+�w\�t	���cLJix%Ch����M��W^�����K�ɀiM����zrC<GLa�mN�t��x��ڛdr	�O�yF���g��"��y����}E�$A!����8��n;��ϥj��>����v��0� 4'���g�c����*�o�0�ZTMP� ��m�<)��k��4/.]z���Z��_ӜG�0������kV0�̙3Y�?r?��Ʉ@<��ѓϨ�E+!�pf�dwU�:��Q���, �"_a�*�e��38�݇��>�~�%8��"t��7�����tꍳ�u�C���\V�2�2Y��Zg3E�x6.�����W�,�U�pfo%��n�w_��2���pD�ykk��~I��|�K�Q�{��n;O���ڃ�}+}��!�Ud��uJ�%�(Y��Ԟu�qi%�K	BiPq�Tq"+�h��e����s����R�Y�ў]�A����{�\FG�L%�F�5���+�[�;�����N&\�(��5�TL�����{���1M����z��K9�@�XN���wvYt?����ҋEK�E�)����6y
/*X�˞uE'�'� �|/�5�n`hC�І�W���mhC�І6��Y����W��=3� ,���!0�(	.�XE����_�|�����dG�}��x�+_y|/q.N0��2�!L	�z�`���ձ����,����M8p�<F/�Z��ZV�/Q"W\� �������V���/�r��HU�׳|��5�I�3��_ם�0@��WnD$ث�f�������T��^"�}��#��\Τ1 �[pL�A�]�O뚖��f38<8�:ƛa��<�W�Ȁi���J�Zh�VA�>t=2I�����AP �@p�P������"X��?�o&};�s+����h})�^-oaQj	s��"bq�3���<Ԛ��2;PG�
r�A�J�	h����ş���}����_ �e�R�֎@O�W��Ȗ��]4�`>�n�>@´�>;:M.����rY1�J8�_�Ii3h^9��+�2�� ]�o0SR�Ī��j3*�������7Q�3��j=��-yC)����Q�f+�v���D'ʨ� z�kkT����hį���D�vX1$��*U������k�{�u�eM��mۈ?����	|�s����3Gj�cŁ��LȈ\�L����h�~<��&]�*g<[Y�ud0���I�����_����~�K��@A#]N<�� ��R��l� �ڗ��T�Y毜�MuL��Ĥ�4ᤖ3ݻ}1Z��
h1�E�4Dʪ���K2�}'H��iSW��LΒ�GJ6�2X�X4�8a>W^���:"m�?߬�֞:N,�k���uű��-6��/k���Ԭl-u&�l!�y�wD��E�uv o���G j�~����;NseN��X�i�8����d��R���!lll�AZ[�����������'��W��z�����4GWa4��:5�\�'��8���߄����{���� �\� �Bj��'��z]a���yEX���
�ig�{�R��q9V[�;*�;�|!�Q��4Ǚ�w�>8�?H~��֫o���u!Q�������[����J�:�7�����w��&������+����Z��T�S���h�䧴�:�CY�]<�����r��y���:�O%��A����z�گʝ��@�A'�#��:�/��������tM|�����U8���]�
����y���A�kuw�^Cœ�!	���_���`e�<l�~7L���@0�*��er�z�b1o�g3�J�fl6�ߡ��y�$�%΄�dr��T������3;>&b�[|���[.��?���gRb�����{��t�j5�x���6.��k�}��H��5�		���1he��h���4<������E,�c$c<�|X��v��s�y�lR�`E �_��X^W�2c��|����z�[���11q+�3Ξ�b�b͏�Y�+Ҹz��K�H>���6:އ��u[�q�Gk�g���=�t���S��(}��h�5Q�n����J�"z��I�#���\���+���ph8V����S�?���??��mh�6 �6��mhC�ІF��HS��4�kcp Ay�NjCR���H�k�$HV�xdDW;���p�c��[�v���x?����(�����a-��vp��Z�w�|�,�
@� E�?g���-K8���� �*�׊@�
���%0P9
 Qt�f�.�	
��{�-�e�vRg�A��@s
I�,���B������uݝމ��w�.��u[�jߔ��G����R�_3�5����v,"��M3����B���A�@�	K�`�e�T��2]Y�<ÜQ�$�H�[��u6��C��5�{ *g�ˀjqT�d�z�r<�#�i�o�W礜B���crOG���^pV�E0���5��s�h�w����r�	�&Ӣ7�t����}ueZ�����P2��������d�C��[�=|�*�������RpU�v�
��z���vNA{��B_�y�sW�F ��(�h\����g(�����Fq0|����D0��wo� 03����/R�_��d�He,���f8�W&�2����բ�c�v�{q,'���j)�в���Z0�(e��q�WQ�2Z�/:��bF?�h�h��1�Gq��<Q�A����31�L>�����uz�J	�wy���x�}v�}j�"������@!�!�Yp��c��BǨ�N�	�F�w(��f`"�R����!uĵ���(��4P�� �p	� ��ߴr�\Q�Z,�֗6��F[��ш�/���t鿜��9#5�t`�/շ����ƈ�f����� �QrN|w�;��r:G+���������0����+����[�= o\~��'>	=�v:�o���я��ʯ�*���.8>���O=�H��p���S?�w���U�H������g�3���T�σ��Nk����ٿ���3� {�=X?�z������l�;p�~Rl���2�.P���Oϗ�H��xJjA3��g�ߖ�WU���
��et�w��C8><��7^Ic`}sƩ������������f�-N�:6#b�j��|aӵMX�V���+�/`����*���WJ?������c)�#����D>S�� "��B'�p���)�h�ZJ�d>�L"�>��F�� ��^׼�!��R٠d������<�E�u�'�W��k�����#��k�Hd�6�{��x�8����^��{Z���ފ��KY�;?_P?�뻼�_�C��k�bc!*)�v�l[Rz��s�?���P���>��J���c���������H��� �q�l�8.�c��v���%���*"�zǄ*�U����5����xs�_��g�o��6=�~���evޣz��푴>�*�SK��%��'�Ǖ�u �w��$��R��T�*���[��Mz��ϡB��h$*NRƌg@/k��~�a��&D� .��ke�s�?���7+�Dɜ��Yu�	r���9�ud��{'Kr<F��U>^�'����m;����̕�UWu��G(AB��?;�����������O������ku�=�}HKs�]�v��r��wl^0������G}�<��5���w܁_Ѥ��qG�C����6 �6��mhC�Іf�J ` �s�R��2|���~}U
L���E9����o��|:o������������n�j~C M�T�}��L��N[�����93�Q��Xf�8��{���~��"�$���Te�K�صj`J��x%�V���@�V�E3#��8�Y�Z�d\;�U6\�o
D��l���Z�3j���~Ӡ�/�d�v�'Wh��.��!Lt2���+�&�6��`2^�lv�����'	O&p�����;�̙m��:kk0�\?���u�ul�e#�����j��e���_���"k��.������%��]W�`��α�4�Oi
���`0pM  �g��1�����
Q��d�9p��0�C%����z�";�ϸ)sK{O���n���1�1`�����㪆�&¢M6�%s����g�k ��g���8iP8��H ��6�E��T�*]�f�0�$,IĒw%ɰ^\��ş� ��� �D\�󸉰���n��:WK�TF��m��?)ǉ�/XI'�v��̴�z��Nջ.ȟ_Isy:��<5t���(�b1��x<��a�"���6�w?�3B�m`v3����c��ہ�#�NNN�t6�9�ܝ���)���q���\��3��hs$F�	�	�k��2.�����|1������3U��3��d�j�_�A���N�'㑥���j��y!��Klߑ>��u���3��hg^�T� �K8�d?�Hх,��3Wu]�r0r�J2b��q҇�>`�&f��L��֌�G.��e�g��5f�^W|���q����  ���қ�9�ٸ�2��$�;E`'H6z����=���L��u%�O��ommS??������O�G�(�q�y��ҋ�\<�C~��~y�����>��|	^~�"���}�O��������Jc�G������_�����Ƀ?����]���\R@�;�˶h��~?��?C�o�9rO���k�����Ƶ磵��pP�u8Y�dd��	N��KG����A=em��J{՚�j�=ǡ��k���	뛛p~{Bs���)�V��ܟ������(�HR'�E�[�fu�������./�6���ʪ�D�3�Q}e�|"���r��r�
)��֊H�I�N�*ɍ���%�K���X�B���[<��d�@o_I)����� U"�op�	T#8��g;�4+T�
��������,���|��Y�TY��Ҳ�
�,�����ľi�S�|��Ț�Y�lo:��M�����LJ���K���
�w��O��cKk�� x�mo������7ހ@�'R�	�� �;w�y�N�X	[G�G���&��$�]6��6�7hMD�	"�}t�<y�����c�?�2�>�q������k>:>�9P�|���$����*��	Ǥ�L����y�{�Ua�&��M�����t���ʊpy���D�༗��� �ܹ�{{{|=����G /�\	�DЊ�|������;]���ݼ<ˊ:K5�:P8���p�c�dǥ�yO���["2bI|?X99*D��k�M}x|���;�>y��|~6�k�� wFoZ,�o"����~^�x���H�����^�1����&��~��~.����}�i�^^�߻�j��
	ޯ₉�,|�,z�?��{�����d�ǡ{
X�A�-�\q�M$z�Dy�
:� �~�X,���?\Up-g�>���oN�@���]����x2۹29�z�p<v�!T*'�7�?J_;I�k�І6�7k`hC�І6��mh��ݍ���ڵ�B�E�$;5#(��j�T�j���m�ּ!�� �Y����d2�m������bL��{�Z�B�`����L��GVCr������lo��e��g���� ~����Z]�t�b/��gI.�l�� �y��K�B�'�#윁��4����*јj���[��#so$��8	.:�Y�8쁍
R�z�����I�6�"�U#��qC����AV��1�τ|
X���K�a�:����ppx�Y_߀��a{���I�j�5R��n:�2	�VA{�À��:&
B(���G���:V��bE?9E��q�9�%H��Z�Z(2t-*/�㲐R β�4���k�U��#�@a2��HfUb�Y���csfk`�Q�._3Y�Ա�$�#۔=���Ǹ�Y��I���ڌ��lk��2�sI���/�\�o*�-�fp!Rv'�3��I�5VE `�oÄ~O��we	d���i�c� ؼ�6Z�*���d��-B0������E�{h0����_�,E�UJ� �w!^����-�.拆|�x<���A���k�kE��+�����d#R2��g΄wdL�q�@��&�c�ؘ��C*���߅��Կ��hd�� S~��]�/���~3��Gʐ��ά �i�<^�' ��r���\�!�yn���y
%��D ͝.A^d������ Cщ�2$��w�y��3/���3;���R2B��fT�:Q����X�p���%�xQu��:/�7G��ρ+ƥ�_]����O��,p����b� ���dw�juū����a�8��tR���Qн�
���:`6�t
�YGۅ�ׯB۾^z��w8���/�������\y� ��D E��hTy��؄���_��?�e��ڎ����A*;GG',?��:�9r%p�·�i�Hg��t�#��ԯ�O5j�:�JPNN[NPyM]��t�Kv7�d���?�X8+�̓Iu�Z�� ���h�?�����HvY\����3�mn���mi]@h�ҿ6�G�Gk�x�����(�0Y[]e �R��
XF��ҥ9|��gh>�o�#̊lN$ޱ�
H������	��S����>lmo��h}@�	4]k�*42���da��pHR@�^�ר(�`5���y �EG.k�~(t�28�u5��d���Ӽ��A�r7���R%&ў�����/����U~�w#��Ϗ��o��q��ƕ���/�]w�Ac�����?��'?I o�<�8&XמG}&Ӊ��!a�J�tLBB,�Tj�91;��{y/����D�k"�N	��y����{�
����~�㰹�M�3��,G#��t�{>O%D�|"s���|in��&�0yQ���Z�E��S-��Ȓ�l��6�݃+�Ԕ��~˝�q�X~��2�=�
+/�=>;���p����X���둟���נ���T�a�*��`�(N�[�<T�,��ʘ������i�D�&�p/]=EVV�εmww��~������%����^��� ���OC������������/�h�����}T)���J�է��D����Aྡc�mD�U'{��"���]�Tmu�X�MS������#,S�4��m�z>oj�lG?����{�z�h�}<2��-'�x���s�=����Y�3鑘��',7`� �('�V�?��DLl:Vԧ*f�������6�մ���w����oz�7���Օ��t���t�����?����
.������shC�_�6 �6��mhC�ІF��;|�����'�k�AP��Q��@�.g�5I�1��j}���@{0�{���x4j*�ێ�؝dOd�C��f��@U�/֊�,/�2(�ٯ,��e�5�8��hH�@�h�G����7�@.��"�L�*���Fm�u�B3�T����Y����93gs+�4�-���Ю�0�F@����}�o�.�:�q�����=��Mٳ���8�ڂ�%�b��@�k��+i�R�/Ћ�^x�YX��ٳ�(����� #�kO�e A ���ʿe�)�� 2�r"w]�8X(D��������2���c �\�̪��3� �y� O/I@�X���9{h�b�R]`Y朗L��u����s3(���`z��XT���9׽G<��{Z�ó�3�"�1c��j9�9�;% Z�5�y��t6���3���N�O�Zyl�d�������j�����
rřE��=���2�_��`%((!�o �gzM��LZ3�
���5�o+�	�ep}�t�"C���3�����y�u���Zb����>)<8�q$���
�-�w�,N��H'��QZQ&+\��<?c�S�H&`3�Oa�5���@=Z��dDw>�4�6��V�%糤�}�y"���v�!�������8����o�`��T����O�ȒmA��9�첱ťs��H��b^�˄,(�,�˵K>�Z���P��D�<��Ԃܑ3/'���Rg@�@�t�$Tam�Ih�w�0��u�'a��K70i ��q���"��?<�Z^��1�^�-�쯕`�{~�@��g��BԃR�4�b2߼f?�\�٪x���YZ}&^ֵ#�����8����.��
���wQ���|��k�v��^�ݽ���/��|:_K�H��0�t4���魖�RHJ�t������������C�����?Õ54:U~�4&�(����Z�R�{�{+��Oڃ��m����� �M'�"���?X���!Y��O�d�׎$őX����F���c\ F�A_���<��e˩Q;��2T�+�K�3�F飖�i�^v9A+������	�U�y�a}�Jĵ?���Ц~�(�w��HE��]��"La��k����Ե�~��l~ݟ��z�Lo<_�ƪN�p����T��kB�M&�-�]h/m��8�Bxg��p�D�B�	�� 
"Lz��}�Oyڋ4��ցva��.��qtx��^u��d�_SVyGL�tE��*��W��dX�
�t�]���_JTr6���v�}a��:��}�r`������U�P�{N�_��wL���� �=�9���������,����>������q��t�_��y�#p��YVJIp:����	*y�DS���N�S?��ݏ��~��pt�O{'ܓ��� �O2�q�'��o�x�#��pr�G
$׮^#5�6��K=� ��L���5+��1�Lh.%��T��~;y�C�L�TKZk�YE�5���Pz]��B��w��@�C�f��m^��Z�~� ���4�/EUfP̈́�k��KvVղ��V.��K6񵲽���-e@�(6�b7�����k��M"ݰ
N���"�zh�6����de<~������7�qt|<�v}��?8L>b���ж\�.|ץ�E׊����ؿ4�I&�ܸW��@�i�4ԙi}xx��-�qcq�kcrt�t;V�'1-<F���;��BG��=Ҹp���1��,�U���ȕ�R?bI���$.���+�z��b���^��t��	��"я�&�;1J���5�l����ܾ��s�'��ڡ&��5ˍq��]����!)�p	�]���W��d�<?��Es���u���7���u]�����|������mhC�R C�І6��mhC��գ�?�gE�=�5�"�j
T �8�=��/�|0�˗�d:�46��ZS>�4��ț���q�z.?����K��C�X%@���e#�2�s�ɲ% U�`$���^�Y&�������kޮ1��F ,�o]�z,�FPƾb�W7�IrW3���Jp�Ol�7��uzŏ��-�j��d��a&�}��9�,o���.g�!P6�x�
�7Y[�����������H���f�R� �U�k}t���}��a�n\����u���ghr0�8��%l�z�����/} �m(P����* 7۷f%�] �N�K2���
2�{�o�D��$g`��+!�8-Y�3U�6_�c`��"�WP�R�CAh��(�jsMs2z�k>�[�~��)����ެ�)���^ϛ�(��+�@��އ<4Ϥ����:�F��Y�˶�*i�1`��H��ˇ`=f�6��vA5Q�����H
�+@@M�m>���>˝wl�'b�RZc�mh��(�]O�<f0�3�$�3��>ҥ�<<:�3�g���)(���-�{�Ȭ6N�naL�J��:p:��ɖ�HI�����&��r��w�t��.8�ҙm@�J�9T�"���]��rP�Y���Z8Y{��1�M�'�@�8��gp/}��>���� �x\��Ԝm�����B%[r������Y�=gk��5,��m 677�ƍ⚝����y[��^�}���>�����h/k��/�@��\��k˯�w}�w��W_���y�����]w�����ށd��d�^K���_�'�pޢ��Dw�����ZV�A��
LI姆���La4��s}mN�)����эc�.�/$�"@�Yᇇp�ކ� ��w\��QI*Bsr�Y�@w�!f�UԵ�^[Z	u�U&ca o��T�Q�H4�n��ٰ����L��R+L���甔%��L��yg��y�QLVG�!�d?���j�|���ޕ?��8�5ոB��d�#د�?�䧁���3(YI�r/�8$��OӺ�@~�����	�4o�#�pTn�"��mޥɴ�6�_��_"��R�#���󰵹�,1���VWI5�q63�g<W��I� 	'D�M�n�9�����_^��eK"�� �:7��͓M���f֐����s��[���7��<s�����0Ks�9+;��+�RR��ބ׫�֤�����������k���������S"tP���}���� B�tX$D|�?{���Z.�S����^%� �{����o� |�w~���H�A�*9oe�������7��T�n�ͨ�Q�1}������cy���-x���O?+i��8S_�:�d\��d���=w�}7�s�=pv{�x�Ix��'Ӿ{�ǯxFP%|~ah^K@�,N��������:��_�{$~�񰶶
�T&aDe;P٢�����2#,E��!&	T�G!�ǲ��>A���R �gDQ� ܑ��� u��D:)I�~q8*��F�g��� Ty%���2}h_]���v4Bf l��o�������'��')Ge��?�ql�J�F|���xN����`|�����;]�H�̐� Y���rZYoe���ϙ:n]��i�����*�����|��?"����Q_av��u�L��
�ڕ�I��U�!�8^��	dO�J�U��QY2�� q�Fc���*��M~��|�,�E�R��);�/!�!��K��� �`hC��zm  mhC�І6��͚c�>L���s�E��9�ֺ� �FۂFj��S/,�N��� �����h�k }���b>d׌z��g;N��H�!�t�ҭjv�2�|�# �������Ů��Ƃ�˽��$IY+��k:�,]�(@ϲ����������1��������� ���ݢ� ����u� �4���z��4�Y��S��(Y���9����	$�K���� G�4���@0�v��h�P�Pٲ��eV{ Y�Y�.�ÖV_�a&�d����~_�M4�7
H�1q�P�{�h�Q���
��2P'�c�%����{Ȣv�\���K%�����뙰�E��(�K�]�r���i�֪�N�3aU�c���XR�@��`��G�����6�f k �Ϋc�%C��[�"��b��CALW�n]Kː �a����V\�y �c��Hg�L���H�3�غ����`���d�ZӖ�L`f ev�{��yd��W^y0���bwf_��3X,��uE�(�+u���O�?��d"�l��s��?@��x_(��� ʬsVy0_�	%2��BR0ōr"��(sI'fAR���oKP�+�Ƞ"-���K���X����>L��lCP���[iO%���\GY׽w�F5`E|,J�c��bDّw�s�jȓ�s�� r<?��0Ic�ǡ�ǳ����q�9�����b�ǰ��
Bp�^(��n}�9�ϗ��8-_'u�([�(DEP�Rq�y/e��6��h�]u2n@�*f��v���'�����W���oK�VW�Yu#�U	i���޵ 7͜���lA�.\�����/�6֥_ۄk�v�ŗ^�յ9/]�B������J3D*�s��������r��px㘠���]8���ޭ�4��DW�钕�b&ؑ[.H�f+1�� 3P��tGQZm�#�6��[Y!U��2�Tg����:��-�_s��=t�-��f@pӉ������rǝ�@��lJ�@�JcQ�x�1�;wL���ޕW�HS�]���~�U0(�@_o��Of�<����H�B2��V�&|_���"�?W�5�>��&���]��>���%���._~�Ivd��5�R�)$�l�9�g��l���y֦봟���_�&]�Oׂ����4.5pY���W��JV���=�/����6bV�(IW%P�̆�9�sf�ڀ�Z��
[Tp3�i�tM5��\��7�KHX����������ams� ·>��ɟ�i�����4��=�����$�"�����?4��+IV�c��ٹ
W�\���}+6�`�-�p�]x�駓����V���u��N�������O�MJ����c4��y��\~�u8s�]|;����C���v	0��c�w�'��onn�]o��������!{�>��.H.�җ�D�m%ي��Oɡ�瓽�j����D�?��ʦ~A��N_S�3�!
�=�kk�0������1N�0Mׇ��P�c{{+]�����H�����:�:�/��������q:���� ���9�kd��2�$2�~yW�� ��:��8��$��E����i��k���d����8�ͤJ�tLceY{U�p����K{�\ɱ�3A�5�w�iG�{}/
?����ȥQt_I#�{d!N�3>��ga�^���M�Rf"��a+D|��y�U��w�qOQ	a��ByX���sb��,�.+�A�ܧ��^��̀���اa.�>&I�H۸47"��`��+i�Q���6���6 �6��mhC�ІF���
�9N������$VN��0���0����/�����*�.g�� �`�5�� �@
��D�>��y��V�%ZJ\	�[���^`	��{ �j�e���0&�)1 �M=͂��M����1�0
0�'�$�
0�4B?��-x��Ͷ!פ�t�nA�¨vFg�Ŏ�G�@p�@�`I�%}#w(�2h`��(�CQ�:Ȍҟ�mL d��}�
P'��������4E%Wh�����Z��1��,�F�Ǳ�\����
��8f�������I:[�P��3�b��E;��%��E��*s���9ӏt
��d����5q֚dC�D��2Q��h� �W G>�$�-���*�$#����-���:��K\`��Rq�s�dE
 9{ne����cc��w(p\Y�<��џ�2[b�h5}�.;�����,0�v0ʈw�Ҁ�s��}B��u�5���`}}�ưY4����+/�����~޸q@�U9^�M�R��i:ƌ�g����G���!�Y֓b����<\�~Ξ;/�4�P�9�)F]怷9��N�`M�c�O�\����������ii�2;�d����Y��ڂ�}[(a�rq�R�(HOu��f�Ap͓� �zP)fP�гf��c�fؚ��)A{(=��� ����a�X�5�Y�]�N 	�����AD�����	� �h�ăs&�\����=?k����ꠟ��G̈́)�'��O5��V!��
�i�'e�C��t��EK*�'sm�����T��(S��t���F�=hWؗ8i��95��)[�+O>	W�\��}�Q�>s����>�O����^|�b���H;�w��|�����s/�9x�x�?�O���G���i�h��~p�**n�� !r�E���냍��7��|��N����CY�u�m��[d�0 #��3a�]��**Š���_�p'��� �+�����1j4 �b@-�
��.�3\j?�r���D�1�QI.&��n�
�
���D�)�=���z��?�JC�3XZ��P���P����wQ���8�-��+i�I-�ɷ#� �Bt6'��K���+�r��q:�6�6���;�������Z���6g�·�`�C\�q�uE	��E���:�[�}Q��r�͕{(�� �@a{z<�y�o6ߨ�d_��Iޢ�|�m&W*����9�������R ���.����gd�'Gi�@ץn_,f�˿�C3_X��k��;*�`��~��6�����x���SO<�;�p�[[[��;�w?�H� jtq��+x���L�����o���?����^�[�8<�ؗ��k8��gΜ��sga#���d��d��O��/_|	^{���;�+!��\�]�A�go`,�m���=�c������P�E"�az}wgn@�*2�n��|���t:����t_�p���:��/��z'�S�j/���ъ��R�O �ߠ�O���L~^��iϒ��A:��K���	�@
-���c�}*k&�c�o�C��H�5#�" �K]�i��N_C� �%\sq����z?2֣R��Un��X��c�
��Ι//��2e��T%A�I��K���D�ŬR(W�|�iA��������3AdUrHZ+�8P�X(%�P��w-ݤ�Q�������3 ����J@WM�������}�K��1���?��mh�n`hC�І6��mhذ��O����Q`�/���٠�v.q�����r��0��؃(%ڮ! �6�\K�	���%P�p�2~�����0��R�2�(����+��Vo;����z�������KVkY���3q�3��� C��"=���8��ȡ��hCg0����':`<�r#���6�4�K��A=?��׀��2��'i�Xdc8	<V#@4^a�M�OU�Rsz)� ]N�%
�V"���bC�}��ܜ�3=�-q��y���bW�� �T����`��p�����A��������w6r�q�ws�y�]%��/�	��s��P� �z���q��Uyx='�YJ� O�9QF����Yv_1W{�D�.j�.'�<�*��%�,9���}��:=PѠs�[��L�:�]O�c@-@z�k���&�����u|�de6rM\Ǘ]�� (Q��|����_��W��7	�g�)����v����p�A]lT�/�?��$�[I��1��>~�
ü��¦c��2����dТ ��N��?D��F�_�|����0�9�f*W�[ �.^��/s��/{�8��FN�e�+�m��r"�#��:�Z����@ :�T�8k��u�mښ�@y-
LH�e(�(�d�I�^/�|:�Q����b{����݇7��#>��3���<�6�|�2e��ݎHB:�K���hL~A��/pym\&`�_}Y���������Pq��b"6�o�68/�y/;�K����Hn9��tm�@��G,�.>F����S�2ub뼗k��.�u<}�/�S_}�0�>��?�|�3��
QQ�� H��ŋ�w���;��7�����<��������|���ڕk�1��8�;.ܛ�q��3�M�����I�t�r&�W婘��$<���!cA}�!�e����y�#�h{��Ʀ��P�K��+�k��V�_���+H�kU�J1  �@]�ѡ��=%�����5��%JN�=�rΔ���tN&J�'q^D6[�GP�c�I�#Ѫa8�G^�Q���l11 �}OT}�LV���oO��P�,҇�G0Kv�6�֡/41��s�4fJ�c�8؃���̓O�<�p����� ��yL�N�i{L�R���(��V�����̒tϭVI��h?�*s%P(�,SM� �Z���G�rM,�Z�h Y������/�O�_���L�y��Ŝ�j��K��Ɠ�����`o�:����ҁ�P�J���W����=�8sx��%��~x���d���H�9�-��h���qK��?���'�h,t�y<���|���q;���M����'�l(#m	C'HX���[�Zۏ�y~������d���cAwRj��g]K�fж"6�l���%���եVI�ޞmq���g+���������N�`�\�^���o�67`cm&�R@��J��*݋w��؀�PP����{0k��G;)��L}�7��F2Y*���~��5~����}�D�i.e���1j!��^��_�� |�#�?Ԯ%�Yf��t�@�J�s�}z�d��؏mN0	���wB/��!�y���g��4��Q���'w�g�5����)���L|<c'�GS�¾#�~̾A���.�@{Y��Z�P<[�7��u�KS�FU|(a l�ox"���@�ϥX�e4���M�d<�+�i���vT�ޅӴN������І6��ݢ��mhC�І6��Qs�U�Q�E���98�� (+{��Rб�I/:���/��d��MS����IAl�\�SW���i9��������j(��d�O�����Y�KB��` �-��m0ДW�D����ւ>m�4	ſQ�����,)�K.�%&[����Z�QjX��g�X��s�m�{#�D����E�@j'b��POٍ��J���vN2�x��Ʉ�f�.䠬\��`��>���ek�
�G��fk���e�­�ѾX�;ck௻�>{�Up�i�6|��㏔vom����|;Ł,����o�&� ��M�������f�j��$ �QN����We)}DȘ�vr���zer���=�to�~ˀoy�� y�X�8�xrC���oK=�.�V����s���X�u�S�h��q�~M}������0����/�S89:�ں�&�](� ��8�1ә2���U�F� <W�%���?fӱD.�?CX�O���&��j�V̒lb1o��}��\�����q�/8�-�v�,F!���>v�	l��e3ۄ���g����32Pg���*ի���yHQ Jl�Tq*/u}#�,G��N�s$�Q	,��**A�`�BQ��ح��;��|���Fu�Ir(+��q/�ǩ���Xt$C�����"Pl��-�����z��'�E�(i��+��d��+��/�;5.�<���9�$���5�ΝIp�JX":���;>�IRէ�S*��@�_���L�k�w���=�O�J ��#����.���_;==�J��Z�ki.��������]+��.����N@&�  ���	��&�������p��g٬�*��
HT��>�����E�q,lS�j��1�ͷ��/��wV�p���ǉ����6:��IC���O���C�	Ю6�ۨ���^\�Il��D�#���%�m!<jq��),���Ϡ��y�k�[ /s��Ѧ�T��c��%�hO����	�V*ɎKl'G'�kPick{��0%��&�z:'���Sh�u$�9]�e�#�T���/���Cܺ���/���ޮ"!�B�#��u��!��G/�yo��) L���h��W��Xi3$u�ſ�%��`2=�Sɝ</�����/=�<��?�S�=��=�|�#�g8F��
NR?����g�\M$����G�6i�<M�����'�۟���M�D5Z�L�t��=R�~��Ou��.=f�����Ǿ����Y:fc~�(� ���7?��0�=mV�-�8��-�y4,�W4J{���
)?|�������7�-�
]N�*�����eRY����d�X�s?��BG@�%}/�{A-U��&+��
�=+Sؘ��J��~��_�j������F8w֒�|��e�r�
!��,���t��/H�U�{�TC>o�@tJ���zV���-޿�R:@m�	:��D�=�6��C�S�T�[I�����쇄��{Q2!b�>BJ��=v�,l7���)m.G�~�=[�� ďw�|�J�e�݃Qu�����=6I�9����S4���KD"S�������o�a�>�9�ޙ����~�2�L�x4����Q�&�٤�gi��u�$��{,��І6��I C�І6��mhC��
 $P��:'e�9#Sd�1�@A�V�"�=�Y�T��������k�u]5?�������ףP�Pk<ҹ�Kl����|V��{',@z%d�P��1��-�c��޹-3�:t7'#>	�e�{	Z�2����)��J�L�D8 �q�s*����ƣ1I�>��;`k�,T���@YV�K�	gE�1�R3X3��;�i�,��U�q��(k�c� H��d<�/~�$�m ����������~��D��_z�7����! ������N��b\�5���sxݘIZ�(�Q!�d�s��:6'����M��9%-�`|(��3W�K�ٌ߽�o�_��pP�{����!���s��-qr�^y�vfB� 41��5�ޘ�M`��(,$������@%��C���˙,�r����ѕ�����\o ���zIMR��eIS��v�K�V�	49�ɏ]"~܊tQv��ˆ����>�ت�.;��L.Ȳ�`@��d/vZ�������⇉�3��9���4��j��ŀyG��\�U���ӓ4��� ���"gF�$G�D�`ʥK�cĖ|QK�u�m�ؓ�-o�/��2�O���u/h�rU+ Q(�J�7�y�����<c�Σ��/�%&bD�w���3�e��� ��F\����v=��7[�u���y\��)pr���h�p�>�T���WVh�9�d%���Ks��l[�ƶ���F���U%��D,�*H-��-��0n&���_�eV"*	��>� 5�c�˶�S(|�~���ؤs]�t	>��߄�o^�t����C�P�?�|,��� ��<4f㶜A�e豿�s�����}�o�������S�!��{�^~�e�Ɔ���%�?�IwO����2@���W�zV��p����� Mh�����F��<���dLL�YƇ��EC��	��|��J�RP� 'pj�]V2��S��X1�`叢��:�2�E�4��̂4Q��.�O�Z���`�9H~�2��h��;�o{9���#H�Ԫ����R����zԅ�cE%&[VVA0���˩�J�d�#�r5����B�H$������v��`I��N����s����*U�+$���<�8mf��w`��k��y7���5Ș�����]��g���?V��-��1]���Q�x�зG}C��}����c�ًFGkXE��-�� ����	���g�����Ns��W^���z��7�|!i'�lKN�5�d�c?y8><��������>��؈��dɴGa{8�݅O~�S�'���Ҝ����9�B�ȥW_����E������Β-�H�>>����i��}�w}���/��?�Y�v�˪�Wy_m����wt�����%�#
k�M��e*+�֖k;Z�LA����9��~@�umB��ͭ-*u�v�H>�#2U�gܷ�?w����W_ř�D(�� k@' u����J���D⤪���D!����&ҥ�3�. 9�2ޥ\�B��9y��~0�RJ��[^K��zY}t$B��5�T(�UJn�{�>S�$���]Fơ�t2� d���7��E�A� �S�2iݱ��� ��9J���1����2�h2!����>[g�Ws�&�����9ُy~�1e_����3��3��W�ӧg�U��r�郗�0_��N^x  mhC{�6 �6��mhC�І��u�S<0�Jj-�(�)Ív~�*��"�Y������ݛ��|�6��b��������z쥐�>�S�!����\
l�5
�Cx(FQ�
4��K&���ޛ�Z�dwB+b�3��r�*�f����ݶ�Q�_ZF�4H���xFH�!!���ղ%���4m[�A���\�cU�Y�Mw:��Ě�>��j^ kG՗��s��Ê��o���h4�I�nN*�H�+X�;��7G E	�!&`�o4DW�b���Pt@�艱�D�>y�@������i�:�`rqqI��h0�8�  ��}&J���<���{Q������(�b9��FN%���	��_.ۿ9`.<�y@�1�ؖ��k���!|�K_�˫K�ѧ�������R�J���(���%ר�j�� ^D��������@�n`l�nB�2
�U{ ̇&��Z&�$���2�����4�����t�_�QwObL`îż��Fǥ���b�d\H"��<�WG��.�7��U )�gJ�̀P�L���{8�'eЌ�L�fѸ��[�
��QJ���M�Q�ʞ��8s���tq��y��(����E���'Wǀ�:{��·�����V�!���������� G90���յ����̉B;N��N��'3<F5c>_����w��{Dߏ��qI������,+E@�D:��������;���E� �d���p!�(�'zƤ�93��yՈ�^뙜�R���A/Q:c�1��w}� ���]-��% Z��3�iU7]qa'1]3�C����� x��9�X>�uf��}���.�R�*�o$���xIdV����:�����y�%z� ]W�ה�[ud
��z�X�t:�.\���z�@����r�����`�*p.�2Z�̽�#S�D�3�t����:`���	��N�i�K��^���G�����k��0�u�5�{$��m�o���i��h�2&q��N��30}��t�(���y(�DnU��CIfr�&sS9u �J
���|�̇E <��)�Z�g�
�ŵa��ߨ��ʠ��(�\(���
�#v� 59��`��7�Yj��2LNSm�1b�Ř#��}�����{҈Ut�ܕ���d݅r��q�dg��j� ��s�0#iZ
|:�t��9MEC"*��Xώ7r�y�40C�1ݶ>�aZ��S8Y��٭[��xL��V��N�7=+˹֗d�r83�C��j{�FO��]�Sy�����Cק�MaA���0u,�%yE�&=0���Wm���?��C*9g��:X��pf�VPz����~
�����+��B_x�m�V���Y=x������w~H��F��hEǢx����_�W�w~���+_�*ܻw��ǷuqyN�!?x��2�7�l�8g]Pj;��̎'�{�O�
ƽ�LN<���˄��vF�$?��ɰ�P�*�4���h'��.�����R;C3E[{�wn��_x^x�eX���� ݄��8л
�͞���0�쀺�� ��tPn@r%��*le|�J4�Ao��g��H��&N�r*� T���G�X&��,�B��yؚ�Kq��k�w%M@1�Ls`�=w��m�u�)���xPp�uY�c��N�x8퍬w�9���_����r�wS~OF�G>�eI�Rdl������a�X��$�?:��F�r6����;�B��&��������뾝��ۗ�m\/�=�[�M����=�l� s��\>�� s��\�2���e.s��R��|��:�V&�D��`�{B�j)�������r���ˋ˫��b�.�5�4rPaX�K:G��@�R7Z�yԨ��0,&��{N��-�n�u��� m�j���W�\V L%F=�.3��3�W=���4�D<K��0���M��W1�h��(7�I��fsH �I�ҹ)�o�r�aٳ�oΚb��Q�6
�Vq\���/(�J� b�A��@]�D�#
FB�{�t I"��>ԋi�xʹ���L`eG`d6�3�D�:|��1ԭ������t�U2���?{YM�L�3�:q0k
�T�̲&�!t�v�j���g�qPԢ���em�����c�d�����mq�B'���ӓ�D?]L QH@�/���b�&?�Ж�Aܘo�pPP��ZV����@$���E��	B+"o�H@h��a}ȶ�/ܪ�WJ��� v�"L��l
�>�[X�͍�Y%AqҚL�TAÜA�Hf�x����?�B�/V��Z-�Zu1p;C���"��]2I����*mh�^�W�w��?����� '�,N �e��XU�NQ^=u�v�����&�Э)���dC��.��@��P�+�BUK7T��:N�.��$�T����ӕh/ӵUk��@O�ft��=m��TLdo0�=x+� ��i#���~'FwYӤۛ�F�hl����=�n��s�>P``��p��- �݋u�#ˈm7��EG���X�%ǂΐ�b5ȧ��ɴV��KD��ӒF��8��(}�rx�xKr�/�pq���-9������X3��v��u�t=�?��ҹ=�/���(3�E��#sF���XǣkV,�=QoN>N����r2��Y
E�3Fۿk�����M�ق�2��m�INXz�u��ʠ��]��[�֝jp2�J�E�W���P�4����/D�*�e��+���e?��Kۻ�~�6}@��W��-���,8����B��s�dY�:���W�~E����/���VZ�,F�sz�
�
�gG�2K0�"��s�v�L�=�ur��sWמ��a:�G=�G~�n$@��S%��f������n݅G�;<[���^8ʚ�2�Ȍ0��ag���A�Q����E���gL��͋1��}~{���fX'Jك�mh��G�=[�>��D�R�$L��X�F��Z%t4�
�k�K��ԉ��P��������-x��w�L��J����g�!Y�*�U�ݡ��ۗ���������IFzd#g�=����%�m�����Ȟ�.��u������A���G�W���n<����b��*��,,�*��6�><=;�����?�,��ҋ���/��/>�n݂�;h�,�� �܆ku�&��y�9��gr,�G��	��K�Q��Hp�K��Q�=|FLy3�����U�KU�K����6q
���}徸�E雮wy����̉�of(<��N차��N�E\k���ڬ�PU�xp���^i���Tq�ZYx��II��Tr
�TĚ�,U�oz�@�������u�l�be�󏟹�[����+:f���}�`����:���㦷?����b��W)�x||z	�c.s��\n��`.s��\�2����'��*1JWW흴��!aiG/����)Ӊx���#>����-1�5�<?o6���￿ޗr�^�Wc�[9��N�" K �z�:�L�5V=�9�/�o�4��ЯaJ�L�PK�!5{�$"�P,0C6�ȱU�l(R�6?�?8������܉��2�3A�{ CP���F�7�ӀD�e-�3"�l�����ݮ�4�j\D ¢�Ah��q⤡c[=ZDs;� �a �v���Ǐ����$�@eg2�AP"+@�]������(�C����@�s�r4�ff� �
�[�!+~�П"�u]ܸ栾�{���b��_��Wˢc��Eͽ,k�r��1YA�n�w�׀F�6)�<�8:L"9><'�O yc�=E@�R1��sj@4PH�YC�X��f@��8�0 ���T�DPP�ȹ�_C�F
���5�3��H;?
]��<f:^U��ŢO�nuF���ANjMQd:] ����So��]���F����J�H=���|��%� �Z��j�e�������gW����b��q�<4
� �q�r�m��;==��r	��fr�4' z�G��Zt/��L7��^�������ް7%�3�e�ԕ�����s[��ު�m#Q��oe����k�� b�f��^W���8Ѕ=��*1n��#���j�g�� h����1	.����✞CQ�":�vA�u�B�F	�&:�@�#��H(���$򭘃��~V]��֜ё���Sr����PoqM����m�y�Ɓ���v$*iJ��d{��{��/��ބ{w9-E�^_���ǔw���r���0*#R����9����
F����&��f�NA�Q�C�ܢ˒��A#mǜ���B T[���D�J�	[���*�I"8�i2�g�N�UiPjqe`�t�m�U�Q9��)Y05�I�m'���m�?U�QTчΎ�N�E24a���u��]�^|�X�����O��\�����-\]^��B��Qɘ��rN7�^��L������hP%z���#�Ae��͞��U���x1'�n-N(���	tX�o�v��.����?�Xp�ڎ�_�~E�<HW�� ��H�K{�5/��yY<��A�� ������*����1��A�y"�y�ק�I<�4P}���w�~����i"_�������U����8J������A���L�J��2\��kb�Dj+�"2�z��6�gxJU�!d?ҸÛ����-�O|�P��Zm�&?�>]J���P_�eilzj�l�<#�Fs/N�U�~���㬎C0���4�I����(m �������;)��� �ww�b(~'+z�ŨpuR��(���/{8:^���	��Gp�?���_��[F�����+�����k�Я}�k����z�����ǆZB�;ݟ��١z���&O�Fk@ҏ���^4v(U�@!��.|&�[�qi�*�`30���Zu)�T��� ��7F���&�.��+a/8�t���/�0������~w"�<��WC���^֞Sё{�CǗ*.�xM�2�zҗ|���߹�:�i^Tud�a.|hgq�j�Y�OY_R'��Թ3U�C�)|��m�*���M����d�����ӳ����f��z���~7�7��{�|�٧���>�% @	5*�e.s�˴� s��\�2���e.s�� ���Oe��rd�¼�b|`G��W<eA �% %���'�,�a����~�n{Q?i�J�FjFc�Ez�<a�+�ar+���n����ҿv3o��5H<����?�N�a��� F�'��U�5���Q��5�M�j�ys
GV&vF�g�H%�R#!���H��ײH"�Sj_��Ln)��YV�f!��P'�(c�O����?��C����4Q�a")`�E��XnQ�)
��IIP#���σĲ���-A�2�C��D�2���.
&&�!���2���d&<Jc���O�I�G�A��.�
�p�N���F�k^΃і���������O8�L��� �H]KJ�j �}�7]v�;ٌ��S�N��I ��:M�}��U$Qۺv�b�NG�+�옖���d�o�\n�N��{��O��d��¯R��#Yk��X��Pϒ!Tj㼮<@I�Tפڝ��,�)��,wj-i�	p��p4g�Qc�E �{�ea�kUGt�B^Er��$�'�k(����0u�k��kToM`T�ʜP�P͉#�w��8�E|.�o����i $J�rV����Q�z� �j~�Hn��ۡG�Qt�(�S�lr���j��xgq&����W���^�/��h߿� �*� ��m�GZ{��}޳<�����S��I�@�l�z�}Jrk�z���~�������7�=I;u �8�X��0���n���?���O~��Q���F���5�ʸ0e2RU��B.en��0�=�S#m١D"�%RمSo,�v����8��fmUC��Kp�gB;NF� ]^��5Jד:�%��S8S�O`{�E��wˑ�
�bxn�)R�>��)3)�����U"�C�5�%���=��_�UȔ�{�T�nۜ"����cx��1<xp>isq�T��o���vV�Q��<99&v�~!�o-Č�^�9�W�GiT�{X�Vtf��tGG��a�</��H鎜yb�u92G6����<EB�Fڛ���`�2��tzrv��/�|�����H:���#5�#_���{'C��oA�"s��P'�'������L���'w�2�5�	>�t���+�$� ���`�\T	�-7$���<(w�[���[v�=tJ����F)'���39d�w��(�/2zȤ 5Ц#K	���`�uљL"��G�s��IzXОVebҫyah���(��v��aC6�R����|,N�~�(�Z9:Z����y�9r�"G���G�³O?�fO�A"<JO{c6�6�m]��8Z��o��7`���/�h_� ���((��%\���J�Z��*�dY������H���T�4��F�l0���΅�
8?��:�it:��}�t6���H:5_3����;ѻ�����̈�̙��8��:2��ɞ�祝��CL9���B��J7,1��B��۳�#�F��B�V�Z�.Ñ�x����~�GGGe�۶Kk��Ć�bY�4=V���䉂|��B$����v͢40�+������>�~1�:=�'��պ�����n�����x�����xX/����YS�i�^�������}�'�m.����M�.������A�G9/��<Xm�>ܺu8�3�?����ǔ�`.s��\�2���e.�� �*�.�D!1���`�^ޑrx�d�/�h��4��b�V�ܿ�(��z�[m ����Ow]:6âK)��ŸF�p���Q$v+F�	*U?�F���3�y��;����'��
������h�N�HP�t�ԀGXN�N�WѾ&}��	�%kRF7F+`ai��f�c�=O�/��ń�1�k�<����6(C�2��a'g���c92(,�44�:�U-��hA)�l'�,b�����lG2֑��:/�Il���wY^��B��8v����:�����Ӊ��-�h��:�:PD�/�
6��xE�������Li��x�b���x��x.�7).�
|$Ҿ��0�E�4Y��s�#i�3�\ul����I����h�4�t���Iۡ�I�;Y�����M�&�3u�я�����|�q�2�E�Z�m<[��W܇��`�ɐS��(gQ�$1���r@�h���>�l
|���:�С�F�5�Q� k�u�5���1�ꄃc3�P�~Lf �����T0�N�ǗҀ`DWap�(M<��%q ��p����Lc���,�}'����Pwhq�5P"�[u'(p�^G��q$�<�D��:��[a���J�m�^�3��J�N�3?2����iwJ�A��8��v�b���ɀ,�f����\/��h�[��n�(v�� � ����>�te���ϴt�X,4�����D����n�H�l������!��Jkzفv�=�� ��Z-9�!�"�d��=�.H�]F����.�m# ���l�!:{���z�S~C�(� ��#Oi+&�ye�b�AeB�c�x�ǰ��������s�W�eg��8��W�F ��F����ⷢ�\u�Q�?����Q�5!qj$ճ�i�Yǋ3���쪎Qm����c����у��p���}���M����~���v�9�}���]�s�>C���!Dٕ����^r	?��'���}������&�Ղ������zّS ��@w=��5;�A��~ԑ���C��@��.�e����y�[����8갃1d����绾�ݸ���s��Z��i��(�Q�/��gG�8$�	���J�����q��3��1[}���z<�C���!�W�HH����|���׵�@$R��	�g©�����S�1[v��d)T���;��s]	g1'$>�e9'���"����4i��/>c�ku 
λ�R`gm_JV�9�ZN��ݯM��"h]�ލ�= �i��}_�������~����ભtvY�=���އ��c���s�ܻw>��cx�g�ޝ�pv�V�u;STr��T1�c��������{��Sٌu����vƔ�k!�"��A桐�R6��r�,�F�T:g��Ϙ���{���C�������^,+9D"M^^h�o2^��MiAZ2윍��Za�w��ZU8=�8�#6޳'Gn���Cm��gu�gǀ֦�b���m���
�/����/zR�]�~2�~���yAB��m���Vt`H]W�y�"�k����]7���zU�~1���~�W�5z,M_����y�̈[W�������7vЍ��C��k�#�֏}�GM��}{������^[Ҿ�����w��m����M���"/�%����MӦ��s�]���e���;w��X`����3�?����Wf���e.s��\�2�������G^�������n�^�ۻm�J�<�B�.��@Зl�A����?|���s�N�1�un{w�캳��ū���k��3�;�eL�ad��Bs!�[a��Rꪣ����h%��p��	|��!���_x����'�"1 #ᡇr���K�^2�$Z)KthF6l��J��-z�-���aZI���PP!�L����e��Rt�(�䠐EFUF�j�aa#pb�h��'�"��d����D�cHu)C�O�-K'�=2={�� 	�o���0�:�|�\�(u:�0��d5I���(�2��j&���bt�b@�[J�i��rq����7�|Vܦ��cQ��׳�B�걸pG��-�*X���[e��?n���t���"�`[!��2�ԟ){0��ut=�	�O�2=��Nṕ����Ȉ��:�qO!fY�Qy�1��G�\��Zǥ�,$|�\4Y�N�� �Ă�Q��%pC�/�S����>I��=TeS��*NkPC_�r#E��.��9'����2G�����J�j\�┡�
�)KD�������o�f���Ut5�(`NU�>z�0':�<� �S>efu0)L�8�q�Zu��z)�^��trk �kq��$�-R��Y����w��mX�Kx������.7p� �j���&�?�E7���C�J������Nf�x��{�6�̷~�>{��I{�̋�nS ��7�Uz�ɹ j�>�.��,��>:f��j���b��N���-%U�A��Ձ� ��4�
�E��{pV��d@�B�(S����]%z^r�;��_l��Jc0*��Dv�TV�ي��t��)�o:�/���|������h��Y�Ł[�O�bd:$�ve�ncAL�~���*>	i�1B7c��vϢ�о;�`��8��U��q��� �F�o<��6�����%���B�y��g��_�292�9��뷈A�jsI�f(r�h����6�#E&c�w�����W���`�ْ� �o-�������9��۴:�ܶ�(_�
z����48V�E����tJyH2��s�#P3�m��oo=tx.�	o�$�i�;Y9̴ �z��Ȉ���m������Z��p��=���V=8��-z��b�g%߿��H�:»D	g�bߤ,�$=?Jڕ�W�Y���)��:�=�7eIc��H��H�F��	��U�:�>q��<�S6�N�G��C�����p��Q}_��vJW��~E�3~�;�א�ERO��'��3?��G̀���h?��k8Z����-8�u��w�Rt� �k�t�O���W_�W��e���qfd'�5�9$��*�0��EX�a/z�Y���q�?~���~����r�Xm�'��/������"-��M�J��"wâ_#�]j���q�/�������܎�Q�7}Q��M�z�E���\��{T�8_&����'6�Tٙ-W���5��+_��Jk{_{N�F�U����^��,u�������i�Vc�Q�;|C�]��ZAr��i���A����O:9�g�e�U���=;�D�
B� ���r#� ~߃~F�.���H.eh��~_��q���j5�wÐ���S�3��%��\�2���u�� 0���e.s��\��T��>��_�V�f���K�[!݆�V}{k����w�,�v��݂���"K
��WL�]ʲCnO@v�j������߯�O�ٟ�����^��Y{�ͥh�F�
��B��"�!Kv�89X����+H������|f?��e3�'�Y�qN�5�k�	 ��+��B"���>�5 ��X<��%$ހ76rKd0jcP�a�s̒������Y!(����fT'ӧ��2+8��>U��2H�`�l�pT�Lh��*ґ��(��U%Udu*_�U���8��63��4���+Ul���8��E�|�z�
���	h[5�
����D-ݔ��bm�:���d5;ߌp�WЕ~8� x(�� ��������ſ�g�5���l�>v&�$m(�:��4_��e3 :P�j,�l����Ҁ`͑�9�����%�QV{D��I�u���6NNK�����Xl �Nt8�J4b�ʆa5�i�P�T���0��G.t������a�����姶I%��D���|�%_�	��2�T�Ь�]s8�����h����]�	 *�~�U�P#%3��ʩ���OS]Tյ"?E�m�S�Wo{��B�<5:1�(F�$�k�i�) gt�}F��T*9+�it���zP����uJ[�Z�x�	0�g`z���5����� *� �����G��"��=���Dfp
��H˻��Ai{��{wA��T�}�R� l��oL:�������uq�SB[%���a2r�H��G�Ry��:��*l����|�E����HW�0D�D������$%*kV���<`g4�E�?=I�u���em��+a<y���h_k1@���dfiL��EUJtտ����*I��@8T�&uz,�r���=B�C@?��N8J��e�#%dxp�Gp�8������<^ç���TA*{u�H씃}B����}ꌭt?J�T��NNN�Rp`
�>���9]K)���@� �љ�kc�\�d�'�Pbʀ=\\>e2�J�?����U$w̺��KZ���1��4�Ѽ8�Hэ;�����Y�������~��n�ڜC��>��pvzO=�X�~Vw_����؟0C����;t�Xf�j}�t�Gm��YS�,|X�(_]�}_dI����`�%݁�|^�'�tp~9�Fe���Ou��3���΍ֹ�g���;�0˅�Ϡ�N5�]��E��+��y���-ר硪���ǜ�nd�5Bg=A���G���r<$@�J��Q]�Ł\ׯ?'<7�È�E�QmL���*��x����/`s����������y<K��x��{����Gpvv���i[���#X�u��O\��~ծ�8���:�(�>���~Vϝ��C�kt�Y�:"�\9{���3w?8:>yk�}��G�r�/�{ަ�qC��5m�x�������}{6�j�U�c��6�j/n?u�'�~���m����R��5rx}�ώD����"��S����p�|��i�M��� Ϡ <�Ϗ??볉����?O3�\�2�����`.s��\�2����'���}��G�ӔN�}�����n�vge,wS������j�T{u�W�6~�z4�U����A����!�w��v_O�e��jW�������>���̥˛M��:dX��?���ӻ��o������k���q,����D�7��@��=�L�,��įn��+�AM�q����Yi�⌆>2�ju�#E҈U��L�dxr���
�����E���N����P-��0ưj{���q~c4��Q�뉺R�����L��l��~� �P^ʔ,j8+-��U����:XϯuV@}`�B�-0j�QZn2�A F ��I��mрnQ�.$.i2�6�:9��T�qI5��I�S0�(H�9Q��S�`>-6_ڐ8�a��J�4�kx_Ud�C䯎;`31YO�a���4�T��<C�]>
f��|�f�r)H
`�f��s q�M߸V0bQ�I[{� ��R������M4�m�)ƈq�;�'��tuE�؃{�t\�-��0&��*�\���잌��Cӷ���Q���B4��@R|]�o�1GX���cK���?'	�ɋ�e�h�1�����e4m����׳�_����& ��.Sՠ��sPm���I�2���`5���@���r��e�1���`8}O	iX�Ϫ�h
���{��s�V˷[3����Ls��!�5E��<&��d^�t['L4Y�_���.���WQDm��XR5M�'QI�h���Ax�3����4����� $�#�v_�?\�L�O�t~l���tթ��$%���c�o����	XԽ`�<Va�(���S}��\ ���~�N���^�`^�s��N�����9(�,�G��p(O���i���w<+�S�_�kI�L�}��Ge��d�<�s� �I#����#�NU%�l����s���2<�`|�����7_��G���S��.����[��U��b���\�:B�y�i�svG�'M�O��O×�ju��"� �~��F�N	����1�#F��a�Ѿ�������Qj�v� ���c\'�7�.`��GF�/>�"|�чt�~���՞΃E��G��l7�n���Բ��5;��H"��f����q9Z�����;_lkz���A� /�������W�����=�<��+p�ދ�I'p���$�l"x�����*):H��ꀫEA�m���_tu���#��d�ee}��nȫ����([/~�3��?�<�������h���T��j��9��	y�e�gH]�QW�Xg�ٱQV�����[z>��ߨ����]�a�IG��9�;W�����/�9L�C;����W�mq����}�K�܉,ʷ���To��W�T"�*W��F�ʩZ
3���,tz�s'l�䌷���~���Z�w,������dLVmM��׿t���������W�|ut�/�|�^J�U[�;�QI��~�ht���
'p� ��F��Qj�ӥ9x����ɋ�#�0x�ݱC��~�tܞ����g?���7��(3�?�����ev ��\�2���e.s������o��߻w�^�[�����������Ǐ���k�=����O�7�{�n�y��/~��Ǐ����D�z��|���=�r�5��I�����b��[�����_��vݾ�z?&�~�E)��a;���z|����x��G��]^�<�c����)��a���"bZ0��Zӊ���6z�Ԑ\#�fw��- J �وÄN� s���ςI���ܚ�� KԮ�7��R��c�Gn*`�ѭ#E-��W��f�0�(fs�O'5$*`��!�&�R�F8�	�`ԨI����VΫ�9J2CgR
�T�┍�^YJu�g�����G�jc��0L*  s�H��W�}h�|�����M{��KL������ܰ��I{���$r�'tೋ��$�K#�£�?�A�
@J�dI� �{b�Nq��|id�ϟ���R�BrPޝe�õ����Y���#f����Ul�u7[z5C��6UpU�]#���d��o5�W���l�Y�k�ۓ�:��s8x�^5��%�+%�Y��>16��U*lq9ڔ���P�"s�(�F��1�1:ՁAf�U��I�`jD�߳�/)(ec�7;����})x���,���X�����͞���
OH���(�C�!�^g���1w��gq���c��\��8	��g���a�����
	�Dy��9!�F&���Uq@�gp��s�;���d '�~G[R�㹁8�=��룥 )�b�I�d9�i��<����|8 � ��:Y6�t��QM��P������:
�OUv�N_�g���S'k�~�5�P��ԥAeT�R��dg��Mֆ��l���=��@kނ��� ���º������z���5���efP�N�G�	>�4�7;�p��"�	 G rJQ�EG����%����'prz/=s��]ö��?��#��>�<��+p��m�wm?_�c6{�v�l�`�o�u]w��&"O�_h,0J������Ϯ���dv&q����6��,:L�3�Z��w�,�@ತ(@0r�� A��g��~���
ZA����#�=;��"��f����5�?>�?�~��}8�����K��cB (�k�S��c��v�b<�=�g1�j�Vwa����_�{�^v�}s}o��:��ƛ�Λ�&z��38~�6<s���~��{��m[{z22' �Ya��}T��=8ӄ�#�ɺ��*_+|f�u��`�.LD]"OK갣N	���1`z8��ǃ%>�S ��Y�^>\{��{Mp���b-��&R�;�Dʹ��� ��t�������0e	�Ĵ�`(;a	����Ӛ̏�DϢ��r:c�w�ֶ�+.�3 3�
߫.�I�ޘ�����C�,c�<]=mI�g�{f�J¼����V�;K�B[pӟ��q�@G��뎾����$�����c�Փ�x酧��[gWw�?\,�?�n���>}�6�W�V~��2�����]f���e.s��\�2��iш�w�}w�^�����o��o��>���������3g��n߽{�護�^�_\ߺ}����NK��Q�4F����puu�������~��/.֏>xi������.//��ۡ��?|���hq~~�h���?X\^^-6WǗ���n��n�l���N����熏�[G�&Ԓ�U�l�ǹ� ��bP����LO�F�C�N��h�� �)<���GV��B������-�n��f���n�<��t�l5�I�kM	k ��H�"���+ �����ߕh�#�p8NIk���!��MU�\U#a��':i�9Fcrr���aQm�"N�U�I��"B5|$�mѰ�)��5����]�&_/�S�YH�!��qx�������\�'nJ@�:�a�#��@�eӑ��J��u%�[���Z�P'�`ffI&S ��2UX;��K4TA��r2���H�nR$2������T�ԓ�?��W4�Rf����*�J�k��Z��rע����8x�+�L���}��Q������H�JՋ�
��k��)fX������mz.��cC~��qq|A����Bm��c[���Q�	T��`z�y�=A!�����Ԡ˨Y��>Y�'�����9�hֻL ���P,+��{�h�.�&諁i��a��WT^u։�:3�T(���ê��&MY;�::���^�Cŏh�qFi��2���%�+���7X�ؑ�r�S

��f�@L1Sl�+;W_������� �w�N��ޤ����U�C�"�4���d�� �r�;B��{�n}.��X#�-�g��'>�G�|o��TT�X�,G�1y-�*��`w�=� Q�5�:^��A�)��
%R���)�
p�n�Ȟ��=U�7b�)2�����y(\ۅ�M�­���~�[�������
ܺu��o|VGg�<:�:�Ö䳎	�]�n�%����a���vƾX��P$���֓@��1+�|V��7�k�/~&�m�t��@���c��n=�G��_�V0�����3 �ql��(W�<y}��V�
������;��{��/��"�k��	���id�h�xx~��.�y����6&��Ԧ��Ohg��=x�?_��_nk}c{yp�!|���Wo~�/��^�*|���=�����"�����T?����~�|-R��g�68&_���J��'��H�UM��O���z�mK#��1F夊>�Q&G�pX_�o�:����q���H��"���#��Nc%�[5����p�4YA�/�IuR�0f���J(wc�w�?u ;��~5i~x^FGA�O`䎳��~�M�Ȯ�~�=�'�Q�O{/���:'�;�M��#���T��f�>�+2�J�}�dP��Q�uo׳N^ �@���Ӑ��X�m�
)����\�2��� �2���e.s��\>GE@������|�	�쯻�;���z�7��ٷ~���]_]��������q\|��7�K_�2����s�"O?Y�}Z�2�%4�,%��I-p��UkQ���yg�;���ϟ_�ߺ8�ޕ:��g�e��ǲ(������~��/c�L�w�J`�F ��?�]4 '�1�Z��<��S�I��n��dK��uީ�����H�������N򬪩�%2�A�G#\��W��	F(d��>}�^�4R�q"�Dȅ�T!�d�\�Ţ'��m�Y#���|K:5̦ �T�jȴ9�[���H_�A�	�"!j�9,�����}���>2�]� #�R�V�7&'�1����������'����(h��h�0�͂JQ�j��� ��'����F�"�%��l�
x�����-�d�D�%5VW��#n#܆����]"0���
0�s˃# ج��]N.T��9BA#���>Ot��F
$�86b�Vp{Z�g;`��Qā���%�?DF�1Q�I��D��%� 1�G��R��N�`cP9h��Wl[`D�[0g->����  �D�iDzfж�}��m���>�������_�)����������j3U�~���)���[�O�D��Ä�B�r(�[\�o�12Р�t7ŀ"�s�^<�LQ�������@�K���ub��Au�&�x����(� ���h�Hˏ��D�F�J$s)
Ԏ6W��uYp��;�I�����i��o�*E���B�=��
���-�1�iҽ�$�����'�aJSCѬ�Z��qP	J�9��n����aZ��S`G��X��٪�c]'rA��I�]�
�%��gY&;��5���'���U��e��[�F�b}tg���+��V1�z�?�ϝD��s�6I��}���Y��u�3��m6U�`����.Sq��s�F�k�;E&9/J�5~Ok_�4I�Qd���(VV䀙A��ܴ����d)��J�}�k��3������B~�ݧhadŐ�{X0�I����ay��&��~�N��y����w��Ҿ��}�]��U�{�(��1���ic�Ӻ�;Ƒ��lw����wvDY�lȞ�e��I��aG�S�V��;wd]��Â����D�Ӛq}��c(�t�ڽi�D�H/5]���@����c8��<��Kr�cNB\87%ÞtM����<_}�%8���<~��*6#���'�C�������l>�(ɒni	|��5F��:�Y�:��O�wʞU�AY?������G���_"d��W��zP�z���OߣR=�Weݱ���R�s�9Kh�a��fFgf�j:����|n�fҚ*�y�3=�y�����h�7�⌆o9�)��89ʹES�Y�I�x�
���l|���ٲ�,��KU_MV�}��8�)���e��X���,���p�(~г�~��~��?1���XN^��R�4>��#�Sx�X�y���U!�Ź�e.s���� s��\�2���e.���z뭷no?~��ѣ/�����w~���G��\]���񣗆a|n�����d42~�;߁;w������M	[���8���a� EC�0�����k���6�������U�r�Sr�Ʈ"�@��[��{���ĆٚFP�L�"K�>�����BA�`
J�MG���������62M>��R5m����f�e���������y������؅��Y�!�hD�\m��̌ɌOP��x�H�iUi������	�Oj\��J5Cr�o�͐�C�)F�yT�� �Z�:���	(�ٸ��4l��8��CA�5����-�����ɀ\YX֪A �pU��C��SCh��'�T諰���O,���n�~��{6 �Şd� ��'��S�G���(֝$�H��}����u2��i��(���
���P��j���\?
�l�ز��\��q�!��5̽?�g'��du���d>���@J������h_]�|Q�y,2Y�����ֶ����9�G' �����z��z���������׾����܅�w�PJ�G��z��\�Wח�Ek�����7���C8��\5'3�+B�җq##z�rY��S�ɩ��?��XU]7 �C�~W��(^�iԿ!G���[�.�6��BZ��������ȸ/���g���Bթ� �w)ݏ�x΋8PX�ߛɉ �-b��@EVƋ�nx\T:K ��ő��&Tt-�'�_l￱߇�v�u �.G��t��4?<�ٮO&KI7?[�&-�%0�.3`��i}����v��vk.o]{�ߴ't�G�zu��t��׻��=}�O41�a��a�Z��])A~���cϗ�~����5�_�sGH�\��A��ߨ\��%4_'���!O?�X��Mh�9�WדIF�4�����f��K���A!qʀlk�A���R� ���k;�ګp��������=��Jgn;!e��t��w�=,�� �]��ќV	/�Y���t�ø���e$ƣ��売�;�����p��=re��"$U�x�N�F���g1vA�G�r��i��:�������a��.*'[J�v�{�HM���Ϗ<ڷ6߅.q�z)���;'�ð6j������������mE�
%��q��$�rDN;��z�+�����+�t��sЁ�UN��'�����%��t����*:8�ױVZ����la�4�
d�~VT[�f�?����_��H',/���[dII��omXtϓ�����.(�I]a�	��*�$S��%M�alr!�I&6w<P>e#R���.�E>��P�9���+92u4Qݑ�
�2���e.?Iev ��\�2���e.s�������������WWW߼>��7w���/�q|z�ٜl���n�GP���łr+c���~�� M����zί\�0̔�!J�)VɌ6c����n�[��B  6΁��YD[n��R=�͙MDEiqA�����F��`K�@�ԘMT�F]5<��QYo��̸#F����n0;D��scަ-
X�a�u7[9ڱM�Q
K+���2>���8X3VJ�6�I#^ L�82)/5BT��F98T�Q���D�R4�[#�Lh�J�8��Q�Q�ǀ�I��%�R��P�NL��-$�19*ҿ���\�E(������Z�D��~��Xk�M㭶)�Ag�e} ���dn�+����-���i�S�	�ʣ�� 2_)�$Z)Sŀ��RŸ���>�i�`��k��H�Ҽd�a�f,�m��m)?�2W�����ͦ''e!|Qݘk�<z��f��F����7�"tD����
dt�P�Q���#@��"�΋N��ptP��bu*�HD@�_���q�(G&�B��b��%����>�~������ݻ=��?x�޽K`����� �g�p���D��m$�W�	���33h�ў�
��ѲE��SA`DГ����ѱ��ę�=�$�;_C�|����5���Xb�%��_�N�H� ��uAgBVza�P�D�$�=�V/Rs�s����H�2@����� +�8�	%?��u0mì#" E�Z��k�ɮo����hm�b�z�H7�au^��3��f�l�Qt;�h�x�Y���0���:d����<��r0(U�,0�8�%k�D��2�MTl�4-���'�Ԝ*��$#�:Oۧ�,!�8��!8Nf)��06�r�,�\�LTe�ӆ��W9���E���S�JF��f&��������g�#��_
��H��D�LBU�C��O/Gx���S3�<�s��`u��A���,�`�:?Pmlc������[�ȑ��
��';>�=;]�������`?��!ʞDj��FeC��"�;��/�PH0`�sVܽ�o���I�f;��'v����
���'��_@cu@ȞJ���x�1�a���y�=�Nԥ��$;�d;��������{k���T�=�L�T͓b�������Vl���B\j.��ڵ� ̐�鎦}��o!���Dy��:=W�Y�n����'�����]�������JqR+�2D�1L{�d-�.�i�j�{�C<������I�D�˩,o��t*�8��Ry�8��g�?E��}T���0��u�͹|������ho�2���e.?)ev ��\�2���e.s�����v���'�.��~a�o��^���8��aX��C��,Q�c�b7���e��lD�{�W(FPcE�{�P)
	����f)�{jQ�g�z �,'3r��M��������2��`pN��D�r��x�G���:="����uU{���xTϓ����4J� @��jv�5=�+燁Ҧ0��{�舂[j�<�[�Sg(Rp.m���s0g1t��RwK�vb�]J�y����2>s�g{����o�(T5�kN�n �%1W�)pg�hVCs��R����ϘG��QKy@�����8�{7)M���4�C+jU�����/��������T���d&HŴ�θ�7�P�7@'y��f鲐��o��J�鰦S�C���,7Y�\��P��/}��U�7�q�}>���`�Wp�����&��7 `�I �?LG|P�Z�ʎ��z��s�:U�ؿ��\�Fc��ֆ~*}����}����LԹ)1��SdO��`����v-��p��o�C�*|o�}�����J��H�Ɋ�i�Z�5��P���(��,�K#Qy�YjZFZT_�4�������]��H���� �sú�@�ݘ�ژz4`�1�*�"�[�;�@Զ�d$!�j���]�9��(�-���7��E�\�	H���E�Q��i��fD~�Dq�H%Ix� �lPE~:K���t��z%
�m���&�G�V�%A��}��z��s���IEtUN�����1���f��~�?�yt�JhM�.y��E�U��o�~;Lվf�O�%o;ɯ�u�*�v������D�W��=)�����	�-t�h����Ax��Kt���F����8���
1=O���2���Q��!�ߝ���}I>�]ư�}ɲ=d�G9�#��k��FX����!��B' Nˀ���d@�2�2�X�M��}��гp�6��6d�s�b��s��S����������G'���ڒT-�-)#xݡ�D ���Q_� �����z��3�d^P�ӶQd���{%1�9�����Y�7Lu������&=3��K��X���d}jN�床�۞������Cy|"�~p��������k��2�g���RB�R���Xe���3�\'۽IΝ�n���I�HJ��S
���ȿo�ߣ̲�	9����,�]9�˻J	�9�pv1�lU��u��g�0�O��ф/R�`�Y*HF�jN�tI��-�%q��s��%���Nz~M�s��C+�>���I����e.s��OV� �2���e.s��\>�l�0ܩ)}+���r��P����}��K`
f,�:�4Ɓ�'u�CE!��+E/�0#,����}r��� 5g��C3\��R���@@��1W�c�Z�����0�=9���2&��ُ��-���̷߸M�8�K4���Y�#�#��~��J0���'�#Fk�v/�23�T�Y��ю�j���=w<w����K�Oiy{���4�u��̸��3��Vc�k�����pJ�@2�E(0�І�2c��f�s�V�NC]�H���h��y<�lh#g	��#�{)�d���a�:x��a1�e�y��������=Y��B7�.��\1�tp�~/���^S�n�'M�
�.���1�p��o��2�����85�R��C@���el�mY�W�t\���ts�U@�h�%R�;���ܜn�1"Mڠ��&�+9��<G��U��X��9 �|(� ؀�8o
h$�C ����f0���T��_·��-�ٟ�[�������	���}��)�?���ӣG�������|��9W�;����@��F��s���C�{�������C��ȣM P��v�����@�Z���ϟ��5� ��8�3�]�nBu0#�lNElی ��.�*-�g�� D���d�4+�Ug._��lí6����'���hh���ðܷq>q~Ǒ�^��9`4nR�b�[� f6!z�d���*%量gL�a:#�fk6�:i���&ݮc�u���i����h�����Y��hHd��7�]E)��Mx���%�	 ݈ 56�Br1 ��P1�|�4�����I�����f��� ڮJ����Ce:�b�
F���g��0�_����Y�}��!�16us�,����Y�h��y�u��>���v��$�����gE!�G����l{�9�i����P6:b����e:i�lC@�r���]�0�u�/(z��sWJ��T<�������Ƕ�Q�-��g��E}�g����v�
���V��*2�	��� x6��A��7��Q�fe�#�crfBj���w߿���� �Թ.g)�rz��!}���e��̊ �Mg\���\�|�4E��aa�"�C�.�NDs@�ɞ#��]�D"�!��x8�Ҧe�<閤��A��#m�S皠�8cM
cơ��Y�zzVs]��vf�p��ٯx��;nۢ�%x���LW��N���*ph�Z-MWt��/��sx?J������l��67A��;��H���C/�2�]�`�P�}rF�}��3��УO��=K��Y����y�d�?�\�2����'�� s��\�2���e.���K)��������$��#�?�ۑ��Q�@9�/ GG�� .l�)��W�P�86�������ZG�S���N�IH��"4�L����X��Rh��`䆐RD���U���D�����j����b�M�Ǟ$# �E�����J���j7mr��Ĩzӭ�  `�U��E��[�e���FE�KB[+�v:��v�}�6�X�_��λ�Tq����d�&�E([U�0��٢��E6�}Uc=�#���l��t�x�s�ckė�E$��0Ң]��4���a�(��W5�I�k�L"7��b�V�xL&C��Ĉf��P�D���׀"�1����ȥC R�'I��n��&���T�9D�J ���KU�C����S�{ *tg�`45��a���!�0v	�+B$9lP?<m�y�Nk��z$!_�@�T����b�6Gd6'��t��	t�j�`][���J#u�}L��3�m0�BjouA��v�nZ���*z�
fr+]��N^Rb~N���H��N �?����	w��&�~�,K_dH>���m����{�������߅�s�l����~C���n������K@�������	�(:��J��j@2��*�ȲU�`G�
�&��t���q��l{�9��;~ �>	 n:�תr�ОL#!y���䉐�s�MF�5l�1M��K���D-�IG���S���Z=��]�w�j�~fQ�Vvȣ�jց8.`�U�|}�zA��&P����1,�b����9���e��o7W�ֵ�B
�+��8��%z�+{b'Ơ�^|�HR�s�La��P�e�U�	[G�[������hYd�0
{ K���:
-�%�����jI�o6��v֋u\S4�]�N ���AK��Ǘ�#R�{n>���p^�>� �7M\O5��x����ɦ
��m��G;GRP�V	�{v��s��D|JJ&Q&g ��Ǵ�綳Ta ���v{������{�7�E؏��J߾��
����a�v�P�����(ٓ�m��&CӃ� ��F���}UG0���J:��c�������G�O�=uQg6:�v�4j���͙�#�ũ��������}��p�~ȳu�y����<�YD�	��NO�3u5��x��C��r��&k�����3�o,jt/��$��R/�jb����Œ~�t��&�Y��w�w��0I��l�M�	s����QRU�"2�ڝF{������Έ�g{�M�d�F5�����gg�>����j�aX>P~�@�3t�ó2��=�l�b�C��\�%;�b���}������t���1v8;󩃦̃�U��Ď������{�Mn��p�F�i{��]ڜC,%������sv�?V{�2~��c�Ustў�\�2��|��� 0���e.s��\���(���N��v���vs�>���]��5B��&a4$X$�����E�n�1��w9CRbĢ�4��*_G /�)_����^��l��/���eer >`�	 kH?�]P��gjx�~~#zŌxl����
f��h��t 	b�돎������m�\,�hő1dx-#��a�jF*�)
����\��#ή/.ՎH?z2�р90C��B��JJ����)��F���|em f,�*��\u"�ө��^� uPDZ3s��T
F�,�#�j��满���3 `z�XM^����d�ub 4��� `ap!�`6�κE�� /��~T�@H��~v�t!9�h� �U����L�N#� ��4���i>	E����	�
�N�v���u1�AV� � 8�nL�%�>%���L�&���b�t����������M�gUm���J�-��\���G9o�8�7�҅��X.���K��ݻw`}tL���\0)�%���[w�����_�/}�5899���(��H���Ǐ��?�~�w~:�Q� ��Xr�8��d�GsJ�>c��2����q�qC��4�;��	��Ufրv����m+�<��
��D�j�x�#�&�/u�\����O�]y?PֈQ��E:x�A�io��
�:�?��`�P-VZ��}���WE��GF��59]�m�A���1��g�>_�a$�z���z]�]�{��3T�|ۨ�c�, �f@w�$�-"��R]G���ͷ���#�Y�������~����SX�s§?�������~<�Ղ�pM����/�H�����<~����)>^l��o�	���mx�h���o����{P������s�ń�	2����� aI��r�y/�&��%�ȑ�GU9'`�c��sM�+��c�ӂ:42�Ċ�D.��rG�gg�N@��ͮ����f�n:���ah�N
S�#�P�F�o�4�������H�(yuu�k��z��m�=��N��q���������t ��5��C�e��)�
y���ʣ*aʱ��n��}����pu��P�s�7 ��Vd=t6Ɵ#�Z���i"z�)��D����",,��U6�~-��N��s�_���:R���h`�G�^��l�s��PL�{������P���]���)����q��
�c�"ϐ�{@8�����U�X�:�Q$eN1&r0⎒��5Ց>`�!�'9C����<���㖝�e|��n���B:�����y�ى,�_���N�����!�?Y�+�_��u���ut]6���e.s��)��\�2���e.s�����^{����;u�\J%���-5@��Y#�F�C����Q#F�N�-cT�b1T6��AQ�E#�C䥚8�x��m;�n�nz�������H�0L�;�{5c�Y��� 8���k�`�0���j�N0�+EQ j�B� 47����#���K�3_�
���{p��p4�!$���s�F��J��{r �ؘ	��wQc4�r��ɐ�9z��$ �(�fX�(N <_��bV��G�8��ݶ���G�U�Z�f�)�$�.�  )�e�,�z�w2
B��^HLg�*e����H&��p�&4M�%r5��(KUA!����,mOu�[��\:h�0m�Zߍ�2P��r�$O��6��5 S���_�t�`�>�OܗN��H�jϫ����VG�禡��bkt�]���N�k�0[UO�ژ_}�WP�t�aF2sY{��+	�p�Y�0����I��Ɛ�{
<h�kx6�W�q:3�SD��Q�32�����5���_.��C`��:�6]U��ݒ)��� ���V�E��F{�j�t��w�܅_hb���HW���{W��0��{d�D���DOo�/��蔣�q̃��mKAHJ��L��BU@�,2���oе���j H�[j�(ǎۋ��1��u�쓕��,�H��t<��9������ie�01Ҝ1k�0��s�X��O������Y ���%��$���=k(ئ�_�\y�:����TkdF�����*�3wq&�?W�B��O���)M�:�u"�3a��{�Vo�ݤ��V��܍�cOG8���=��U���L���� ���_�����{�
w��%���ǿ	GGG�������_��_o���n��ï�ʯ���|���[��D��k����_���hM��ګ��+/���߅�_y��/�2���G>�'��FQ��j��;�%۷��A��aul)�����r���2ϦA�T�}�A)��&�KԬJF���Va�pI��HY�&uigpy�8��u4��Ή�F����5��
g/������o��Ӱ��a��GgL���
���Y4'8E#2/)������n�������ޛ�Z�]�ak�s�o�WSWUE���$�&��&EqE�lKb$R~$�F����I����6ˈa�1'v`��c'�IY2EH�٦ؔ8w�͞��5t���w:{g�y�[E���gW�~��{�}�^{�u׷ַ�ù�A2��15���lln�|)�"(�"T����0��إ;��
�ĶV&& 9(z&���^���4$dp��b[��ʸ�8��sY�.CS���e����=7{{zpV���5!��]�J������Ֆ��P-J��ާ����;v�9+k��_i�DU�(�؆ಬl!�ͣv�]M43�w�@?�-,F�l=~/��Qi��DW�`�=+�,c�"N�̥��,%� h�%��KE1c����]�e�`f�"��/_�$��/2b�U��nӽ/K�����kOK�tYl�lA��ךT�P�U���І6���{� C�І6��mh�XC`v����i�=��@�= V$s,u�2ԅ�4�'k�O��q��g_4�������*�H������t�F�'VϸvyS0��U'�:KdR��e���S�k+0��]9�v�p�/�Z+��7kh�mȕS��e`[u�V2��mkkcxۃ��:OIm�Ƕ����?�y]`-Mt�.����έ�8ϣ����ф���Ħ�2Ҁk<�Jѱ)���I��rw�GK�X��|N �t>�,C�	�q�����������	��+�"cT.�)W�hf���)���NZ�<�դ�$��C��\�����x��~�\�
� lq �CB�|z+�(P+=p�깋��n�㎀ȵz��q��ٳk}��A:�n_SQ+���^����H��&�g��B�
0�A:���U}�X���V׷�n�2�w�����Tv��G�MHW���;G]aRur�\�s��U�s���О��z��`l������}���cT� ��۲����u�,+v�#� �E���ǌFc�����A�<_'��x<֭��A �llm}��/i=,����\�~���u�OK��d2���J`�YExj1f��,:�ӣ>��0�� *I��A=��Ie�稟[9K������I��F`����}�Lp��5z���M� .����滑 -�K�ǚ�!���D:YeL��Z��<���7F��&Ӻ��D� ���Z����erԀ������,��H����'�=��*}�+�R뱕�>�|���}����\�>�\S)���������Zʇdв���8��!�j��mZ�^��G��p�>����mo;<p����h��e����6�����h<���-
���e��^x�yx�O���}��e�ǿ��3p���0����g�	'N��O|����=
 �P�7��J�\TY�	��X�$��.@vif���&e���b��YU���GU�2� ]?�Ծ�M��f� V�q܍��\�C�
:M�G�g�� �r��|�[W���s��=��5XĉVz��&�~�G/�@�_�|�re<�Yo(h�dKk�3���ĉ�tdQ��)R�u��� �
 H� ����g�^�/���s߸z/\��g�A^�/�3HITUؘ�2�|�l|�7뵚�Ϋ6���u�b�<���ʢ�����#t>�퉁�,�F,�ak3�g����^�UL1&���L�g�k�s�O�[m�1����#@�2P�_e$y@����){�˗ȣ��=��ǃP�浔[��0�hQ�(����8 �J�i���4��`�	��ib5O�,��VAY�4P��G{A&��.rZ�F�Ac�i��2 �}�l��� ǆ��UU��z�zQmlT�'����}hC�Іv��! `hC�І6����i�6X.�9�&��9Q������k.ܹ��:J����tDA���HY|N�.�$)�b`�ɝ��L��HmŠف|�$�p)��Q����^����H��E�\�-�N�H蝓�z�����V����;�
�W:�����eT���HNYh[�ʘ���𯛧�#���� ��	e{b-���&;���1S3>�Qc�Itγs	����Yhݒ���Oܓ�t��qc�n�����wR�'�o^�B�� �iF������Z�P�$;_���b�c�c�e*�9ͩ��7$�ʯ+NX��Jr:�K���%�1*X"Aq�S��BVp��ѐܛ��y�^@��n������(*�Kr�>H�����xj�Pv^jfR%x���Kz7��zk��]9�{�h���{�����D� "���Qf�'g���
Tk��>�89�!�瑱�6���j�^�~�ˉ�\��1Ui ���#Y��f@�c�4���SЀ3�HI�Xg�.m�\��y&X����͝��l�ZB9  ս�p�ec�l9�4�}�����z10"�����8�!Tc����7��'y*�cmqw9@3��GK�MT80}���6�@9�����A�����E��|�OAP�nނ��.������2�K�U��`^��#���q�8�@���޷{������k�#��+�I9���	�G���/�&u��� �J4�ގF]L,�z�"��
a�>�Q;"��~���
 ���J���:O"���|N�pX�da��tM5��R���?�5��CX���`XJ ေ�0�D�{�
d{�͑l-����*���A��m��i����^����1��mG�eax��,N"�2w��Ú.�o=���G�lnLlMo� k�_�tn\}��B���u��0�ml��^�Xd�~ �z�2����K�,a�N`^���u���G`���M]�n����t,g����a�
�pj��qY����ݗ��2�� ��,A�e}c�pF��nI���eG`�&��yȒͯ6(~n�	��b��Ib+��S�u�s2�uѕ��"<�u��u�,K���1�X;���k���Ed'���r|C��M �/�h)� �h\�����5Z�8nKB�31���C�|��6����HS�E�ט�w�L\ ���q(��d{!��
��M�'�eyuTdb:�~��
�=��wљ-ڐm��4��E#d~�l�3��K�OQ��L$��w��{��ɵ��l�A�@&�%�Z
�b{�%���G̋�L`
M7+vwY�EF�q��"���V���੍)e9� U�AU�@U*��y
�d���?�����c�K�}_��c^�a� Yw����/F\���Fnf[/k�)�A�A��F�e�5���(z('����I�m��&���(�^P��HT���oɞ�q���Y��J%r�2Q��T�:2߹��y���6�T�9���A&�Dr^�S��(�e���r@-Q�e/H�22(�]�!Y��]M�mhC�=؆ ��mhC�І6�{���ڶe�C��)!}u�$���a�'�^�5��0���R� �5g�\�	���Ԩs�k�Q�5C��0��IJ��^��� LR�@�;[8[=�vԉ�N�[�=�w�?9 W{]��w�K�c�@���y�d>"���Fz�e�fr��;{��.LV��ކ�3۵vC5��vKF,�t/̖M�� ��n��'�����쬭���&P�f9���� �ڳ����z�~����?	��.^��o݂<���pF`ff�1XԑcڒM(  ��IDAT pq�)�C���gl�ܵM� �6��M�Uk�H�d>X�e�y	�3� $�Cej�����¬�U��׮�~��՝��/�s�����4�D%2��j)䪻�o���X�������M0�v�$�cF��O�n���u�R ������ѵޥ����C�AK�:�1�q5v �������%�>���H�T�dψ�@��];C�O��A�ϫȍ�*���M5 ��N熾|����%R�^���s)s��zH,c���,K�����0�.����=q���%�6��'�/�3��bP�g{k�J4���C��Q��GG�@�N�y�[�����o���x�%L @��;;ァ
��MǊ����\��l% Q/�]34�׃�@�D_{��Tk(0�D��{?��.�?�1�"1� ֙����'x���D����ࠞfT�8����I��C�d�lGP��{5�76�	�5����X�K�/����0`�7O��C�����G`�</�Z�� #,�P��S�N¹s����.\�~��f�(r�k �qV�a@�A����E\Ǟw����ol��h
�vB����>|�c�7�^}��qx��Ub�8<��Zþ`p���{�L>���;����{���ڕkp���vn\�J��Q�nܸ�Y�W����6t'��e_�Yt=׺I�"���ZSy��XI��$�=���ZYfA	��l:u���P� ʶ�j$��`�_�<��}���rY�/�M7��G�����Y��#X�����?�7/��|�}��7�u�lu�&-$,��;�쵖 S�ݨ�o��\�/ 
0E?���Q�gaD�}٠�N�w�d���&���XhZYb�Fy,O� ,fc%2�{�1��F;����߄�A3Y/}�y��ԍ(u>�Q�����,q�� un;�UF@����B�u�vIm�r�� ��Ӎ��@F* ]��׉ ��r�l^f`��wj���[�neh5v.���\�
N�Ok�>�zD���5<�?���'�g�!��'�w?��m��S�]]�
��\uQ� z^4��MU0�uά��N%s4`�˕� -u�I`�b�����{m�`0a	����J�.붖��#��8�c�=
�<�<��#E��P����O�1|���w���'
=�h�L��䲫�������!��RN`hC�І��҆ ��mhC�І6�{�eJ�jđ�9���ow�;���1���+�}�P�  �%q�F�2����r`��fi�5A`5��^_=QY2[ݑ���AţTӺS�|| N�>�^�n�j�`^y��mΘ�V9��9�A�x��t�������ѥ��\�y��ǔ���/��SOF�KL͊s6.�(V�I�\t���A%�iG����y����{�\{bېq~�\X#8�#��!)�<��5+�co�R& U��ܭ�+H�:"����T�_荗^ہ|�Ϩ �g:G�/D��5Ck���e��+��wߙ���p���wmL�{: ��L���Y
����C��<N%׫�)� /�P9�+w���&е�z@�J��սr�6>u�[�~�ȷ�{����X�r��U�Y��Ҽ��8�W�eyV��Ě���, �F�WzX=2�V�Y��
�A�Np� ��:+A������[�֚���|�,A2U@/H�uI(��Ey�Y?"{� W>-u�?��B|�t�.5���ב��	W�K\\�HO�\���,�(����7H���ZCz8�sf�9<���O�������=���ϴ�Ȝ:�-�5�8�4������ք�5P��o�Q�O������@��|�:�@�`��:��lӇ#`�T�L�z��Z�����T�`?<�2,e|* �[0�����>hk�����
3@�:��j�,{�6�N��T�Uԟ�5��Ϡא�'�t��KյM�h��y:S��O<O=�$��|�3��L�w��
�K¶���n�^Y+���[o�Iv9h����ࡇ����r�	l����ޠ�������3gi�a�P	�9��E��)��Z[+�?q�8�����|�⚻y�lmm�5���?˹d��=
`�>T��N���G8�W�Wd�����J/���P��p8s��
����X��^pP�N:]+�1�̨4d3���y�)�!-�!�!��Yl��ґ_�6�y�1���s�������_z>��8��ټ�m1�l�n� :��BGs�c����S�>�.1:٥��n'v��[0�?��vvO��Z
n�H΂K���e����2�c��$�禆������B�>y�-2�(B�NA�����Ev�l�h�r,p皡�y1��7cYw}-[�a�YB6a���\�}ŕ6�H���Y�pR�EG� l�&�k���� 등>}7#3���q �k�Mƾ�|^�e����Ynmo�Ws��?��a������O}^��jy�r�Qی(DmY�|��Ls@��� �%�0G��_�)�ͯc��T��z|�?)WpPǎ\�˳�,������(\�q�?�0�����S��o}Sغ�owb�7�}�'y��>�c���Q`=[�6�n���І6���{� C�І6��mh�X����~��}RZ�-�u6
X�����H�7��e
Bq��%�Ѡ5��ټ�8悁I�5�.�=�gx9tgh&�\?�&������[����*���6#��(��}�v����諻�@�a���̙~���i���th�QC���Ǐ�r>��o�Gә�A�ߥ9���&��1�)��Ս�f-]{c}������5�>~&�

���@f�&e1bm��R�v�9�؞/��� �]g������EvȕW��j�n:��R�|5��y�r={�ث�Us5�>�R������X�{�_}q
�}S����sү�j�	�$V�e�	��a?���NX���#T{���!+Ӏj��\��d�����K�V�G���J=�a�/���+�X��m����J���wu��N�;5��i�b��#8W�T�t^Y�, I r��)W�z"��˃�c��2V��ܩnhy�L�n�F��z�����q[�J'�]��
1�-Y����]��^/�jA���D�R1Q���JO;U\���=Y�K�e1�o���CX�a���H}�2}?�k����{�
KC�Q����`DCz����upP�0g	�H���ن˙�@��Y�8��g~�����<?��u��Aͨ�סmM�2��I���	jhG-[���;�@5#��(����Nu�i�dC_��1�=PoU�U�8R]�H)�d�ۛ��f�(�������U:�n���u��yԱР�ﴄ����ƵkW	�Gp)�}�;�'�(�eu��l���޿�Y��������y��}F`u���Nh7lmoQy��7oR����(��\	0 �v��d2��ϵ���4���#���,�2d_` �XJ��˶�������I`j�&�^�z�6
ca��E���b����"�Z����p �� ��D�t�t�غZ�J�MFU63�wԟ��%������o?o]x�8w�7��2dE��#'�×���ex���X&�����h�%a0
�����6�G�=�G�eMb2��H�C v��"���"fȑ�B��Ө{0p� �7$�8�y&�7o೿�y��N�}���~�`}R�[���(χE�M��٪�����׌zӧx�`e��=�q�]�l���s%3��;�Sr0 <8�����yj2��Ym�� �L��;�>�Q�E�ҙJ��ԃ{Au�G���
b����{_0��f��tlu�Z��lH�zՅt�h�CAub�K��k"��a_v ��u�����uA�ߠk�m8ԯ��Ǖmh��3�d<��G=@��c����6:�ǆ��ҋ/�xk^|�E
ĺ��Ix���6^/�w%X�?[�6�K}},=
!�hxW�[��І6���mC �І6��mhCڽӐ�_=��9��Z,63�����R0���������H�Q��IK�
��Q�V ��a��R�_>�k
Wv��m�9�����e~�MW�����?r�� s�=��$w��O��a����,�>w���z��_��|>�Q�G��7��}���t6%�J�շ����"g�"�hҒ��-�Q����76`<Y#�l�`�F2��1��rT�7s]X� �>�ʵ@¬\���$�*O,�����e�b`�2�NmR�2�k��~q��+���f�>ёm(U(ؚ0����*�Z�*�A�2T}��I=X>^B]W�W3�ep�����.st�g�����4՗�{�]��U�߰�$7�:�d��l�|�+t�U�lpyW*gS'*��_宵gul��b�tG��s�x[wY��-@BAi*�"2K������Y�����z���lNo��=���WG����zQqs�=dwVkb��� *������;d�1=SAZ�������y��l�q�a:Zw���TS^h��%������XI���pp0� � {�ғ�&�t�h�}��2��n<s��.q�t�tIf�)���f\�l�	U@��+�-�����3�Az/�/|�>���'�z����Q��,؄�:�m4,UA��(r�x @�&�[ϥP�7\���/���k�Arc��̲�3{�R)�~%]L��W�3{�� ���3Wp �N�[3:�+��䪔�[��t��j[C�n(��sݢ*�߱3���v�J���	=�l�(�S��#���,�7�s8�9�kܺu67����FY?��b��������f_c���p��@�۷�a1��({b}L2��Ec�r�
�����������=Д���
�/kK�=Nק�()���j`��j�}��?�w �t��"D�O�S@>8M:*s�y�yb��d� ��l�C��-K:s���S$� ��hxwj��&X�q`� r\�Z���o^��{��~�ux�S$ۇl���ۅ윇�����_�����f0�T^���Or��5���Aё�ɏ�G����l�ҡ��mOd�����g�񱁃A��}��ݢ��D6�q�7�b�$2�1���m���,��	�����uXs���7o��y�n�Xq|����B{����K���F[Q:��{�� �vp v�{�����Y�HK	�.��>S[>f��5�_�9X^8�Ĕuv�$�����6|� ����U��A��M>NA��j ��\�F`��*�6ԟ�\��,��2�kJ?-�LK�5v��Y8<:,v�>1Qd{�����}odnW��������We���v+ W�s��β_��K��1�v�*|�_/��������G~�C��/>mvA$��� ���@�}�1�<�l9p;U��'�>\��H1���hC�о�� 0��mhC�Іvo�BH!���V���0<��Ԕ�b�i����Z���9&�iJ���Y���6X]���M�$C4wB� �d�@�,�3�P�\�]Rws��%W�zL�i'�Y�+@���/���W��sԎ��u�a�����������}gD���/%k�!'�r�Am#t�t^K΢������&��>'N� � ��)���ExN�Ns�:K�.Ft�Y� i�D���P�;m�<
";���C���9�`�C���U�R�PtF�-�Pd��V��ʊִ&�F�T�Ik�Sw��}��+9�U���P������I��ªL�3i�m�L9�,�X)H�+�,���9v`)a��f�3���z���_�*��n>�*�&���ܜɕ䙳/]}VV{-�Z������s6��q1Wk=��� ������R�@�mr�0_��J��S}g-��){�ࢂ���K� �fq�px>��~F	Ω�
��j���-��T ��AH�]�����G�G��>��p�)KR~f���cQ��ف[{{�������{�Ex��	T�ۯ��8y��+��)B���T3�GG2����e���I�8�^ٳ�>���	Ȫ��\_�8�*���LXH�ٯ��&����m��U��ڸ�PPB5�>r���t�)DOU�d.B�טō�/�/2�������rq�&f�c�l�8ำ��,��%a��y,9(��9��nꪚ�1�s��w`M�jz���e=)�j�م����6�m��/��K`�w=.:-����NV6ȁS,�&�d��s�Y�+�ă<��[�@=�@*{���Td�!��l�%�5ؒ��w�Q^p�q�����{�0�e�
P�e�:s�~��+��Nς�?��ۿ}�O��Vq���eݽ	?|��G?�q�g��x�;�+_��<�큳��q��^��D�ҳF_7����g�l(��8%پ"_I�bK���.3�@�ۦ<�jk�����#UN�2#4�s�V~&�@9�� �Z15���GW��dk������)8Xb��|z��_�>�P�E����g�g��=�,<���S0-�Ǣ_sCz�C� ����l�d����t�Z	�P��Ae�;FJ�D ����=^��2{�db��f)�K$֍�q@�m�v���/��7pO����ƚ+E[(W�����n^��;'!�q[J�%�SdD@���>Y[c�Xbq���<�n�
��{j�鞩6�~���2�jb6}�}��:��.z��!E�Ⱦj7� U��C�z�λ�j�E>��M
Ig;�ohɚ�5(̟��n�s ,�QY�Q��q�����V���_�-�ې�Tf��{��ai�Qه�;{�n�"6�����?�~A�������R��Ե��[�B������Qw��ؤ@��*���Y�Zn���ue�Í7/K�����ˢ�e~e>�;�JJ��t����ӄ(��Cs��t\� �(��7$�!x|Ӫ=��mhC�G� 0��mhC�Іv����գ��
�E��;f@W��\���q���Jǿ��*g�8\4R�u,���|�wx(<�Y�����e��������ߣ�.4����.��=g5+��]�_�,{���߽o:�Q�S�:��~>����.,gs�kD	��H���f�F�U͠	����$B��!��	���ѡ������H���s�w�~��˝9���9��F�m�Mi�.�S�3�Ͼ\�`OT9��i��ڹ*��E&�
v�o�Y��[�8$�Mu�if�_�o�͘�D������2����F�`R��:H��I�a��;e)�w69ƃy��j�<�F������d[��9V�_�c5�n��l+2˘J&W ń��4w�;�k厕��J�l�-3�ܜ��
�.�0�� �<�6
��a|s'5S��0ӺvL���r��ݗ�� ��o׾����Vj�T�^�.'�c��9�Es);��s�������0�lx�``����~Rs�dA�ct�MG�3z�_���d���� '
"@�z�y����3�Z��q�q� -)��|�{݉�z�;;;��r������Jb������ϯ����cP]��T��$@_��^��
���rF3�S���W���d���2干�%����N;ba@*k�r׌~�dNt_d�
�(�A4y� Fa,�vE|�"��T�ꕪ���[��w6�(7]=p��.7ߏ��n�){��!�h���<��QFp��OtQ�Lm1�T�155�i���(���9(�Ȫ���p���N��){�r)UUF=�?����t�E�c���������+��򥷨����o��/�H��=gv4����p��}Ў#�̿�����e�Ύ`��!�����g���[p��X��ܹsp��=�LJ��?���un��B�����eφZ	�
�㵖��Q�@U��M	��Β�GG'�B%��G�X۾�㈂#�hSu�F�
WU鼎7X�� /���?����l�蟁�b��P�b9�3��-��s蚲;8۲��
�a����2֯��<|��?	�"'����aܖ���#�sb����7��-1s��}H!�|H��c�z�l@}��������&`Y "� �0��)ln�7.\�_���=�v8hO��>�ؓȐ�O``��ܸu��SX�X'�%ʑ�$Ʌg�E�KS��<�Qt�˂[!���_��X� {��"�U�_}���Z���4�~K��E�^ն��"Q�ϭK?'ª��	�M��z��P�~!����ސug_A��v�2Ǥ�g�n��_�Z�fb�:�J~p �x
�@�: 1�ln�9-���a6=��},wr�
�Gh	 4�ʎ2d���4��xG������:��P���,�K�5��U-�g��3��ҧ�,�!3ڬ��ܶ`�KI�{��u�/��K1����rD��j߿ÝF�І6���^oC �І6��mhC�=�ʗ|b Oz6�l �RO9mXF$gfgv�Wg����q0��A�&=�B�� �+H ����8��>ssz��r=.$#�]��yo ��度H>��I;�r� ���x����W����j�?zr��879{r��
j*��= ;�0�k�4� ����X���!��o@��!��I;�����,l8����F
X��$�X<3�	����!�ȹ� \G�\vw�3�6y��g݂��vK���cU�u^i��5�x(���xb�
`@��!��+�Y��/y�>�=V�.�u�������t�����enbq��,�<���9��6g�y��5=UЍ(do=��dMM_�\�T9�]�t����=C��c��&4�i�|�Ѭ�s�S6
�~���ߧ�z��^��u���/�%���~�ܓ�z����lk>��C��	թ�Լ}��y�����Lzs��>9�	@���hsd��@������~'�yHٲ��8}-��k"�V�*�K������%���-�L֚`�z��`���-���~?�7[���#�X3���?�8�%Sfc&�!ꔛ����=�?��NZ�r�ѮM�,�	�1P��w���<�\�|�lw_��ДܞF��k.��>b�?�L���ճ�J����T� �I�$�Ph&�����P'g˞F��m��7H��X����V`���PhS ���I��*�,�D&�WJ�q*�;�� ���Z��R��.������*X�7�x� M��Ze:s~+�� iЄ2~�
C�5��c�3�ܸq.\�P��c0���x�}sf׉�����aI���z��D�X��fT2h/��*|�?���'����?���_����Ϳ���·��<Δk"��/���0<��y8}�,���?	W�]�����/��	^z�%���a<�׾���t�"�FS�.�tU)g��#���71='���'�z��"($������Rs}�۬�Ȭ�.B���(ۋE���!����d/��Q�i���p��������?�W�)�=� <��'�fהq�hfeb}�EY+�'b��`V~���6�B��e>��Kp&��S�>�"��2Q@m����ƣr��/�B=���8F�K;)����>�-fT
e})z����ʻda+�>�܅�_� ���~.ߜ�Ɖw�x�?v
��:C��#�9G֑��;��6������*�8s�tla�Rd[�ڕ+p��iHX&�� 	d�� �����*�����ge?3S0�.ۿ�7�5�bf��^�a�P�g6r�Ù����f)QA�_����r�*�#.e�0��!VOU�c��f��m#��&6�]��m�*�2��dש�o���k���v'������Y�-��@;bzt��N�AǑY�(�+����;�ˋ~w�v��xf�������9@��֒��I�G��Y,��D9�te�E��,d������W����1����{љ$�~��w��5��mhC��� 0��mhC�Іvo4C��I1��3��N�ui�R窀9�Rǽ�wzYW�S��0qB��L?3Pל$_ΑW)����什���0 M]Ɩ�g���KxQ�����W9�܁U9�l<V����j���հ�ՠ����\}]'T#�N��	HC�`sk��*LgG��	�d�߆�@[���\/�C#t���1e#b��x8 ����N������T�sqL�v��2S#�%��Z[����O��[���7oS	t\�z� ��2\���f؃;��qAre����sv���j�B�* �g�9��9���M����.��к�Ii�@u�X8QZk�X��V�=��d,�J>9Tzm��m�9�<�<��de{@�:��S`�9p������Y�B_vu�2��~kw*�����,"�+;�Q(��{zW-�P���(�='PI�!8����oca�ׁ3��Q��$"쮠�l׫=ɣR���0�f?G�8����5Pfe-u�f�z��jh��3��Qc̱��$);��}��0���ͨ�.K�0nG���H�t�,�	�Gs8��4��f�5K�79������}~xxH��;�� ���*��\�D~wB�^1�ܼy�n�����\YY �J�?����3�´��d۩՚����ٸ���00���e0�_�G�H饶6�8�4�i	sd;0?IFeƹ���x#pK��0E2��($f`�"����P��t@��1���Jdyv����e\EY_j�W+ޠAC��j�Q�,
z����!��{)��?�g�# �Ҋ� ��spp _������h����z��=20��rYdy�$[�9Nf�b9 ��/�����7����$�F���w����o�zĠT+�����������~��0B�����GG0��#=��7��0e=v�#Z���љ���}��\��ٳ�D��������Co��4{�#��\C�j���&���3p������؆�d���΃�B���2�4�@�������UHӷ`��	x���E��:��q�o��u�/X� ���זuL�U��|7�~^�����Q:	W^ڇ�<|j�>��Ü�NG�q�e%b�"��r���֐v�J� �k.��0�e6[���=�>�\?*Ͼy?�x��09v��!�i����
���tWCS���������o��.�����p���K��ٳ����V���Z�����J<�7���lKh,��X$D��mxO����2Y�\L�6l`[ j��B-�)���+WU��r5��#��fs�\KJuI��c6��b�$ݫ4("T�beh-6*��Nr�ucP��w�Jj�8�[M���Ƅv4��F�>3�?B���5�ȫ��I����J��j�t��/�A�Ez�U���|(�E�!�Mb���O.#B�����b���)��`�\zP�t�J]�MlA`�u?Uم�mhC��b �6��mhC���&��L,���B���vlU�k;@FN���Z���&��:�%�n��g3j�(A5
�8%�|_�����[S���� 4�Au��5/	�+�D�QN����?�:��;�{�[�R�3�=�>/��!��ハ�8�v�O:D���Q8��	L�R�	A6�#m,�3��l[<�]�h�e*�,c�u���0G6������=x�T�6����%�Q��H�z��I��p��5�/3ܼ�O`f$*�e�>^Xe�W��	ACF�S9'*��A�\�T�b�}� Vfgf;q63;���1p&�$a��%�	�@�D�:SI���OP���U'�4�]��3x�Ȣg��Z%�ɫ(2���<�l2�4� N���V�L���A�V3]�oCS���$�#1p������D��eWy) ��d��=��*�T�C�K�Da�f���@#�͛>��]����͑�Ϝ�"� �΁�@M Z��+�
d���qba�Z�d�.�у+�`���7�<NN�˲��L�����L�he`�jge�5$�/�B��A�)0P��Q��<�������>��_��!�~
P�u�.Y�!g�Z����8�oD��x�����}K���7�������K�Q����z9��,f̜F����ٌj�O��{{7���K/�/��
5?q\���n��PF��B=-�5��A&e����LZR9LIuY�8�R #C@���H� f5He���9�氹�&���V���/�oD�JL�0�{�8��x�c�#�o1�,+���k��Á�$R֣�:g:���dS��_R�(��{9�S͵�jl�,�%[? ���.��z����j;���>nD75j���5[6x���top����rF������`����-pO�8�:wQ���Q�oo\�_���/�l~X�qn�:�!�L�ưV�Ԭ���_}�e]�u���ֵ�t]b�(k��B��^z������4��:��>bм�Ù�%
�:	@�`)���Lw�(�~���z�'����F �D��Ӆ'�wtyf�����=DupG{��Pd��p�aV�R��<�
kׯ�[o|����C^L�`3��`q��p�]8u�;�����v�E^�9��8s�O(�U[棛.��w>^��-��ge��G�VzB�`�A�
��h'���� ZTX> n�|���<������x�C���w�Ƕ6˼M)��cE[ƿ!�q�g���ҕr�x~��?�˛0�}L?س(�r}�6��+���[p�ʴ\g�g����Nñ�4�I'%���qA{@&9iXc�Z/�}�A����W�����V�SPK��bRtUW�����`��I
(C+#���F�f�x��}�e��zb�ʢ3@*~x bb&+�ge��;EfR!��� / E�Cjd�'�ijK�e��T�u,�WѾS}��(�M�G������*���L��#��}��1��U�%�u0C}��"����.W6`(j;�n�:�K��ގPC딀�䶧�|<o)���a�9�ۜ�˦��@״�T�D�vfò RJ�ln|��1�	�0���7������Lf�[ `V)�j���9Tb�kك�ϴ�J�j| ;R���w���,@֓�s6�3�vFG5�7�̦�6��mh�Cm �І6��mhC��Z��_	`��.��V� ��A1�H�b�2�����#�:)�N;8�G�<
��CK3k�鑫��8�k7�!����?����S�lg�UJ?����W���q��u�8S<�� �~�
�덭��%T{���g���]��2�F����p��UX�Q��:�JW�BO�h<��c;p��i��ށ���`kk��!�,f��چ��8�?��
���Ɏ��lNY{{�`onܸA��z�
\)?����g{T_���K*#�5�A�1��^���:�` b�0���!g�V@� a
)�΀��:4�A
������a��Ͱ���"��ď̜C��)㈎��&�:��*K �`�Af�|��>jlf)9B(���rn��if� X�XW$Gfd��bk8۩�ck�C�`t���Kǻ�u�lR���S�tPt��s�Sf�x�1ŷѱ���0v$F�t@
����U�ѓ%;�{)�$��r�R��u�D��u���/`��6ˎ3+�8�i��ة|�w�S�kUe��C��B�
�0٠�5J�,0���0`�=b��kH"2��/h0�Z�L�t�����U8P��l>%g9a�[8yj��9=��d/�P嬅��n5+�f�S�@����?�u����C�8_H'� 2VّQ������"V��<�Ʒ����Rh<��e���	P�`_y6����yP�e�!�?@f��:٪��Fw�@�Ƚ�I��9E��u*�ǯM�D!�D� �W0׭�!K �gbF��1���]��tR�Bk�@��#&L�c��!��L��T���X�0�3�X�n�����@����*�Ҵ"�XT���vAo&AS1:�5ȣju,Ŕ���}��ɓ��3ϔ}z
�/����gioG0kZ��۷o���>\�qn޼Q��#�/f�÷x����#]q{~��C�;�Ġ�Z�~g��J�z�A^��̒�m����ඒ�@,�g
j����~O<��Q��V�fqʎ�	L2k�i[���������^�ٵ� �/}��kp9tum�8�RZ_[#ݶ}�lnX[\��Y����./x=d��b�]�px������8���9��u�w�J.p���f�j�KM�$��=ʲ\�k�{ ^�sx㛷��kc�+}��&U�_���e�� ��$���-���q�z0���5�׼蜫7��ҍ���߁KWo��C�>�a�3��s�'-��er���2�m�F!
 �6���p���s�`wc^}�98���pT���֨�T(�or����0�)7�c�����!�<W�Vdv8�k�E�5�NeF�W�,���}�ߣ(���X��43<������jPFD.�E+���5�)�q[��#��D�'bá���l^ԟ�Jr��L&X�܀��1�#
&IK�״����#Xt���\Kwa� ��e�xOӬ�GS� �}^Uʎ@�.�w�l�����ը�Gm"��@eC X���Sy��bc�G�z��J1`�m�O���Qh�>V�`�d���Q���Zj-Z��0�噪�U6Np١�iH��(�������)@�礊yIyf�`[�]��e���W�6��mh�m �І6��mhC��Z�����6p�Ўv�v��Q@��Jى#�cP�X���sS0 PKT���Ռ�������CÜl��X ��d}��K�w,N���*PI�?�}2䠝3狎��u(�jYd�a�c�>��z���:S)�d}�;��r��C�2����M���[����`cs������S�(���}g�{���Z۷�������`����p
��o��7�߇$�/��1���*� �H{�l �rk-�����̑ZX䠓�QG6��D��q�q��!Z9ٹ%T
ȉ3�3̓�X�,��PPG<T���Q�)9��=1C.��Tq�xD�]|�1e"�F[��d����Z6s+@��Ҧl�Ƞ(g6qf'g�I�3dų��B"9:c�� �p������`�H�/G�c��sS��4�U`P�Lo]���s;rnNgGD5}xxTd얀8Kkp���kk0�Z���+l��lkT�͜�2n,;��s�`��X���5@+I6�d��<P�dh�����f˵�	Sd#ю�ߒ�(������TO�@�	�<T�vgs�S��lz+� k�K<�Lm�:Q?�����M���\��f������la����߳yY�H!-�eՃf�z�p�����T���"�ٝ��%I]_|g��d�s��J��s R��	�60��.�n�x���"�m��YG�ס
ܩ�W�gt{�lf�i�����zfai�5�t�� z!�H�g�g���%��t�@��/ζL�8�TK�XX0�l2�P�J.�X(�dEj�g#
X\��:Q����
Q�R��ײo���E׋p�8f�,g��;Nko�Hw���S�W r}����	
PCu^��T��6U��ع��Ho�ވ�HǏv��:��y�W�=J�`��_������t0�v�U��8
�`$�7�ʣ�{��DS69);��j6�t��%��� jVUh�GFo㲡Cmq%��&��=��6D65*��*�fW��k��'H!^>i���ė�ݿ��#��>a�7�n�W��5����~����Z[���Ÿ���/�M�еdf(��#��Gֆw��I���0do���uHQ ĝAj0�3��,���;K<?����!{f�/˵��3�K�uhۅ3�}��Q���nR���)f�w0�i��O����b����n�������S��q&���#'�jХZvuÈ�?r �Yiɤ����O*_%]���O�����~�w�ч�����Z��e[�<�x�A�:�>�=�H�䥓�4}�r�RWp9T�Iٲz��ږbu�E1��`���f�k,xAk`�3��\q�k#e[Ц�M��}l~���'�x�;s�2�lǵ����^�/�����~��9ֽg��q�^�D'A�P�gL����?��w�����P�F;�M@�v��/^������?��-^Il��	ˁV�k	Ў�{p�B=D��A�2b�$D�=;�Ñ���r�|���0U ��%��6�u�)앱;�E��%ؗ�D��XV�!������}&�]K��3�^��w�ئ2��s^X�����v�LO�3X@�{�.۳Â�WwwfOP��>׿���ZpC�І6�{� C�І6��mh�XC@A	���#%��	���a������ǚ{k jO��M6ϵf��s6�D/����o�� ��=$�����n��{]9⠑l=e��F-s3T���ft��U�*K���� �='�wu��޹=�C�
va�̩���0�M����2{�����:��#�3��a�:˸��M�ҧ�,��8�k�{�,l��7�L%�jR�_X��><�㞤�1:)J�rt(rY�z�#����L}~����ăf:�~pkb#��@{K���
����?��p��q8q�$lmn�x2&Gk#c�T�q�� s~W�N2��0;+E����O�̚!@�w:6�X'��8b��usgucg/�;�}�~>�Y���8�T���0*  f��<"�[ޛM����?��_&,����4��H�ʗ�'N������Ic���:�QǙ�CiŃ ƚ�F���˄�Y*�*8�2r�0�'jj`F�ލ�n�]<�N��:��Z���(P��l&�=j_�-�KF\qȞ'��UR��躪��9�9�8t�d�3�d��+ }�yȵ	���I�ݨ�=^\��5����[���$��TD�iܑ�9[9XL\ݔ�G��<H,kK�$��R���{��S�˄�D�lF�V�5߰n�r8�D]�/u��+p�����P���Y�����[�P]#h�U���M� &��9͗�,	�>��}�� ˸]'%�ǐ�,���1_.�� �Cb}����o���`��d�@)��jtCb .I�I��x�5�-�{v���q�����x��R�u���ƾ�c�پ�c ���2�Ve"�w���o]�܂����ye9���S-LZ[���*[H��x�L����X,9�<+h��ڙ3�ʒ�j��)��jR�u5_rfq�K�3yQ[��K��Q?/�g�VJE�U
���gswBЇ0��N�%:3@�_�A�{��|9��L�@V6Gf���-�\j�@��冞������ix��H�Qq'x ���3�?�qh�3�Ϙ���NlN�C�k e7�Ne"}�R�qE���C�R\f4*��뼋��r�p���n�Gh�! [�dR�Y�Sd��[Eq@S�����Q��Q3��$($usa�1(3�sP ���Œ�K����ϖ�DY�U��f�A@���8��O��>�#?
/>�,,.�	��<e�g�vكq?=�C�����$sMƂ��=j�j����e�˦ws�c����(��T��}� ��@ɶ2o��s�5�D��QoM�c�/����z�Iz�@��A��Z�ps�<x�!��~���%\�p��?����ߦ��b	�"�d{�������W��_��`Y�~`I��۹F}�~�%�?t~�?��p�S?�W�6\�|	��})��A�4�{eCA���qك�c�Of�%=��`(��Z��.�0 T�� �X�]��d�j��>�i��L�)1��n�D��:BZ���D�0;�R6��W}�mU�*W���V&s~��1cAm�v���w��C��w���S�#�߃� F	�L�mhC�о'� 0��mhC�Іv5,2�g�=Pޝ�� u�* +�u��wp��a=��>��'�NVݑ�lwX� �?�rķ���a�Ŕ*gN���ΘU�_|�Gv���ι�>����ɝ��d�@3�֝V]�_��ݪr������w�7";�03��^�7n�4�B���/�f��E�'�0�_}6�s�U��
��F%0��4�B�Y9����4�>9�_2�QBh��j�y���Q3��xB�b�i<4W�gk�x�V�%'erz���=�agg>��O���c0E�ު�׌ Ơ����ܱG	|�W�a��&�9*������yf
�����(�W=y�H�K t�վ�x�:P�0�k��c�C�9��e���`�R&�8"��wz����p�&��#��/��/��@4�6g�kű��u�rE�+�e��	r�VeP���0��|t�g����g����c)���~�_��2V�����0�؏�8�8y��}cm���xb��a�J�3�]V�ޡxU��賵��	f����t��`Fu���O�W^���ϒIM2�z�*\�D�Z�_*���(�",/`����y@�8�����Y��h�fxP��m��������1-5�?�S<�R��;�z�]ƿ�	�,�>KA�{���}�uS��QRA�N���O���F���Hpa�`�L�KG%�,�G�k
��9��I̦��ِ����ڀ��n ������Hh��lC�:�1Qv�j���m/�1� C�uM��T�Pu"�EA�c팬,@p*U3dg�PpD�+�)�67��vVݟV�|� ����^� 5�aU0R�{v��B�����Z�"&�w���\K�&�����aۙ�'
+�g&���A8g��n�Mj�I�cr�k�e�4T:M��u6�ko� *a�N/⓱y����t��/1(I�?>�/1�Gp��9�_½�������E:d�ǲ,)m�V0D�,3F�ߍ�� �s����A�$����jk��h�)�\j�j�/(hg�L@l�\��~G5�#���^3;0,���ë��%$���>g�����	 �Y��2�� n�
���R����+��
�~�[��C��ƱX��]���oL`��d���m�`���st��xj�a����4X�"��b� d	m�����mON��6&�7E8}�$��/��p��9����bGM�E�d'QpD�� ���ٳ��9�����{����<�H� s��?�'��1l#�EM�[2�*�����L���"w�'������߂�.�iu,���V����$|�c�x��61X��k�>�q�|��_�o}�[F�����*H�oV����G^������7pi��-��H�%���h�`���(��w�4�^���n*l��%\%�X9 ��)����l��u�����E�4�
�3����DwV%�t[�O�Hv1WQ�C�І6��6 mhC�І6���c�bu��(N�J΂^F�f��;�Yk���\�������W��	��Sj���,N���ݚ��@�[B�#(��ߥ�6�{��{���TQ�P��V?�C�Y��9���nC����t���
rRv�'b6�hĴ�~�c�>ؠk��;�|OVIR��ɹF��!m�^��Y�=ǝ�
�h��:�b��@qz�؏��@���3/�q���Q�A�z�N2^�<1�������t���0��NJD�R:~��-O֎ư6���%���'Ĕ&�h��4�L>�
�+ �`��>�<� јD�j���E:�Y���;ET�)#k�n�Au�ژ��:`�`���z6�;�eKYk���nh�,: �=�A(d�����:�on�����g�A���E-��`D�(�l�HC��U@Z��JuR�# ���7oޤ�?O=����O�����E�g$ɴ@:YMٽ�Ո�SX���5?��X?�ÏϺ�p�&.�ώA�}���o\� i�Ϣ}1�.{���VE@�J���en�n�v�>��F�^�"��	�:B3�c���sR�� ���ʘ�J&f��I� |�첔�6��W� �;�̈́ҤJ��d��]��Xa��^��*�1����R������Y�� �w�"ޮ�F�4��	y$ɲP�km�Tƿ�A7PS�.����ub�hTg���k�����j��Uo��`���0���.e Ԗ ��_z_Փ~SePۨ.�`��U� 2o��Ax���zc�ǧ������:�Y��A*��K�U/�Cp��D�'��t��n� -a�׾�\���:E���c'�L�_�)�����X-�:9ԗ3�i����%��r��vf�k�lcG c,�� ��vD��S����}im\�,"��_��p�ڟc%�Oi����®��g�<I��Ӹ�J?��������E���aıj$x$�
@E�hyGe�ms�m�t+4�&��@lJ�^�e� -3��?I�}݃�a۟e�u�Sy�3���&x��_���a��Lƛ�@�U�zz� &x���#�L�yksc{h�HX��t��#,@���>��f�#�5� jօT�)H���3��fV�l�,FM�'Ϟ=���;�����������_|����W^� ����{��bg<�k���T�?�����_|�]�Jv)N������쫲�`�������0=:�=��������}��ԓ�M_~֊�����������-y?h�c���ܿ�s�O}�������Z*cq��9�}����/�ѯ��p��u
*�rIt�k�U�춝�PY�d'�O��a�Ւ~?q˨�UU�0QZ1���/m���;" ���٤6�HP佋cܢق*�l��x�*��Z�J(�3�zv����#% / Z}]���І6��}�! `hC�І6���jTO��K�ߑ-��y�r��&��ݹ��lԹ��骎dqu$�:M�o��t��=�����
\��5�@?��S�W@��x���"���vHeq��_��{�s����9�����[V�:Z�n�׶�:7%�.7�FV�/��[�I5&�٘�g��Gɮ��j�gj�%�݁$�}�5h�c�@ 9D�hN�F��+�A���&�t 
T��ž-9R)���8����{J�,�y�UDQ ��%����6��D�e��2Ms�,ͺ��t0i�S�!pנf�{E��c�/hvЫs��Ɩ�Ou^g�A޺,���k�Xn|�ޚ'u��8i{�K�|z��K7P�xdn(c��A�A���I!i�pu]��]��#� ��D�Rkı���g�FC, �w�NIH֣�?�,���@�k���,���l�VtB��x��/t=8:$<�L(hq�V�Ri��غ0��ϯ��4�E_���Tg��c?�尃�|Y�l�aR�dM7#��t�D��eLA@.j�jvП���Y�:���f�;_�Z\�r5+/�67�Y����.(��^d${+Q�V��p�#���`z
;g�v}� ��������W���t�
nր�?LNYg����#0�93�2A3X&��t�/e��F�x�}O�������^#�5sR�D��O_��Ж5��Rt�f�F+�ӈ~RZ{bU����I(�«�;(Mz5^�r,P��@��+�S+e�OE�=���G��Ad�uc�~R		���+��'{l�"�ާ3�9H�h_��K<��|���&�SX��u�m� ��,Z��태�@�3�֔�'t'Y1V����Ft��wE�SRt	�K�Ҡz9U3�z�oպL:vb `�N�չ��%����Y��XZK�֧���\�x	����!�J҇��C�9/�1��kQm<�.�$A�A�Ĥ�\���Qc6�~�h;5�w�v\�e ��i�I�P'��4$&���x�Z$�#���B�|�`�Xmc(�����Q��NfCf�=�U_�8,���50	|WbB�r����'��٧� {�]�3<��1X��2���� �圍��
^��I,�i�|�ޒ�ݏվA���P��f�+@�]�� T����ĥ}G�0��Iq������_��_�@{r��^z�E�տ�w�������._�g��U����m��O�����¨���@�ž�s�?���������y��$΍�7�o�����"�u�E�ї/����W�#�}~��~��Ɍd��1��������H�ۼ(�?�c?
?���>G�v#�lZ[/�@�[p�����O>Ul�m��~�s q���JEi0��d��3C��x�uX�`��]�IGP�͑K�ЛK�̾tbgk� �t-rI��P��*<"GV�I�z�N��Z:c���/�w0��)z��W}F^!HS�+��mhC��H �6��mhC��������LEv&0�z��+��%EgU.���dܫ�C���t!G�֧����;�ѩQ;��T$�r�!S](��?:���]/We�U࿝'�X�X�*,�4(0�L����%�:rru4��鏗X}q�OuV�;y�)D��r^��/�Ϛ���cM4��F���F��b����*��|n�L2fr�7��c1�Ik��C\��v�7�Emp^���cg�o�N�ɌWj� ����ڪkX_[}��w����>Lg3��cp[d�yE?僧�!͊�ω��16~v+�)cL���L�q'���������f�l��d���` Q��&7YS����+@] �Y��8�{�o5��/�ֿm	t�`��S:�%��I�l0�|�Z�-�O68���?{o�[rՉ��{�������ҫZB�ju��f-����/1�28������q8<c;bb�c�p`�aL�I4ڛ�w��~�VU��o�7�y����c���������d�<���~�wʒ�SZN�(^$u	�"�E�]g�H1����xQ-P��d������x��|<'����{�զH�ώ��B@�e���wN�	\�A���b�V�2	(�����q��?Y# �%)�i����:���5�ü��� �Ք���@���H�٧L�<��q~�o�?����P�m�8 ���mB��x�R��
��
��/y��h�x��q��'-�k"�i丱�s�<�ڂc�6�"i�,^R�g�T�>��jd�����a2q�\[I�A}t���>+!x����T㬔
��d8"�]�U� �=�|P�l�n��CXh��&=vj4H�C���!>�'#��2�M�L�C�\(��&7�������Q��;�wV�Z3 ���>)�8N\u�^�8w��ҁ����C���P�+�(��K92��"s���x'�S�M(�,�'%���d�g'��;Yv��q�-e�����0m|Rg��9���r2�(�@���>��Ѻ���Օ��?h���^cܕ�}�x���IN�/��p\��`�շ���K����p��^�3����|ƶG8�3˲H_21����҇�F+ ���]qb�I�XU�����u&c%S؊HN��B�����b���h�����C��y��Q��DZV� %�PQ+�a�AKS9Z�U�������v:�@�q�������'�����n����f'X1����#�M8'߃n�f�>��$B���썝jL|�)���ZJx!e�z�{�Z��Ⳃ�Al&�|컾�Ԅ`:���^�
����^��F�܃�ъ�JX�q����8t���O�p9�c'��~d�X�"��U�[���������4��H�º!%��/�w>�X9p��9����>_��t>[M����Ű�����Ɔ��Y�����>r ��z0���������'��? �<�d�{LX�A�:[���H�W*�U���5�0 �*�����Q��{�;��0�=���g �J
4�gޱ4�����jܐ|%��e*ZB�1�_c�<�����9�;�<i����Ze����.�iMkZӚvǶ� д�5�iMkZӚv5R 0�;� _���;H���	 3Y&�hh�0��ق�`�8,,(x�2�Y�r<K4,�gȮcg�e&�-��5\LY:�N}�ͦ����E=c>��2s9a��w�����]�}+Р��x|a�P�ACl���A2���� =�V�����5g�F;G���6T*g��dA-EO4����_�f(َ�t��BEr���(����HWP�F{�,�d�9�L�X� a�;�`�:��П�6��g���ڭ[��
\=�\�:���a�}�	/��gxbT�3K���5G@�ߛ�����σ�N(�[�ܤP30����O?/>�lnm�p4��+��+b�� $k0��5�	���]!�ߎ���nSV?�WWWa����=r����TYr�Q1��S% �y�`�H"�5��m+�"ɡ�2x�<ݵ�5�
�w�Q5��nG��1
���ؘH�����ž�%�#
�WC�ף�E���Rz+���*YϘQ^�a�M�\�_|�7��8_(�dd�SX��Ē	���]n(�AD�b0n�	���a!w����F	^�ҧ2����N[N�Y�:g�3�G�o��N��^�È��[,�v�F�e)��`�ڐ�y]c/L���;���iU�ɏXq����ֹ�>lmmE���� 
�
`F��Syg����B�������O�D�Fdk�KN`-b'�>�k!�E���g�^ �y�>����0o�U���w��!t�]���^k"AR6���������!�BY��/�	^�y~Z�X�D)�01@}��Z����g@ы������(a�kts�i��R�����	��18�[f�K������jW��42�:��F�?^��G�e�lT�%_Own\��D�P]@<-b�N���<v��b�Jp�_U2EbQI��t3�ʧ{žR��j�Y���@vU��W�F���_%B仝�o�����O<f��%<;'�a�A{h��&Ѓ'_~N�밆���<���A�77p��9^�x�p�2�Q1�Y�V�����F2��9m�g����.���xoe]���ר*�GI�U6�^����}�o�D#��T� X��+�k,]b}�/,�`t{.�A5�3UI &ۃ&��m�!�"��M�4�q
x1������;~>��ix�O�����:�úf�+�6�`�ѻ��P;��$b��Y��H�]��� �����*���Lu"��<߸|�'_R��9�|�^v��I���ϝN	��u	ןVف�����Ί��ԡ�V�'��nj������_�g�ΏP��t��sƛC��u�Ϣ]]�z��tU��[��`�Y!
�����׾�5��g�����.>̇]{v���τk�g>󣰰0Oj4H,��_�%�yk��Ǭ�m������w��}{i��D��[?�<��4�"�}��@ڟY�a��nD��ݞ�l|�z�x��7�ɇ���OT͏����i�����qM_>���_#R�K{���M�IH84�P�����y]0�[�=�-�Q��N�pĂ0���y��5�iMk��@Ӛִ�5�iMkڝ�|���`d=Պ�\#\�ঠ��5�e�5��N )~X�������.��L���er��3"[���1 I�~&`c�@��)@��d�h Y1W�N�	���c��J&��<u|,σ�QN2ň�1c�O�T���	�w��
�0�3f�޳% �3/)�V�x,��HOXKI�%]�)�0������r^�eth���
,q))���a:1CK�#�(�ʤL��j@Y���2ٳ���洵���3g�H�r%���0�/h�JWhi�X�z��,ׂ�L@@P��'0��a:��}���eAo���9C�Hv�cI���i	̼�t�(kw��U�
�f�|ˀ/�oER�Ux����ʯ����r���ц%����11�i�R�� ��+�΍��8��Kp��=���|���� K*�xN����l�LW�󥖀��%�ׇ�*~G��W��-\�|�\���m�w;1�Y��N�z���tL�4tH6�r-X����~�)ĦȪ��0��@Yk��k�8v��<j��EбQ���{���` �֎@h��`0������Yv_����p *�8R`qY�z/$$� b����{J����_\���x�)S�l�����,��~���h�w*Q���K@��u^�|е10���Z�b�h^^ň�d�.��R0����n��R����R������\/z4ɁV���VWS�]S#�N�"X)��D�J{�j�# �m/����bUuE|0�z�t�����䶽�*�x*�`�k�8E-�c�6D!$���9����Z�҆!� �F���3�~�\���k�Gd
1P��S��Y$��53��(R��e������4F���f��`�����dy3���*^ϖ��IH�P�؟�!�"� %���%kf���<jP	����]�/F��S�
�����H���s�w����^�!�'pIgg�k�����>�����D?i=�'
z2ȧ��-����Ke��VI�	<6����Ѳ"�,�{%>xv�z�B�p3v����M��D��aB�
��&P��lߒ�p�6�Z��~1���� f3I��!p�r^�t���9س�B1�t��1lOln�`m} ��u�=�}05-"��x�9j��=7���|���)��J����O�:^�`RCT}��#]��ڪ~-*\2\O$A��#��n��ڰ���"��H<���'�3�į�k"�A�s�����z��<��B���Vк:eE���DE�e�L��e8ٸ����`�����믂ۺ�� ��?o��Q(xz����b.7��X�~ʋ�#�ܼg���e��
1��4c��(ύ�M��A�́��5��@��?�Q� ��p���>ֲ�(����Ѽ�5س��;x��'�
�ο�ɏ��Ç�??��y�f�Ї5�����D4�V�F>���_�7ہ3g��aߎ��ă{����S�&����x����K^��g?�e� !{��p}���W��'���{�?�{?��Eh�/������?� �%���L�U����d���sx���>��w"�(�Nk?��B�#T�����y��:�Ι獋*9LA�� ��j�&�V�or�g�3��ۈ�����`����)Sˠ�k�sȳ���l�����Ԑ���a�Զ��E�Lݹ�5�iMk��@Ӛִ�5�iMk��<7�D�g+��1�hx�Ogf#��זIUS�W����.c��bȆ�)�ϧ 1�Z|
�����x��Qg���Db��{^��C��ě1�z}^3�|���@CJ����A�A��A R�P�������X�dA���d���hX�3�eZU�
|
��09�Ο�Q��)�q��@Q��*7�.23�����n���6~'�0����6e�[�ʓ�t����V��kIc�����y)�>����8Yb�.<ʥ�<~��*��5 ��2����7l�rrm�!hmT��!q��P�z�P�d,�`��3OTC]��hO:�����<���a��\kG��1�H풾�-جf�S	@ri|Q&3��������$��2�o�C�e<��q}�7��f�+\�hX�g��֛o��k��� �f"�HZP�� 1�L�`�K�.��4����6�z=��?���G�~�5 >_��a�C���(��~�}���=�4I�C�"�Ck�;9g�~�+���w�����˒�Eu�`#�"��eVv�����'�nY�lق@Tm ���N�Ŀ�����5�-I�qE��;��f��@;�̎~[���:�GR�ዘ��k�j��G����]��^�&�/8߮^�o�}�^�lĳg���sgi�a_�\�e�*�;<F:�L�*$����1t��~�P�v�������'?.�Ȳ��_D�j�l�ŗ�x�v�8��8�oe�%~p���7x�p��P�-9#��a^ 0�V��vz2����4W�'PJۍ��q��`b�FGe������u7]��z���� F&[�v��s�ݎ�u�"ߧ��h���e���@o5'b��B��b��=u� �qԓ�ex����3���t!M�.�����v���"��#!�=�z��œ��)4of�r��ݬ�~��>.�*%��y��CF����Z@�M���΍���Ɏ��T���B�\[ܐOG@�Hu&�-��%�O�zi?��W^��~p�ڞT0��r�p�6ǰ�p�߃��B��V�II���h;�c����X���Ԡǭw�=�Y�V}���pL��Ł�4G��8
-g�Fe΃�[q/�l:>7�I�F����g�ĭ����ɂ2�5�.�ѫL��{�`�ڷLh)�uTv�����,{A���J%tЯY�Ǯ��h*�����j�a��{����h�6\�q���Gx�����N�������K�zT�A���g��g�L}���+�O		g1�WUE;��|�}�/��|��QXÕ�WIA��
;
�3T��	I��~�?�ͧ�W^��'O���M"~�d++�B�:d2a�d��x��yM����:n޸!*K\.mieeE��=������A�c�S�p��9s��P	�z�H��~�v�:����G$�Lw��>�s� ܼz��0�R���^����Nh03NEo����7xo(k��C�����.�Q�	϶b�����y����G�H�ҙO.<�<��|���$�O�fk���|����M$-%�-7惟K�s�i�<O0�9�dk�ִ�5�iwpk MkZӚִ�5�iwV��ZJ4��Z��1 � �$2hޫ��P�G��gQ����б�4�GLL0ci�T�[�v�����hM0����eiZo\Tŏ�1L&�#�OAd��@��9\br�Bs��.H��G���vҗ9�U�nG ?�;�~E�W�0���c�K	�irML	����dW�&�8�O��8C|U5��S�&8���)_�{��f�QB ���B�
��P �Q���^2�LBp�{,+.��������5��-�- ��2�j���姣�%�9;�V��`�d�cf�W+�i�e��3�������RvfF�#�	lk���68��HXW,�O�f<���2����FY�4�T �}��k�^��%���de�T���>D��s�̡�*'�5�F5�R=�[kk���YhY(����n���SX�@@*�C%�}`�G�KX��&�#��lmnXƊ�%e�,��� QƘ�����x2���n����L)��K�`$�h�; ����ujr6��3/�. �@hX��e�	�:�P�q����&�Ma>��>x�%�6��8��wɆm��k�v/�����}r�~ey���|�>Dsk4�]a9�cB%e��޼O=�4����<��:����2f��Z�D�A֐���oLʪ���t~&��L*�k�ՖMpc��0r7���<����1��f?)�3y�(X�d�p���(���B���Jp\.�ʚ���e����9C��܉�z5���в0�	� ?���&@��S��� 7:��~G?��}��i/�����د�9��&����0C��`���Ι�:�����BL�� ���ϵ��u��뷎��B��g��.t]���F<�(<(�T��H�fU�y�kg�j�2��<N��RO$wx]�峚M���0�Gg�]`��l#���=�]�i,'%�>��1�t�F}��|FIs�D��(��q�p9�)[��C�a��fnLl:�\���d:�.t1�k���a�-��·;tʹ&�Ĉ|&�<5�)�=�Ͷ��]�Ik`I	�i!�3��]C1S݆�z�)�� ��I���	YL���ׇ�%س�="�HFhɸx)u�PI�PxO�1�wj��
"�z,�9ݖ�.�)^{	���y�I�֫ZJU`O�%��p�i8��T�)�Pc��N[�1��k�i�ĕ��ח�����ک�>�g�=J���+��٠D�(���}x�k*�FDTj�}��yV&���5�H�eZ�¿i����~��U�l��c��=�%�E��U���m^��� �ܸw/oo��ϽH�7�1eihNki)k?KJv�Ox�@�����0��ImJ�|��O���4�Ml�7n܄"\�Cp�J���Bҍ�!@u��g�9��A[��� ����kD��(�E*�J� ��1YD{�������Rh�I��`>EF��y���f�1��d䤙�:�~z��~?.u;d����$��r�6#
P�:d��X�L��Ϭ�6��I�F$3��	c�li��ߕ�;�fӚִ�5�n�iMkZӚִ�5�k���9����\w��*�,M?�}��C�Պ�@�WK�b�X.�P�NG�Y0%�� �<�������.�(8'��RW:�e�� ��"9E�l74P��;�Q�5r�4��S�J+���}j��"��A���"�^:�"g$t�|���nK�P+@K�X2�J���" p��HqB"@��%k:�)xo����z��U��3*Y_z�R�����4P ���A��/0���+���[�`+J�pUZX�������g%`��c���) +�D�l�.e�{���ϖ���*	�%�W���D 7��UF��A]~j�٢D�
�jv��@b���{��d��	Az
��V�Hu��׏�c��E?)x����d
ۃmhk�6����ϩ2��(�!o:Y��{8�v��I m�y��s07߇i�a8�>BpX��&OǔY���H���5+�����$D*���P��3��N�������t�RN�f�����D�d2:G!d�į%Zol*��v�A�؏:�L�BIk��/�C>����l`��̜���e���ئ�R�@ T%��3BZ�Y$�p��ر��3)��������\�v�:s&���k�w:]���Dʰ�������0OH�a}mr�g��G�c�,x�'�L�sL2��}?$U_j ��W����x��@3�p���ۗ�
V21��w�|Б1q~(���A Z·Ǆ�Z[��W'ա6R�(d��b���k���Ӽ��lEĢ��m&��|��୉�����|����d�v�Lf� 苤��&�L>3o���L����{�\� ���0{�y���ӜVP�"�g3W�~O���kN�<�*��>7��ݠj��E"hG���C����H3�N�7�%��}�wG2(Ȟ��Q����G����9w*��1>�OʾC_��6�Iή�*g�0
�ҟl�@5܄� ��jKa���NL�?iw�7n�R����ϒO�f\C�u`���pj��Z�2�����4`%"���N��9�+4�5���(�T��1�A��,m9�PT��w�"Ɍ��	\�(i�R�x�x�:�cd���!�gX�I�)ᵖ'��$J�}δĦ��L��x,?�Q�M�s
��OYV��[myOR�,��$����ªִ�N[�w�:�%^h,�3�v���d�m��{��oD.Ž���H�Huy/�0��e�z\QDJL��tOZ;�d��E0܄�~����c� �>}��O�=x�O�����֭[��l��z���ދ�"�Gy���V�S����:&C#���J�5���q��}qg�Mk#�`�,��;��4���I1��j��?Dr�x���}ܧ�h�\	�}���B��!����otF
S��s��M"8��2��f�ԡ�iy�T��af>è���a���ꨔI]�
(�/�N��,@���Jk,R��u���R�/�z�;�=Nv�J����r�<ֆx��Դ�5�iM��[C hZӚִ�5�iM�Ú��N��e�C~�f�ڈ+����DA��z���쇢��.ʠ����\c��&p�R��Š~�V�k�@5GB((A��NKx���Z��UNQR���9��`����)��G��o	j�s��O)���CF2}M&4:�5���A,c<���n�b@Ϧ�ӈ��ƻ��I)�M۴`a~�����(���cP<fΛ��gҾ\s<e#����]��J�� R*��]�����2�U+Y��:)�>��9� -�M�}GpVjԗ1���v`l��[e���>���s0�j��*�>u=v���I��4��'VҐ�ٖb�l.#x�$[�G���[ڵ.�W���K�k��
�R�3����/̊'y[��	��ٷ�w<�}?���\��TOTUH�s�~����4�ݹ�����Z���E���t=؏<n&�!��O�4t{r���J6f)R�a�
IU��t�Q���1\K����(��+�U�K�s?�spꮓ(��<��Tﶆ_~��������'�ƣ����Ʒ�w�}<�c�j�<q� �~�o�?��o�$w�`#�! ���sƬz]�e�T6���T���,wOY�-KJ ��<��e� ��v�5L�)l��lW��0�J2"���s�-��G5�������S��wi&�S-��_��O5f�Q��?Kj2
���g�Ƿ����L@@;�"M��J-D����O=_���IR�l�b�d"!9&�`�O&_}������b�O!}�9��]���Iˁ��㵱� ����E�lE5F�s��F}�._K�8���>�L$��Z��;(�a����q-5��!1��&���̿𕶕 -�Y��\ ɇ��K�7��;�;MJBN$����^�7�qp[�П�-���	�<Csm��_/���d�Iʺkt(y��V��q�U뎀K�e���y709��}Td�+g��� �U�$�TU�iW� ���j-h����I�ű�����Ե��L��n���۪���H��9��1���H�}�R�*�Q�о�5�����>�"h嘼��轀k�/U2�͈$�oZ f�E����a@�@AB�^�J�Dpk���P#���.8����k��'���P�`I�g��M��ߡ��&́Џ���	~���y�q��W���%ZO�ЯH��}��D#U�{������'�2��Jz�
β�����q���񉃭�&�yXZZ�b�j�vI��m#$�kf1�k��1�n¿��?.R�L��yn�����=:F��Z�ڶ��ȰO�&5���S�snSٙra�j�d#Q����������C5
�㸂�d�3�Q�~?��\��D����W��Ɖ�p�}��nId#kHUz(k�����}m���_&B�Uu��kZ�~[̌�s.s�r_qy�b���Sj[H^39M���kT7��P��R�b�Z�c��|≿���a/2�/#8r�>rHr-Y���+_�*|���0a,ØMX��@�$X+�m��>#�#�=I��X�f
�����>þ�Lu�a����ݼ�����.�[����s���7߄��~�-u:X^���G����'N�qg��׷�0����k�����ݮ�vt�[\R��G�g��"��J�CZ"��t@�WT�-{��ArĨ¤%��+r�Z�!UGUM�UE�]�.E⮬t�5�s�iy��D�n�>�D�H�ً�׫��K�s-[`�?��}(kZӚִ��ѭ! 4�iMkZӚִ��Ae�:�GX$�\%/	(Sp�����@�@&㫀;J�[�.���}{v׋��յk׫�vns��E�jM�U��/�)�˨U�]U&����RV�5�i��
:�����^��)ę�?^�I|% pA�A�acɽ�~x
��^�q�xL��X�(~�� ��*AB��4��eġ@��7��� ;f�b0�����	��)��� K%Ǘ �8%�N�ʳ�M��gYu�0|fO90��\�tʙ��$ Ș�$ 1���#YU8T/�A;����-�tN
��Z�_���G��Ç���{�כ#P�ʤs�J���Y�	�ex
ʫ�F��=��`P�z-S������\?V�S�<I�$�^S����\*f`u:��vl����hQ���u�t���e,��AY�c��7�6I��}�g߾�g�#�x�<������������g�����}�����FP��Y�3��P �A���T��F +��ʲ&�۱��*�PGA��X�y��}�gE6DU���:m���`��ɧ���{>���᭳����S��������Mx��%�}�� �d<�6�.E�,�^ӵ��J����#mۮ�����x������?�����ܾ}[:�%��Z&�)�y�:��f�O�L0O�}Ty@�|o��
���\�r�l�KP ]�Qu���[,��%2 �g��5��@����H�W�6ı��㟀����������-���p4&R���&Q<x�o�s�?G����M�aE ^�T�}E-$���V�	���!T.�t�H���W��f�c=�hPH9͌7�����s��Zޗ��(��{��d��}��4���%�)aL��^�Ov�D$�Ԣ��䤳��sq���r�`�V��p��������yK%A���oB�%D��&���I��(����"�Sq��|��װ���-
~G�+�%_"�x_�3�s�~"L���D�@�
��
��֝Ns%s�>73��:薍�=�
���9e�?Te�d�;�Yk�3F�+�@|}8BKH`iRA��Nܢ�o�W2h�ka2IO���G%_7f�R�6��g�����rrb�l��fi���O:��/z��z��pBB�����H/a�5����G0������(���G�J�w}�[�5�;\'��w`���ֿ�",�9[�����D�g�#*��A0W���{��$.P�.�	�f���@���_~���z3{��>�w�8�?��v���p�7�8C�f�7n�����}EXw�^�&�E�:�Wn|�1�r5�$-��օ+���OC���&��WD��)�ۇ�ŵF�����>��p-�;�$o��,Ͽ[���b��V7��]�C
/&��מ��'O��<ۛa�W�,+{K&��^G���'k��iI�'������ͅ��ie�Y�{�z�kۤ,@�9!��u�DH A]���d�8��Q��%%{hN�L��/��/�/�W�%���_g����Eċ^X7?�����>E{6T�����4A�#�a���}�#r��%���s��_��f���5:��`��}��#	����{Fb(��<�!R �Z΄T'���D=\Sq��Tr 
"�۬D#{cй�k�1�������ci�:z����r�Lfd,�s��sX�cG�Bv����v���0�]�wzn�W�tA�~���u��0]�e]yvG�]$DxY�>�7�`X�O���U�K��<`�-ZӰV7% �ִ�5��g�! 4�iMkZӚִ��a������N2z�E)O
�Iv+�J)H��(�hc� k<����n���u��?��K�{�^����?�����/}�K��N���X�Vu��5���4 D�1�5��k�R<D3,b 8%���g����L���jmD�����Zw9c%++~_��x��z�/��X�9CФ�{��Ѐ!�Ey6��;V� YDK�>������To\�1�#�V���k�ܧ�uR#6Q�`��Qv�e �b=>�!p�K0�]l�o;��A��P?[V Yb�O�ǎE�yn~N�<�=r:�9���`ii�	��L&̞Ǹ�5�G5��XK�U�2��NY��ʒ3�)�7�%#AC�lžܵ���� 'e�W|L/�LE�&�v<�����A���[��^1�����/�H��� [�G�����*h�c�Z�{mmν}���O��{�{?<��sp��ux��G�+<��? ��}z��w�2lnmq=b��N�;�.gr:���'��a20"��uG����$�^�A�L��@x�����l�R��/_�7�|�W�(9qr��x{mH���6no�F���������>ܸ��{	����7oݤ�]�^גuΙ����RJ����.p��y]C�����'.�}��u���h�`>�K	t_�pv��@𹰶���p,Ǔ
��t8��c��?�4fe���xM�� 0�D�c�?#��T^�%���%��*/3T�#�2ɌĬ�V��P�a^����{��%� I;TFF�p�g�0��� �����0�=w����_؀�|7,������0.�p����뚰2�s%h��U��Yw�OD��t0۱Ա���}�.w��9]�fd�3��t�R# �!�� �GV���N�_P�}�$� t�f�
H�9�D�>�?��(+!BUQ�Z� `��*P�	�@s!� ��׺F�4'�4U$�ùdg����5Ľ������mL��H�����"���3��	��y�t�)�����N [%�3dOXD�A�kx&#�y%D�Z���e������f���	��;-�w	y�J9�ߐO�2&��܏���v��^v�^��p8��W�x�d���-W��[7o�軘��I���i��%��4+*	��DR��tl�gϚ8d<gm�{ZCꈖQ	�
Q(w������<���	sK�<wH�G��{G��a�m�C���C�3�`�u�=T)Bߋ�r�s��kĵ���a�/�kj�⯝cB��qC}��/�^���/�{������p�nw�&�p����L�y�:)
,//�����"�µ�a;����
�6��7������`쯷{<�⸗G�ۻ��"��{�H+'�Ҟkk}@j~a�8���E�!�஭Fe���?�����KVr�u�݆}�ϿLY��>�>��9"�M��  o\�a��c�7$��,�$)����><�a�� �s�}��/�G�)�����<ԨXlg��#��������/o��F-s̳���ݸ���ie?M�%Sí��ǿ�����������ѧ��>p���xʾ�Up��Q����Xد=�?�<|�_���<3�z@{
��1p�iO��b�к�kb��3,�z{�v�k��^��7��	�1\��Ɲ(��^c��g�n�Ժ�|4E��	����_p�ԤX�j���JH��S���=�� G �%��r/^�(��6���V�܄f����"�_ч.���魖A"��~�ϻ@6�|~�J�5��%��K��ⲬM딮3�>T?gҽ��+����hqa~V�de޹�5�iMkZ���� �ִ�5�iMkZ���j�f�[,��!	Nc���<�#I�4���aʲ�sӿ��:~�����ŗ��/޼�{����C��?���<��3O���7����+K�(;U5m��9W��!],⸘���[�Yj�1y=����>���]��N�?�X� ؜��cf��}
�0���$�,j��J��Ѐ���H�>e�^	b�W4c�n)˂�����d��G�g�� b6J�D���hP0b�)�ڲD���n竳� 0_Jr�z2	)�9jSF!_��F��㦵8��yW�W�.i����7Ơ4��]��P��Iz˶�²�;֪%8�s�T,c� �`�,�:%��tx��W���p��Az}iy�noR�<eK�c�y4���%�������G��V�%�YU��pB
긱s���%Bb6[�jXT���[kx���k���Σ�m�ݡ���p��=�������&?rnܼI�(��%P*N�(������!��K�πʢ:!H �9��E�Cr>ѧS�._�3g�A�"+5�ۿ���u$#ړb ���3�*ʂ�t�2��-��-Z�d4����Pyk�
^z��1�����>�bTn�,�mI�Ǯv-8w�|�{��w���޿��x��G`��6lna���������z�����
c���Xv�Y��E!�DkP�j�+�!b���9k_���Ĺ�D�XWJ�hpZ�9�c#�e��{�X] 9!�(̶Uňd3��P�J\�� ����>8~�.XZZ����� y���p���A�)��sg�_�3� *�A��=M~�W$�΁ ���f��먨���J�"�IL�{=�O~��
+*71䟂�.�S���,۝�L�f�*��B�fT#�?��\�Ɛ����̾��Ҫc�0 � }� _H,�H��D&���P�ApX�gU����K1�]F?� ��l/'�}ɮC�eڡ;@%�K�G��k�����w�7�,���<Q�X s����=�0�H�3��ɴ3�1�]ck�Hr�ZԱ�e�����C���P��H�"�~hKT�a2L!���zv>��	{��v�$� �0ƒ<H�+PrM������/������0��	��NU6��D�T��Аu��Y�t���#u�T��jV��� �@'�]HP�c�?�gv��o���]w�v�􉂔��paݰ8�z�	�5)�POK�	�����7K�Wc9٣�I<E󞙸�v��>.MT̼����y��8�nø�"��6\��[S�:ha�*�/�p�i����U��߳�0|���ο}�:sRs�v@��=�����0L�x�������:˻�С���qi�n��'��O���ґ���SSy$O��=z���C5?nZ�UU-��I��S�a�9����î�'`s}���jmwR����?~���=��ϚA\�
IS��G_��wp՝��c'O­����^���E��wq�p�O������#+������ֽ�>�ڨ	si�4���<�� ��`:����[�����?�"�g+*U�Q�0W��P�#G���p��?pN�����&L�q_ͥ�xM"��4ᢟ�L 4E�Dޣ�\�͵�^�1��+L�t��� ._�BwW;.�}2�H�
�~$-����p��i��k~a>�[@$_�)��)����҉�#��U.�?��J���lc���6��X:Dʋ�G罈5Z�M�C�܆U�q}�u_�}�]�#b�����+�[I!����T��'���1�jy��Q#Lk��$��Ӄ��ٴ�5�iM�#[C hZӚִ�5�iM�s�w��ƘQx��7�p4��R��1Y�C�� �{1�(\�]V=�����﹅��j/�֞��4֎K�:��s���W��{�w�G>򱕳o�q�?���^{���eY�B���1o������~	�Ѝ�� �]kZ�@:7�L�:N���p2+� �,��d�'H ��k$x��p��V '��h0b���a@F)����@��}H�S�D�$�7%�V3XR�d��x]
Qe��wd?��x&H0xhU�W��y���~����n���Ͼk���
q�-�u��L�/I&��^����+��J��E��~��[R�����u$�o8X���W�^������}.�zۧ�_Z?���c�O�&;Cpd���={�^��{V����d�Kˋ$�]S��"esO�:w�sV�V
/2���l<���P	�8ц� Pv�	������c��٪BR�z��e��B�ۅ񰦾E`hqq��#�^ǣ	ՙG�P��R>vK��|��J��$��@_V��	�O�*% �j�R� x�����E�2�;���p�*��t�F������z��PJ�}P��#@��͛����u�M`F+�۴�~����o�G��`@J���:�u�8������11��������s/�>��Ѓμ	�.]��poO=�"�/�������^�V���_}>��C�[�� �5)MHf�a���i�j݋͘��$��#��Qi��$��ߠ9��?�;q,f���*X(X�#*̀���A�B�<'r���8���.�w� gP݀��P3�q����׿FeFal+�\L�!���9L�9(�u>s�I��~x�縬E$���$P� ��|5��� �!ҿ�G�7��"�ݻ5�W탿F���b����D3������d�
t�5�LKH�|"�g-��s4U��L"�)8�K'�AZ���$;�
�\V�,��?&���(.�e��Qɏ&� 4sT��3�w~6_�D?)|�G.c�ߣm�ԯz^��0
z��t^F`2��V��N�����]IL��ב,�j8&�Ń����?�)X^Z�/H.��������z�ln`<��?�I����ac}����TH��._?�#��\c�N��~�'�>�����4�q��H�#�8��r1����~N�5HY���3�2ؐ������6/x	������Z ���m�׹�0'J^�����k�CՊ������"��N�Kk���[��d)p����9d��=�;k��ϱEG.\���y�څ�wh#�U!
꾒�M�D �5a�qxs^D���2��`}kڽ9B�i]V�(I	 |��Ck%���5�VX_����G5!2R*A2���U��p��(.Ta<ڻ�V�0�T��c�d �-�ݭmls��k/@��#h�R���q���������Ľ0��G�X:r V�o=��:��� G�Lw�H#:���I��������9�/��NT9J�Zl���Hdϰ��R�.^�˗.��&���p?;	{���'���>�}�#�z_ñc���W_�>�lV ����}�\�q���W��e�_b���*�3��Q�µ������W^#%T5��tSH*���Ymdia	���x�Y+Y��u)����Yq�0P� ��rl�{!ܰ�E�(z&�&O�ǎ�4&>�3��@�+����QYyyM��,���-�$+%!{!��D*J���&O��!'s+�N�]�u��rD�`͆V8K]����z�!��:MkZӚִ;�5��5�iMkZӚִ;��Z���m��A�ۙ����$��*�18[O��,[��b���s0J �n�o������iu��t��nw�>q�[{��3h����g�v����޻N�>���d2��/��������\�7`ZuUQX����I*���B3K]*I���U��3��}��# dP�L/�mFA�i)��4��t�8S3c���iFkDHֳ��M�>_D)�l�%��j�2���9*���v�Ar/�D`�|��Eٞ��[cV�d,��H9ҔU��!�N_ ��[�*Z��S��orya30�l6!RM��Ԡ}�'��6�e���f�k@$�χ�Z�ȳT��C��ϟ�sg��`�A��C
z�w��Iř���_�ʄ��,��Ĭ�&K�%��<i�O�Yw̫�a�sbW��ľ�x�"<����O}��>��{O��� h&[�0���я=F}�*�|��]Ƕ��P.8���]�	hz	>{�$E�E-@�(���v�]=�l��z�[�鈽N	_�����t��_� �3Ά�d#1��B�"9��# ,����
�fW:�5@�r2���������2Ҙu�3�&�6��������Y������s0n�j���E薘��~��V�.��4�/����Ix�\�,@<y!�c�e���π�� �9��be~c�:+0����
lnmÉ'�s����&��,�=�i��9�#'ׯAo��Y�{Ͻ4�e��iC0u��px�;���tf��΁f�4�H�I�n�����.��X!%��%���ԇ�ۖ�v��eiDm��f!��� 4���t�E�	hC�����%&��ے~�I"�
�w{]�|�,a4܆㇏Q�,尵=�:�0��P�����R���H�f2�`'����à�O��^�>�Z�.T������Ч����-���af5�L����3�2�e:�H�Y�+K����1�K@ ��@�c��Q��\�(X�i�>u~+X���q#��#~o⽥��/bS*� k��d�|�,�qM�4��IoY��욕�dtoa"!0~?^�� �@���' ʊ�g �,c-^#�7���u"�	r��\��G)�됖��H�Q���-�����;-QaD�3�[��18y�T��F�[4�(�j"�O��.܀^	.^�@���v	O~���_����?�C��9!��D���F���,�P&�8���3�+���z8�];��!%Du��O�Q�øY�؎�(�	U�lo��3}̳�1Lߐ^������¦�²�o��޽�g�/E���\��OY3��v�X��}\Ӂɉ蓪����Y�=�.̔��D���8D~�B��u�7�(G����P����-�e�G� ���Aw���6,�Z���I�;�w>��=�C��R8�6Lp/�c+��7/�Á}{�y�x�0��`�-�[��w�H�p3��M��[�OI_��T��Xp�j�e��Z��(�O�2s"b�}��]�}.�<�ҋ�j-�����OP\%�aP�~�aؾ��z��xN���F�UI|�mA�<H��=+Ȟ�~�7���ZM���L{$����^��qDU�R&��?�pج���`>����z=x�C��붴�*�e,�A�.�\%i��F���++�]��Pu�]��O�qn�o��I}�H�c��!õ6���	퍧De{�q5h�S�����óĔ	���oV��ym�<�y.�a����k]s��lS:f���ڢ�/%�!b7�D��R��$���,����^3�?�Up_�N)��{ ,��$�$|f��"����^��g�vI�J��s��w`d�F�aI���p���y+\ܴF��~�Fek~^�s���Qk�MkZӚ���� �ִ�5�iMkZ���˲�L*�1�8w��Tk�Ӫ��ZSԕ���UN¿�-�Q�����I�hM�s}��u����_ٵR�{���������}���]YZz�Y{��Up�������[k��p�n���O��O��/���7����kkG�5�`l	)�C��ؚW(S�,�(�����6��$ ��U����e(����J�&B�13�^�O��ƚ"8�C��1�+�1|F��|TC
��ĀU�2%9:/�1,W�YD*yi%3���Z�@�����F���G��bP3���[A>���R�+�Igؼ�E %g�+�����J>�ɂ�F�:ޓ����݂�Lx��P>�M�lK�B�B ($�8�T'b ������'�L��ؚ��+����zb�k��-�1dp��]{�$V���)ץ1�[+�R��Ȉ{	:����V��T	�����o��w��Xuzsh��)xw��1�V� ��{�]�ާL��H��� �ādW�L������Ї�<t�����}��t���`.f�Z��ξ��a�0���.���D��%��NH&�
_�O���8�u�@$�#5�_�DKY�A�Ձ�qo�������p��~8th������x/��C����=��O�j���?��x��I���%Fj1����D��9��J���@�z�\f׉M0 R }���$qkʂA%�����ph�~��V����݆���{���0����.x�̹0F�f�u0�8˟|�"E��Z�EA0��r�S"�#�_;}6b��dn��X���?P֘�o�7�'A�s�H�E���5a�z.�@W_��>ͧj��z�. �@�(���ػ�]tZ"��>u��?�3T~�	 �P	eǒm��[���N�$�g�{��.�r�*)s`y�7���N�򘶀RN3�w�/�m� R��S�v�S��9��?I	������l��3�ߤ*�i��zѕ�D����
��-�j(F�;+ ��3�?[�W][��jQqQ j%^�cf�������̊7��̇@��'� 08r�w�-f��MԬg�	;��쵦/ �-<�s7��o��KlӚ�j���bW�O�y� ��X=mP/��K����@P2�z���/�s��u�'~�'��x�7�m���O����'5|�N�É��>�W.߀��O��K����2gΝ��V�#}�\���}�M�,�tL;�Q+{�31�P��J�)��I���6����P���ߙ�������������m�Ug�q=#�������r8B�!z��k��e��\��.�����|�WU����0�6�U�!]ǀ���@�W!�z+DY"�B��'�WR�! ��--�]/��r.��2�J=����_^��4{�-4.�/t}GP�r�%K�2��! ^e%>�fSa��$�2�"��=��3'���&�s���Q�*��SN��7��;,$N�p2��66as4
�����_\�+z�v���D�;w9)J	vLTRNi�t��q؃y�SZ��'R����p�mx������σ��DR&�r69ӆ��M��?����Yp���8/���MW�^��L�s!��B��g�I�HZ�d�c�tCd\.f����l�k��2xhi1�kDw��'<�3�|q�����G���E�X=}ʋaD5��?��{��qֲh�L��v���u� ��)��=
����5i�FWɥUp�b�vq�*I��I�ɪ�
@�e��E�#
�	��������]�'��`0
�
����w�����,�������(�ִ���l�iMkZӚִ�5�h������v{�я~��|����¾�laݿ��+eQ����5lwڃҖ�eYnE�1��V�(����3	�������g.;�,/.������T^���v��KW�^}au��՟�ٟ���3۷�omw;��ۣ�9Jբ'��Um������ue�,Nk�ҳx�N��M$59��I@#�Y��moo�'�]�ʠ���A�ɴ��Q�������5t����l��p�e�7�jU�X���r�(�H��Hz� �"��0վ%0	B%8�3�����D�����~f��{� C��$�!9���1{aKӘ��>e�	p:�N�����`2��.f�!0֑`9J��Zڗp�L^�{K�˒�`%l8M�z["��+�,�����!�ܦ��Ĺ�N��ul�_聹���<�N�r'�ﻎ�J�s/�Y�<�7�e�9�u"�kf�ڋ,DQZ~u�n���p���� wl�Ɠ
��.��,�<.߁M���؞�|���߱���L+�4M�;�R�غ��3��7�0���矇��9"��ݺ���BV�� E%͹��=��k�x��y��H@��{��0/��^40If&�S`=U%�`b��O�7�*0��s޹��E�$�����_�Sw�����#{�l��y��s��._�O=�,�s�{����p��9x��(coyi� ��߾ �7������.%��?�T���%1��)�S �X������.��#�@�¸��=�pk���	�^}�A�u�&\�~`4� ��^w��������ܤ���0�rX�I�%e���I�`��1X
�	��8p� 7�S=n��B�p#�E�����7qn{'�V �4ԥ̿��:t�%�;^�����V��9�#&��Oli\j"� �o*�.$'�|��9�ZX���B��޻���A����J/�5������s�ׯ�w��� 7su���Z��ůj���0ޜ��+P��� 8�$e!�h����LV�r��%'u�);��%��g�~��}�����L�:+w��#|,��ߩ&e�V�G.��*��e�+? ���u�R�U�|�%�!��%�����wPQ�n��r���҅I$�g4*�&�E%�l��C$���g���(��/�j᧳h�?&o��v�wZGp]V ـ����7,,..@؇���?����ߘkw^}�e8z�8����^�U��RB�Ӈ�ۛ$�����G��dc�6t[=lq	��{�J�|�s����ux��F�m=�H��ο	�?����F����-�A�c$���T����p�ͤ|`\��*�� !�s�eL��o�Y� RpR=��-㒬G�B�DF�i�U�P�2ש�b��!��fC{D���e��d+HvCbF如X2�
��+�tK����A5�B���`��5i_�R��;��M���<�S9^���e^���o�y��N8�X���5�r�_��2�J�#�U�>$Ca����&���FE\�M6_e�q/&ceX����	��g��|�VJҵ�&bl���=��Lz���{T۱�ρֵ�R6@�f��� ��E�,,�#dP������=!!�Ek��������u��S�r	�T�ނG��Gx�ɘ��[7o��V��[-]��W�H�Rs �7 D[&
`CRpq����?>�5Ƒ�{�n|����>Gӡ���y�V�~M�)
|HA%,+���nP����d�{Y3M_��bKl��}����o2uN�4�kBs�����y��Q��U��������PP�����b8'�KR7b{$r��Q���U,$%���Z�L��Ɨ�}��D�sH���J%��$��p�������^�Sػg�\���i5>e����tj[�m^�ti�}�w�ޏF&w�Y�]�-��,�~��_Ѿ-���C��>��}����ϳ�������}�UX���5�Iy��އ�������!4�iM�vZC hZӚִ�5�iM��Z�߿��~��x|+��b��`����ކ�_9g'ֺ��6<��*��˲�gV��A(˺te�J7F��t:,.."Q�������7�u������<���y��p��3�rm�W������������7�^"���k�������'����O?��H&�U�����3���m�[O�u�*�um����	�礚�1�#��Tө	߷�����}�T�ϙ�\o1����*<omkW�&�qP��hB���|��p��tR��q{<�77��7֗\�V�V9���ä́�j�q�>�M#�L <�!�`;ɔ�����h$P���,q����w��-Y�(q)�:֡�*7����$K�AG��]&LQ���8�E5�)�K��]�b�I���/R�w�?O����k���P���IƱ���|l�&�g���B(��.�H���,�m�t���2�����]�SQ	��\��ˋr_
�Q��E� ��A���A�Zn(�M���;�S�|��ν����������0��W)��4��;�^87g�^�r^|�%
,��ط/��$�Y:�ơ־�شjB5 ^�����6�>౩���M|
b�������o��$�V�J�"`�m�0�.�|p�F��Gcx�ŗ����B21���	k7��6��[�4�^�\�&�Q���hE� ?� I�3��o~�IX[_#�ؿ�կ�G�	��*<p�SOv�Ag�N��?̰àt�ׇ3o��TR������ܿ5L��V�,Σ�<N$�|��|u�Ƹ�	9F[���Sµ  `���aBu�!�I ���µ vK&Мz�g��ǿ���I��x
W�����H6��@�Y��$��e:�B�e�r!RZ�Jf^��AL���n���G��ϫ)ϙ�^J���Kͻ��JP�B{+��}5��$��
j�ీ�	4�yP��>)#L�쳱/��11�0��w����E���`Cj,�TC`� a�H�{�ύi�٬H�@��]$M�(=�ef� ��9�;vE"���C��dr(���{��%�o�z�;��@r"�)��!�vփ�M�E�L:~>�CF��P��V�NY�T��SÁ|�����^(;-h_��	��裏�ѣ��O ��f����������߁�}�+JD�kYZ�M��v�z�����w���ǎ�s�us4���M��>t� ln��ŋ`qnZ���u�	8v� \�tΞy�ú�����7����>�a�~������<��6�%ͼ�����g�<�9fI!ڷqlD%�2ni�p�s0	��R�MdJ��KIUR��H�d�-��&ֳ2���%�ɮ��p=xR����Y�F��}��&�jr)!�k?��@�)]��G�P9S�����(���B���ltq��fF�Q�}&M���i�n�u���~�3���^	pA�R�Ĩ\��Ȓ��U���%�@���RN*�����C�N�D.EC�d�l%�,��L�&%�H�$ �����{w�׳���� �S"�v���w�C��ս��gq��qڣL\�(�@-k�dK��� �8\C\�B�q�4H���b�8H~�1���G�
>yU���UZJ,|�,f<��o��٥a��#�,�[s��3=� Y��:&U�鼷t�Ʋ}�ko�z�O	�� y�J#���S�Y�5�ۡ�Р�)���χ�2J����S	{'�0���ٳ�pZw�_�>�O��/��q�RK��e�l}/d��}�vVz��ꝑw���@|2V��$Z�R���݃��l�����ᑆO���M����-��tI~O��8��8Sҵ!�b���+�$1"��LFِ�d1o���cQv��c��v2O:�\H,:7��p2xnk��\'�KW�y��:�����Phb�s=������ @K#�ǅ�,�����b*hi��]\����������Eʥ��^���g!4Vi�ȳ�~�U�>K�~��p����엾�Տ=p��A��'�>�(�jն�I���mZ~:�p+�������QL�o��J�F*��y�V�.�U�*s�ѫ�J��ף�I���!�\ k�ٿ��k���>�c�m�m@Q�$fO��-��u�V�#z��(MUG%k���6&��g1p1�K'���HC�������S������-$���,3���/�i�tªj��7�o�ӰLc>�Z$�[�y����a�&��B�z"@��ַ�`�	 }�[��ַ���oE�>��C�k�'�3��c�s�_]�F����fou?�~_�����k׮�k.0M �Qx�����ӓt-���wk���:7�畗7�G�Wޯ�u����w����wB�y׶U+H���5�ߧ��J~o]�=�����������Z����^v�����n6�KM������������|�i�!���0-�5p*�P ���l��
��4�eW��i��;oP�����!�X�V���䵆)N�;!��%
xv,�4������YD�.�	���N3�c��H��MOg4=��s8��-�U��O��H�{hz��d��*��C�m��ڂ���`�W��#-WK ʜ9� �g��e��?���5�5�La%�MBh��ޒ� �|6���=N����?��^�(��lD ��4>�5ٓ	��Λ�����3�79O��5���x��?�s|E�����>��O�#�>L�}�;T[��#i���O� ���@�.�c1v��G�B���2K���N���s��M�2�3��Q������}�0�͜��y-�؈>��'�H�;w��iio'��f'G�n��R��4���4댢�`�\��~2���eoY�'g�?��#t��Z.L�����\� ށd��^庹�la/�X�2��;{!�ۚvGB�3<��"�AJG��H�5uNE��h���T���|����B�^��g�}�>��'a�w�ܡ��@5 ������(���O�Y��.������%=8��m�N1��6.ۀ{l����n\�)�F�r��=�Q@0�i6�;zO���,ݹwH/�I��fӪ
��_��L�Q?���I�����|x�۲tp( |�`�6�� H 0ᯟ�=r�r�V�����̓O$��5�B)�>Ǖ�I��Lfk
��TW��Yܳ�R�,;^�(��,R	��}�3hNJ�*+�����1��r�h�Xwk`����ɨ|��T :9E�7[���@�������-b)��	�B@v�dx���Isg�D�+.ї��%Z/Wtpp��ƿ�7��k2٭�����ݽK���1�@���~��2W�
u ����ۡ���۷o�c�=�|�d�F�1��N�0�{���tzB~�!���>��f:Ͻ{B>x���y�{t�Ξݣ�Û��[�o��+���ob.q�p�(�[?����d�l�d�Z�7l�:�k��jP^[��F}x"RRV[�^��K��ÂW���=	@##�p�7���W�1����"����?����xY�p�,ُR0>�����;��0��V��S���AF&/E�oU�'���PV�OX�_�)�������5�b��,s(MD:q�j#٦�\rx��� �k����@M+!�C�߮�T��`Div�ցHY�d����?Iv��Mk��zr�
���im_�Y��'��4Ę��&�tqȥ��~9�ͨS�5�D�Gw��� ��^� ���٪����u ��R�J�c������"z��������/���\�NgҞ�7ߠ_��_�ô�1��ۗ��ᇰ-�����Q��G�i^�$��t�n��:d��21� ���&�sG�B���O>I_��:)2==��7MG�UEP��֘����s�����Y�1�{:�l�,�?I��Eګc�3P+{qgj)�=c#���m���P�F,6c6"�0���B�G&�-30���Թt�h8N?��H� 8��~��{T5�.��a��T�Q<�T��Y����@�3rQ�=��*
)���q��ymgB#_?JCA�
�����z���l��7�z�׃�X�.�jFɼŞ�3Q�1I%�����I�]���᤯4�=�ST:|T�a��߫k�q�4���OEf��������~�b�m�7i&t�%�z�~��'��h�v-����W�����VP>N]Q����XM1]O�8Y�����K�W�n*�7Z�Ծ����_�80�f�n�gz�m������`�I��G�z��O}��+W+WMǓ�iNf��h6ܝ���c�߇z#uB}�[���~�' ��o}�[��ַ��k��oQ�x�{��S�ﺬ�����y��{W{����=���]�F�Ni��]�8�:"7H�yc��I9
���b�4�JI������z+V�vZ�q�?�����oU�vY��]U�M|�~h�����z�xӶ
&" \	�)ؚ�,D�kl��*��-˗ǀS���G��~��[&�]w�2��Bֺf�� �f%Dҟv)����Ԭ[	��qpP���²z��1�ZZ.N�����z(��@)�
��#����|� c+�CC�i��,�(�hp?�"]��#�n��\�y:��o�߿M=���pr���d<��F�cS�1,�a5�@H�_��~�._����A}�k\���xr�fP#�]<~Q�����ѐ���>�`Pi�֚b+����"!�<�����ͷp�y�&�|��Fɂ�>n �(V����+ d�������eT.P5	`�	�+� rȏ=���o�V�W.����*����9��#�s�N�3������:::���/@������~����� ���֕�N�9ơB�[5��:�UN r|M�t������>��}_m�G�7js��� ����ߣ���dNw��h��������G����Q���<4Y�\�e [�$Kа����L�20��=4�����Ǟ~��<p)�����\���!�N�t��Y�1�6�W^��������]�|�Ν;�s��� �������.U��kdIl*W�@K�A|5LV�2%��՟T��0�U�ɚ����ޣ��ܜٸH����Ue�B�������߁����,kRVA���2[H�
�9�����Ņ��Q��L-@�7���,Vp�� ��q�,��,��fP]���fg���[܏�fxf�=nA]��N��%2�*ǣ��֯V��@�ܯ�߻��+r�݉�SgX������X�Q�?$�Sh��?a�8�N8]�<��;�j@��<�ڝ�g�:�`$�'+y=6�+9�֍�z�ύ�F��|_�6��+���17p�2*�?� ��tx�k;�Y.�4)���s���aEg����?G����`o�nܸK}��4�B�� ������o~��q�������Ξ;K�'_�kyTt�a
27CZ�eܬ�FTrb�L!��W��t��U�ؠ:�p	Ѯ�����C
�@Ba5">��ڴ�f�2'6�0���_A�f'��dH�,���=�,Jz�eYt��QG+�� ��I'S�p�<ҘOs�u�:��t�7�B��qO�9��w�`�2���҃�ڏ�ɛP�9��Zr5�+��%�D1����H��9?��ґ�()[�yɫ�߁�<`*��j0P�YG�����KT�G�v��5TvzN�r�~������T2ݔ9Pr*
AJ���6lNY�m-;���i)�ڲx�G�B������.��o<�e���N�y��^J#x%�,�zu���?������E���Oz���g�=��5I�
����O�=��sy�7^�3jYu�gD�:�|�����կ�*�S�w �L���d7�����矢�����e�o���kR:�Q����Q��3i?��/H���9-�Aن6ɞx�	MU�'��3�]|���ؙg�k�%�d��w\4�����c�1��!B�� ��3ͳ�S�OU�"� Hs�3��fC�JԼ���e�e��3��t���>���2��d8gJ��J��'['c̄�L,�!+�����gK}2��]��R��
HtH�xަ����E��Y�(x�V�1�i1�:F�GXkE�-�zW�u�Z�+kiD�F�I1oxZ��f�e�˞�����Ğ�H�T+�R�R'�<L�L��3�M{�J�!y�[Vnv
T���x�>/ed����D�\��Ō^D�ن�.��0�)
��Z��qc�]ɌuB#9�U�U����,�����t����h�V�E����ޙ������W���7S�L�V{%����o^�	 }�[��ַ���o�_����u��������߮^=w����nծW�.�+�����5��:@�w%���0Lf�(h�Uce�$T�fmBzU%&-��	E��(�� g�W�M|�dUm�J��\�AV��V����z�����w��:g:��,��׽i�V���0]�xY$�+��v�^���s����T���h�(%�J
�5,�,pg���?�=����׮э�7�G�g���c�%�Y:`]z}�\ ��L8�����=J�����Ե�Ң<,^2�`��>�� �Ad����;�#"Ɇ���fb�#+��Q� �\���iUXn8����9���Hm��V?	��q�����,% f6VWV��9�No��bF{�c��Oq��T�d�MvG4=9L��H�ʲ�%���ݽ{���4���{	nz � ���=@(�C~��9��¦`M�D�1sP��ģ.�j��E��c��doL�� Y���5��1�Q@�u�^�����]�k|����=��B�C��V��5�l=�u�A��&?�0��F��r(��\3K(k��dG������>A'''���M�=����!k��<�cp���?��ZO㑌��t��wJ硔1[��=co��'�i.�B�|�Oi4��t6E�#�-�Gج٦[�.��Q@|��RHZ��>��d�+�ݛ`L���>�Kp�O���&]�Ši�'�w�5�!��ж�����d^���@�OW,�ͥW6"�͸�`��	�5�A`Q9\.���U��\Up۔����.T�	�}�*OM[-����K�����u��k�gJ[���,d�����&�LT����ۭ9b߳{)s�������Hr: �\�^�s�P.h�%� ;P5�m��5��Q;P�R�C��6+����C!�0�NA�A� aBg��\�w|���d���L6����Ν?��^�j���7nҍ{w�_�"��`=���97�_|I�k���^�����|~�?k� �t�/S��@R_I�^�m#R�t'���3۹���B$�X&� :NǾ	.����ද�B����杁���o#�A��i�>���=���o���@�n����Z�k�@�D����m:w�ϠU�X����K�REBr�����������y��l�g��~�'�p����x�\E���-@�
>��%������K�v����i���{'�W������q^kL-}�*���=���읡��}�{xH?�(��ƫt���q��tй�CY�?ﲯ�:���M���������6�JkY�0�!�z����~��S���6�i\ɾ��O��eԽuǎ�|�S���?���PӀBO�?V��������y����֟~�^}�:Ns���?��~�����i���I�+_����*pc2��M2��'�~�'�V��ƢX����޷%�q���_����e_ ��U5J�w>>��ٷ��e��g	���P�NDB�)��4V�I�
=����J�1�)x ܼ��j��^WW9�|J�����*YY\?�H�i�������G��IT�lm���}0��k�/�H7o�N��%�6��𞚷,�èx:�l�Oo$�J
���;��"ÊIB���D��.�'���*�Z�����KY�AJ�/�b��lj?�&H�Lb����m��_��Q���gX���T�.2��/^�#C�G�"�/,A�Pu�hĀ(�0���iLX3��Uӵ�̬��*\k>���'?D%[H�
a�9����l���Q���{��R�����J��9e1GW�&�'c�ɽl��.6���'ӣ�;�U��'��x^�Q��ַ��w�	 }�[��ַ���o}���E����qm�~=NO�'ՠ^�f�r�J�d�����\�[�\"YA�h��؀D'�LRBZ2��q��_@FҠ����y����Z2 K�G��K��f�T� ���C��QQ ��:��4����j�"kz�X�b>G��������LpH�6]p�m�9��`��~e09�9�%��(<s�,����,�N�{�2!��I@��EF� g�[2��X2H|B���������s�z�l������K �e�Mv;�_��3���$楯9����%�3H%Snw�@�%�{gP������\f�ZlI�R	h�v���N�]�<���tQ�:��o5������f���l�>P�Z��Z�Ym#p_d�ҵ�E�x[`R�|e�!�Yxn�T�������rQ�ЍQ�/�\`I]!u4r@UKD	F/`�6������Z7�ٽz��)�����M�:�nx��
,q/5�蝦q>؟���׾VbFB���4���������E&s����'
VIx
��!�Jjmz��g����?ŋ�}�)��'>�`9����� മ=f�%���d�o޸A���4=��ô����߫hQ&���l:��E����%��N���2�c3ԟ���s�Z�5`n��:�"]ۣ�>J��޳2�A	)�!,�^32T���p��3���`�zk;ҋ5F%Ϲ>qk5��I�k���Hp0�- ����g^��<�X���ߕ�G�[��&�n���x� {+�)��V/� �P◙8�,�bj�G+2a�����L*d���NN�k�5#�Z�]�,S��[c�ig�Bȟ�� :�&�뾨��E
��3 ��e�붮����U��
��;�A�ME%%D�y^��l_�;��a2�t:�UZS���ߤ�����+�z���ׯ_�+W/ӧ>�Iz�����hJ������ǟ������g^{�:�)�r�Y�w�߆�9��ݻ�@(��H��
�
��R���͕i��4����8�����t��dX�5����"P��(��4J�����u�3 $*Z�1�c�s�	����>&�D���|��Y����7��$�	'���c_�F���� ݾ��Ʉn��ʦ�:�NJ;�(h��+NM��7&?񾆕\G��^�J���I|� �<F�t.^�׋%�����~F��i=m�%5nC����z��v�WX����aO�i�W�y϶�{�G~2�s�Hq3�0=��cB�"�~��z^^�`���IJ��k沚�����P^�3~)�=J8�6vA�AUH��(WC�����}H�����U=J�]��c�^\K���h��;3b%�2��e��o�Ï=J�'~<�c5����Ҿ�~��d�ޛI���W;��o}'��#��"��{^�kn�>�n�_�k��a��E��l|�7�Z��o}��x��gy$�� ��"	����z��sZB�����2�3)i��� �e	�_Q�l@k�M�F��M�,�;d��Kc^t��Q���oQ"��9���Z�j<_y���&Z���4 �����8����������p�k��_�ɍ[��͊��R��m�U_h>��e�n�L��y�ֵ��=3l;4�gx6���$��>Q�	c���*_��*{y���#R[QI�r�dQ�iz�N�ݲ�UY�F~��ABt^�$��D�hC���ix6�!?[��֤>�,�(��VJd��� ��C!N�
��a��OV�N���E
Qm [�3!��'����l�#ND]�Z�,@�w�YL��:�Ӟ~�����w�i7�Y�����'���>�S�&�Wf��'�|�WU|'}� �������o}{�� �ַ���o}�[��ַH�2
�n���NC՜F��*�,W� �;	�K�e�|])io��[Y0>g2��~V�I�i-��w���Q�؀��-5VU*W#]Z=��A���he���EZ9�ÁJ��} `�q�R�Z�u�7��b� 8K3�2������7P��$��DjpOk����9 �97�
AM�wIP�����������kƇIc��� RD0>�l�
�g��>�'��_�2;������� �I���! i�(A��P��m�����j]R�$�`'��Vp�����VP!3�i[�[H//�+ �k��e]` ����}�r�l/N���u�P� R���7�J��!�
�����^G�z
 �D�˦�i݊ �DM,��Y%��io�O��|!��4Xϗ��j��i�D�w�D�z�Qn�m�M�G"{�6ș��}�DD6�9�����ƛ�_�|�N�S��f� 

��������@�c�6������z���{t��Y�(��4�4n#
齰I�7� �x "/|n+{R��N���E'�� {��oYc�	+�B�K6�� ��zs��o]���_�7��+��fr�-��#+J�ϚI?"%{={���O�_:O�z` )�ch`C;�]}�2�������S:��1�$�՞��F$����F	+ �d>�+��g�)�3��u��lU�Q%Ë1�5sшP��m�vΤ�U���ri�F�}���zG�#9�NHV��*���a���W���
��D���H+� �FI���!�Ȥ/9^8���ϖ��ftd����-�Q?W 8�f����v-��9��+��ƌ��3�.p\� >��#v�+�[�=�R�+q�D���2� �M��ɤV�Q�r��0��@�����+�1B��9�c�X,ᏚM2+�$���3������w�^y�^�?�O���KtxxL_���h?����]��?�:������G���o�C��Sz����g/�L}�c������g���g��ߦݝ}��ɿӛo�N���Nw�����J��X��ԇHɄ��T�6g\�S��e��@ �5B�~p�T����r�����هQ$�i!@�:�a~ԃ�~NA��#d	3�����4��A����Q��/r_ K:�ڑTe��6.izx��hL��>��5���ѝ�8��[7�/�]K׼L������յXT@ؿ󹆬��ZA������o���u�?�X��D���J3����P���h5�ә�gh��֢�V-q]�0��є�IV�c�p���$���3ߥ+/$�:D\��~z�.NS���^lÄ�({��7(�M�\�f���:f+m�dB;*,�/\6[��'��F��e=��Fh������j�Ca�i���';u�����g�^DT��Z��'��;����Ghr�<�6�ۢY��^mW�f�'�������+84��'�6+uܽ{H�����5r	G��JW���p��������/�
�1�e�摙�k�tz
ۜ&;�w���!��1z�Q�T��91��_L{�e�wOp�Q��fMC?�=�E�/g�k��{�M��H�3 W��ԒIa������>�m��U.��<�w��U �E�!���u5:!���W��˕�d������ �s�
�w�"�<��@��z�U��ou�ײ��Ge�HחJ���d ��糯�������a�G��9����F�{� ��7�{��B.���A�H�2PBt��%/d*/�m�������g����&���RΞkU���j/���%�/9�)��Z�a��B.�Ս��\�� ~�;�/�QW����bkL��D�J��++qA[S\��ZDD�<�3Qw��%��,i�k��Y�M`U5<�3���<L�f�<���;i/x}</��l\_�o}����� з���o}�[��ַ�}��W�M!�?�Z�9�"��8������|�x�J^�r�����d�m�#*2��@��3��I.���M�t��+Cd���׌�����z�Z�� ��&�Ax+ ��?1F��t6|���7�3 �>Wh8��dL��Mz���M��
j �b���� 0��t�P��gP�2*����s�C�����&�J�N@=�5��M@F^���$@� q:�7r�!#�rF�����Noܠ������Vo�
UJ�Y �좖��1�=����G?Lao�˗à��,=��i9_hG,������D��"�)�d�G)�����:]���6��>�K�s�;:!Ip|�˿OO?��ƸF��)X���!�(pMx�+����
�@��lp��9��B#�ޚ�{�{�6M���MD�Ed4��gEgʥ�������d�E���@��tJӓ)�u<���A���.�ə�a���hz�TE��^z}:]����{�{ ��;W���� �ǟ\��%�Ma'P/��O��7���|�V	�n��dQkVl�-�^�� �]H�*�4�R��U�@�}���L8��#��ޤ�^�>Y� ��=���h �rr|��pF�y�O��K����o���r����#�P�s�.��}�=�G'�c(��·9׈JE�n;��k�8X�wE���~��:f�ӡ��Z}�6Q����E:p]b�M�� �V�%m;YA�@	�cs}�JUXZ+ �'���a٩�a��ޙ�h���uΎaEq��a����C0I������	�z��@�0_\@��G2�Q�l�Qɤ�}f�5w�58U KQ+[�3s?t��u΋�!(a����q?�g3�|�Y�*�u�,���\̅�ʑ(dU��>���G>J7nަk�^ǚ������� �{�7�-Ng���oү�گ��������3������}7ɸb>�f��j5��έ�����qk�>U愈!�����Q,� Zmd/�|V��9L�#��9�d�{.Su�"w&���rU��.�'>
� w���(��rdň�@�JU�D��f�Q�p�p���|�ѰJ:m���U���4��w�A�x8끔��Z�b�ֲ���4��V���r5�!���6� ]K��9N$�q���ɧ��O���{����O�������N����}��>�U�xb����9����.�?�݅� _�p��l���������O�>�Ǽ�-{��g5�'+�R��I�?�ry�� ��u[���&�&pJg���t�;s�Z�;��~Z&B���c��/���Y��0ͷ_��_�����A�����'���J�Ν���:�o�w�i���������<�邪;�N�.�<U����C��������Hgh���&Gn �)F�t|��g�O��������k|���ͬ������u�O���:���[71��J7�����Z���;oҷ���5�Ϟ;K�n���{���tm����ry}�O(�X�l�K�|g�(�Q��g#ߑ��g%% �6z�ZI�Btͪ0�;Qy�J�q%N
� ���5�^�)q� ��%$�q����9]ls!��r=�*�ޓ�_R?�g� H���@����Z"d�F�Ik�X)�rɌ|��|EA��=�PԠ&�l�	L>��&��֕�'��	i��{[5�L!{
�D�L=��}�=EeD!#
�}2ּ�%�H��!o�Hm%�g�0OV�'jr�˝�%�^����!�J�#��mjc �ً��H�cc��<[�]y��\����L��i�q:�~��_g'|H}�[���紞 з���o}�[��ַ�} [řXM�>Hp��%
vd`~�XLn��r��YX�^w[ 
 ��&��z�WA�V�� ���d��|��8��Y�|
����A�f�b9$�j>����m�O��{�	�ݐV�;�����9	tJ��@���}��ߥׯ]C 2K�v��A@p-$��X���J׺�y���2�����0�L:�3�9;,j��y�u �<��0����a#:qT8wv& ���$4��Y�A�p����7���!���������qv(���!j��RiM���4�bbA�l��^y���c"��·Y�3� B@z E�!�7��{PsJs�Wu�_��z�����4��u�%�Q�`��`u��p>+ ��!*�7�79;��1Zd4��6P�8�r�嚐��fh�����h��R�\D �B���$Q�`�n+΢c���k��I7v��m�: Ovu�ƒF<�Hv���i~:���V)g��v�Sٶ�ǁ6�U�� �ξ�*�-�MǺ�ٰ�����F�٠�s+���b��.v�rw �NPQJ�O��
v(��)}l&Q���H �өo�����Ig�Y��p�ٻ�۹����39�i�;����Ð섉-�o��2������Kc�9�0�cz|��V� E��N��Z�k�Z�D]Ix�C	d�~5�H���d������;ZJD��h5��f��b+V���IV��焸�vƵv$1�A��k٬�xa+`>�X[&b��oK 1a�^�3HcЌxL��Od�1_o��|+��!P��L�l}��ť��#�r��l��_w^�"���5����V�CA�d�P�Z�m�ٜ�{eIyV٨�b��`0�Y�Pg����	�`+��f4�/�o��;o�;o�I_�ʿ\��D-�b /՛�`���ݧ�ޠV1g�{!@,S���U�BF]u�aP�ђ9��L9���}�S z�Orgn�$��RW<�R�z5���#�=b�<��d�x�|�㟦z8�M�˶֛��؃�y�](*��e5�B003��K�x2ʡ�S食���~M��L���GR�=��O�4����d�UJt�x���2�%=pmB�4��҃W@cr��Yd?;��H�w(Q���98Kz�c�0�,}b�@7��W�__x�!z�'rIV1`b���
%}����S��_O���<�x�e=d �I)��d=��B��Lw+ed���R�G'Y,s��w��2�>���mQq� ���MRN�= �f"H���:�>�T)�>=2��Z׭\@�l{�0_ J+ⳙ��I{��>�L��4��`4�8��c��X̓�~��RT�6R��:���Kv7����z�~��GW�>���D�z �;WY�W��(4�*��H�+dP��DG�����;�e�'	�TJ>QV���N�i����~D\&m��1?��������	�9��f���i.���"�7���Kޯ��AY�U!�_�u�d�h�(�$�+{�@*���J�8|U2�Ym���c����d�הF�xu}J��OT����FBXs�L���B-���t�kⱩHI����cu�� ����`����]�n��е��m9#�P�JQ	���Q��<;��옟Kl<��T?��_���/��I�D��k)
������>Ub�N`}�Cyz%m����G����H	r|��]oL!(����N�r�U��Z�_�V�ϒ �� ��tưq�>"���z�>�������.��^��ַK�D��ַ���o}�[���k.5�9l�9���:y�������s�R��Q�qh�L��f�p NQ��R���9��`����h��^|��ܺ�`��Y59���F�`��o��Χ�2�}pp���I��!�/� *\��C6"�O��5,KZ���G_�ݽ{[e�%�"��IȢ���W�^z�y0�����!=��O����[F4,�L&���z_���j�)�� o_���,0���ɔ�^y r��t=|^s���ߡ_|�^z�ez��(��HL߽{�ΛM�����rm&D�j�OH���O���񫯼���e5���~�nܾC����|v ��fݤ���4�R���~0�k<N�'t�7�9�`�r%5hG�:��B�|��f~mF�c�Wp�FCɸO68���k����"]۲�̳�-�'��鼧 Y��y��o��M�\���:��hD@�g'�nB�n�>;� sv0��-$X�W���2��&��_�W_��g�I߫���5���ǒ��E��,�@"C̒�B�7��� `8F�Zq��5�N������5��`'��$Ά�\G9����(N�,m�P@4*Y���i y�
�k53��m�pX�UΜUv���^CP��� �r^�Ro1�,y;�;wn���1�j�Z�8������� ��w��n�.��,K �����c�s� �m�2��x���B�P�y�D��������Ջ
B18lj%��G�u���>Z3Ye#���^sFyU���lz���.�{�s`��+��0�Ǹ�l��9�bQ��ؕ����+Ewc1���)���ם�!c����q �k����ӣ2����}���]�;l/��w�n���J�N0��&�\��@�Zg��_~��]�F��݃m3�kt3�L�:=���_�uz������txtW���l3&��HCYEc��)
��+���$Ѥ1�����ٶ+�}��nY/�J3���*���tT.<�����l�L�H^�q���-����1�d�'i�o���� �d����7Y��(�\�Gi� �6���%HM���k[F� �\E�u9���Q��>�
��M�QA��ە����B�j gh3��hF�h2�:�L�f�;�BM'��#+ɏ�.�N�u2�Ah������+ �a�A�pB�0-8[WUX��Y���u
9�|�������� �`�|� Bi�1N��,�Qajh9%�� �nwI`Fp Z:�IP2��o�(2�z�,+O����kE��sG�Pc��G����� �D��<�d�C}#}�Ғ(J𲈌i%s�i�ޤ=�:��p3��`o�_nVU��rE J��Pk���~��{��6�����3�͘�� >c�L���Q���#�M��0��d������s��T�T��-��P7��ԓ�j1яD=�άBJ�����_�:�a{��L�ļt��x&~��@��������g27#�S)OVg�,����&�0qg4�0���}H��|��2M1��=�m�+���(�3�/���Gv0�,�&�+2�r,�6ƫa�? �O��~�Zr�}p���ץ�FZ�9Λ�Қ��C._Arݱ�� �I�)� �՚L���B�[�E�k�+�{��b.MK�~Oe$p��<�9PYk��m%�(*\�QR���a���F4�Ty ?��X�z����]�Lm���$R��Vs�\+4��aD��nq�\��f�z`�W]ٽ���o}{�� �ַ���o}�[��ַXc C�!�J#90&�Ě�N
(Q��,�!	2d�gʕ��,�S�oz�.?@�٩) 8����\��ݻ���Z�6J�_*��4�m3�,�C��!�J�ɮS���p�bi��ɻ�K���ǡ�5j#���kt��m	�F˶�{k��1�ȑ>���w���^|	��%��kd�#�:�����h��B�u�_%�m����'"-Z9��w��~�����.��-{q���dr�}��ZRr���(H$�e5��6�9�����0�
i�_Iv�Ȅn@��{9�ە��"1�� �gz���%�������I�:O珨���,(ih`�ea��c���U�[�~Γ���S���D��F��'�x2ַnߦ�����?���Q�VrsI?�!�N�fr���C������1@�{��n߾�Pwn�@���p8�C�ȸGΞ����&����h���r� ��k5/��a��0*�>9|�A�û�i���mD ���$�a���C�  *�T'������<Ape!��և����M��gh�j���%QW E���fl
 ����4h˟`:�m=˙��䪝����� %���L.y�Y�d��_P@��-hJ�N}�5e��\R".�EpIa�N�6X�������н{�R�7�Ĩ~�A��f��(��~��Q<��K����Nk�s4f��d,�����V��-B�ޤ���Z���^�9ۭ2(�1��hiQp�R�>B�`��g�ڝ����l�t$I�W���i�N?�'�/� ��,�|ߙ<���
�29��z�{;W.�˘t�
��M(�"QE� C_Hi�p�:�i�X�\���.� 7VC��˿�K?��Rr#P�h$]  ��IDATZ��Ѭ;�+� �!���\��(�[���MXg���`ïdr��xS,� �`��1�f���\re?@VB�I�Pte�]��mI B[�;]7�֗\*��+��G�?�J��������Z��Jw�����<�*-��%ș-�z�Ԯ�,��� ^r�������Z�Ȟ ��w ��ҋ���I����k��ZUpBQR�LR����
R5J��)��x�����R�����}�T�yg�;/��HH�A"�$��u�������q�}��3Y����U��5���5�S�΂&}fs�|��{���C�r����Z�p4�~��~w��qMx��4i�T�GCf5�z�2Zi�w�ɱr(�w��쯂��m볯St
L  �5��������#�`�(U�PK�GU�i!☡ѵZ�K�ۮ`�ڒ��Z�2��?h��^���^�RP�E�v�u%��D����	���[y����Q�%�B���۝5!7���ㅓT�9x�r�F
ǭ����0%�ٿI��B������~��Z ��F��&��/\���3R���c���� ���;�?��л*��_1���xΚ��Z�����죔(�*K�J��pU��~#cl坺�<�D����Y
}�*N����˲	�1��y��[��S)�Ķ���P�P;� ���GY5U�"!#6z,^���]�����g:�N�I16y��g���s"���+�Lf�����}yS:he��L�&�糈yϳAr}�nà���p'0E%֝E�o}�[�ާ�����o}�[��ַ�����]U.b�jʲ�ܼ�r��d�+��ng�d����_�5N������C�P�m��v�A|��J4܂�-� S5�D����aIJH>vA¨��w"�8�nhvr�A9����~�vd�9H�u*�_lZ.��(S��K�sQ ��JD�x�o!*�B�	��CX�@3�J\/w4�`�&��t��u$@��f��� .K�#{�2�EJ��G��{�>���C���X!k���d�PVА��9C噧��@�L��3��jF�K��L4d��"�6 t�V�O��ߣ��I�;�[U�����+��K��G��^{��|���٥�����]Q��)P"���1��_�2}�_I}[��34_�����f�5�N��>�w���*B�A��,W��Z�l�-~]{�r��aop�͒��q%=�D�� 9�f�z�\���V�T�)��)_B����|B��۫��zr]����`� d�.Qs�5�G��9ۊo�`�	$ ��C�1���kv[ ��	�V��|.�W�-��נr0��m�`n䛀�})0n-sϳ� Q��NI��6+&L,4XK�[}�dv2��_d�� �T.�;��v��N[�7u� ��/dBnZ|[�<��tH����	��L��*�� �v�T��L!�hF*`b�Ѓ����?2�c�5�e�4�l��8b�Czb������}@����q����Xrnq�,2�T����}[����A�������N�"�Uf&�u�����D�'-�Q�qf".?���z���r�|���|.�'s��2���!� w����IF��e��U{�,O��� �m|0�^6J��p���촹�U�1���̈́"2����T 2��i�c3D�kT��1|-��l*7����TT�d_"���R0~ I�� ��� �+jEV ڵ+P* Y�i�9�-�(��^�����$��T�(�� Y�c �o#�˖����	(g ��L�y�rK��=#'�>�����P�`~��ꦰ�k��v�c0&o�x�8�Y���EYB��T��0�[iu��~)���D?B��1Tqw��_R�7y��ߩa�_�v�A4p"G�U��������,��{�<�<�����;���<��];��a�pe��G��|{kQ`؄V���T�='��M>G�YN�*�s�D�*v���sH��tU��e}��8��.�H#	�*�k����m�+�������uÏ;��ǵ�窪3��̿<�J$%���V�l��I_WA��X�Wꄌ1��0Ԉ�@i��wD[�U}�d�fu��d�;X�}�2kV}P���{p&7 ���V�**�V��D��V2A>�����J�02:Q�j��S�O����UUFtBSe�B��Ω����1�g�e�@� ��@��0�+j�M�?�¾�<T�d�
]f�Tʢ�w�v��, ������p�6&��`3	YE���]a�h�6��\y�E!%b�b HV͚J	'��G-qCN�J���,�?�gPM�Z^
l�����,"�i��?�ѧX���2b�\m'G�G��v&wc����ַ����[O �[��ַ���o}�[�>`� \͑V_^�X$@X�4f���!�i�M���Y ����of�!.2���h�i:���?���-�G��������6t���v{
"�ϒ�RGZ�ќՋ�lL��ԫ��/�K'  �v�;�/5��:Љ�.�x��\Ҁ|����Ϥ )�+�(8�@*Q��%���}ɰ��FAі�luq6mh�nh�`�.^��L�1�E�c�P��ȈK}P�t�ٳg����(#0j�ns0ues��g*�b���  >����Kt�z�bp,KGS���D@�9�0�s��;we'�$����\����L}���`!��C=H�ԯ�)tx|H7n� �p�qL>�����    Һ�j�Z�v�l�0��k�u,[ �Hk�w�?�����Nˎ*�����bk( F�A݊��+�WH�KйN���!$'UE�yhkAs�e�%����.��͌Xj���f��2�@#����
���L@��엁��:��S�� ��e�LR)]���$�[X��� ���b� 4+j�!&���}"�E��2� �@'s��J�X2�M>^?��/��-�]!�P>�Y�|<��K��u�[;�S��V��`=�դ1�G~D��b����I=�e2�A����m�2ֹ:����m����E��ؑ��E��eFE�Hds�A����E��&�L�nvm�=M��-�K�f��ߥ4Q:G$���f#�L�$룩� ر"-�  �s"��?�^yM������/��uO���u6Ȝ��p���m-�>�tͶ�30I��s�Dy�t��wd,�FWz����Ȭ�ɥ���ci������[H��(�	J� ��,[���鬫�:ر�� ��,ǎ���T9z���2��BtYx0����2M��%_A���ƀhT�C�G���6^PYtZ�ň@��q�=�5\KGT��L	A��'���HM6+*,�}���� !ȱ��A�2ܴY���6vF�Q'��-����#�)h�B6rjx΋b�C�dQd+K�8��B�����y�X�n^k!��5/%�S� �/�(dm�`�d���x�d�.��9-9�#�N��^�tm(�:
+��ʸ�����x��J�z]]�CTTf�^F峄|����*�/v�3`΅���/�#ci�R���jv[{&���:�Z&��B�nP^�nܼ�d�uK���� ݼuey��1ZP��Lo��A��|�#�}8�+V��/ ,oZ!��;�E���j��z�Yc9|��g�kQ��"�RA���k�֚�����.O�ʻ ^��A��e��(JY��֙�1��:JF�HF>t!�r/V�(���������/������' ɯ�Am������JKfq߲�3cP8`U'��*�9)w2�5�����J�2e�t)L̵g"&2{W�_��.2�I+y���N�?xO�J����,/>$��)pmF��ݸ}�]�����\}\=l�j�P5<����Nv&o�Cߪۖ	 ��o}�۟�z@��ַ���o}�[���AkK�!��sqK�A�ؚ}Qd��ucm.�V�e�n���,�8��_5� Y:^�Q� -�4��e+m��s�9Hr9s����@I��4�=-tj��*��lgqF�o�Jd�/��8���$0�k�6n2*q�f�����Fn�s2��IU�,�v�p��[�T�9	JI�Z��#-Kz���8d5��h"2�T2zYm`2�����ɔ6��N�M�'�;�N��݌g��,�c�ˁ�a1��r�>r� �k�
BD�,5���\l���}=�����>�{.S��y���6;B9G+��_,p��b����t������@�:�"�*Aܰn�b���X!R�ٹU�꼐��d�J �U-�I��`H�}�s���G��$��\l�~��8�g�w~o:�����	����=���(��BAdg[�Elj�D�<^�7
�h���Ҋ�y�s"���ST������ݸ��
�e>�|�2�! ~���L�z��+`J���fY�fcfo�67g�i�o	��B�v�JM��/Y�&?_��e���T?�AAؕeX*hE�S���̶8e!y���KF�H�s�m�B],D�/X R�V�]�0+;���Y��YMf#s(Ģo�ˌլ�q���E=�7?L�LLe� n�y9�8`4���z%F���h��H����m~�w?�P��u7� �[si�^f���ɱ3�[�����@�*DU
	��2��������c;͚6�Cw����N�o�dQG�=O�˾@�g�����{e���sk�� ��#�G��j-4t�%^e�ֆ&�W����M�����a�mR�<���-gie0�*+tH,�{�랎�/{�Yؐ�-�֬S��1n��^���7K��iU�Z[wm�+8��:��ʚ+E�i��{zL�)��0�&ۀ�}L4�V�/��:}��ON	���3b�{�X��L6�1s;o��2)��6 ���y�ޚ\�M6�|`��*��cI�S�|j�pZzWS�/�C��hv�i�j�]��ky��y-���$U0�T�DB�O���h*f����
N�f�{{�ge_k~-�Q��55 S�����e�;ү�H�3 n6`k~鎲7��mݑ���O�2��#�y��0�ק��%!o������u��%�ƣ�W�`2���Θv��P*��x����A��h<��Ѐ�ӺF6;+p����`�}��V�H�,L �};�0V'b��=�:��l�L��� �6x.��(��r�.��k���f8.�q��'-�ZS�nZ��*R���"������
i�Rc�C�q�zKr�\��q��������bd�֦)aO#�@V1KǪ�i���y�R3��*��>wP�:0`�`�"���V����TR�B��$e;��Y���D!@��lɭީ�N���f%s�ҵ��B����F����(؟�?B9!�[]�~ �(�oQ�������P�8�y�Y��hZ3u5�gΜ�\y����gV\���UZoV�e���$�&V�ԓ1 �sK�[��ַ�� �ַ���o}�[��ַX�꿮���N,sH2|I{]p?�$�8r&0u�Z ����Xju	lF�D�Kp��	;��d�Y;�f�[�#�<t��kA^@v����{0�X���U�H���u��� X����Xip!�@CO� ��3�8��SH���r/�����有�]A��r�]�+�+z!D���c�\���}�nݺI'�)�Y����zX#�i4�ָd	��>�9�s�&MX��jUj��@TSW�����{�tL%��)����Q���rEs��龜b�mۀ�fzo�^�|��ҥ�t��yd�/�����	0�S���r�F�b�մ�X���իt�ޑʱ
`� �J���i��S�`�d絭��u
�a���p; �52��M�g�y���vi�ȣ1������K48��������7�@��)m�-��|��"�U�4@���x��)��w��:�u��޲�:&�%J=W�����A�:cHJ��a+,��58AG\����7$��%������K>�Ɂ@
Q� �}��D�k�� D�Q�ͅtrL&�̕ �z��>�wːF@���
���qp���3�10<'�5�w3�-[�#CH
���uU#����|,�����Į��I)5�(�o��zRҢ��s�0�2�O����m)8��qۇw;6�P��������ؖ�KF��lm{�&�v�5e#�xk�����|Ȟ�3i.OS�6@�X�%!
��)KwT/>��e�f�F��/DS(6���%i�nR�����P,�NB�(&D�W8�~7�X�!�n�Z��R?-k>ng�����L���}��sQ�� ��<�΋2l�i���_�"�:׏�xn�8|�J�ޫ��|���{=�M�J�͋�:��ѱ^<���#�$�W��k��<�|$c�aO`ko���)]�����"��2�����t��7ܳ����H�GUo9JAm�v�OAHB�(@A�%��K?��{� f�����ӎ=(Q@��2�e�U��/�ʍ�q\�'nM��F�[d��mWRn�]÷V(a }%�
kl��-��A	M��UΑ�,l~�b�m�{ ��?��:�����B����w��?��bՈX6l���HwB8���4��:ߢ��:���\琨��+��Se/�X���q
�l:h��}�e��đ�\�\'S�Ί���ٵ���+���u�ڮ�fz����ɂ���"�8��vF-b}���Wmk�Ls�9��3Q�����x/ΪV��	���� �]L.>w�<�n��>�%@�H��׆�si폣�(�9�:{��4����N�~�G�Y���$���G���`GA�>]?kR�p�� �ї�-��y4|�aW�!����&�:���:c�Q$1'�m;�Vb��0�kՙ�-��y+W���C"���A�Gy���m7�$�Fq�b��D�m�9Q
�T�"�cGvm8�Ȇp�.���TU���y	���|�>�]Z��_���i��c����,B,FM���]ޠ�k��=�߷�����z@��ַ���o}�[���k�T.���j@�u \��T2���/�A-�2X���*BI�5�A��ZH7˖v��ܺY�۟�,�	Z���*#��I �4�:��"5�	�[�1Q��	w�ILꂝd�X:Ko��)$��@z% ��-x�2��2����,�mݯ�t�;D&�J�W�NU�ۜᆠ�ܧ7�北yZ�=���顇��_���S��Ξ;C�/_E6�|6��.���V���ϝݣw�~��5;� .��~od�0Q�F� Y���ؒ��4�-�uJf	
@!0��,M�)�RN��@�pX#X_*���~�O��	ƌ�������;����4��B��ݽ}�4-��(��1F~ @�=��Wc�:�5��r�Ω���kd���g52�<�>Kͷ͌�ӥ����>Ϡ�j��V4�A���!{<;��lA����:�Ƭ���Fj����9���z �z�P�q�Hq��5�d��drm��(B�E@4�n%s��p
`�T�v4@�6 C.hֿ��,-�RI�x�d0,�ʊ\���rp��$rR������(�)�e�]�^'Y�2VP�@���<��d�������Gde
ؓe�M�_K�s]p�dϝ�2s-�Yi�Fe��7[Q�����V+7�a��QW:<�����jd�j�!�<���(i�ep����n�f��*�,��@�Vq�2j+����G�e���@���}�����z�� I��ρ��u�������)�->_�N|:���a�;�P�=��m}�lH ��(��^(H�5��9��� �_�s-l!��xߧ@6��'�>�ա�~N�� ^H�$��$15+b����v����� h wC�S��\;��L(D��E�5	U5V�fb�М�4�T���՗�s��۵�|�Gf����#�~WYh����R����L��!��Pc���yk!����������CnAW:enb�t)��������i�)o��X���X�W0���W��M���yx|2�TJ�8�g\�BYZ��ޣ*�t� �46�E�B������-*@]�����M��u\��}2�7
Ћ��iN�;�:��UY��o���TV��`����%���i#���y��K��!�9@5!B6�ɠrG�*��<nx_!r�71��$#�ؚ�;���v�x�V�/j���m�Ȼ�an
Y�w�{�M���to��s�'���Wz�A#��~Nx�N=���Ul�H B���:��y��,��C&�:�}}�z]�n�=
ż�c ��ҏ$��Y�
��Dj�~V/Q'm��>����I>�����J7��+�1�W�{���y"�3J�D�t����R�Xp�¹�#����O�Ŀ���G�za0�XWխ���'�S�j���(�M^��c����\�	��Woo;ߩ��O�����������\��
��-������:�{�����6�Ƌ�#��̋����?��A��5�f�m7��ԭc�Z���,=�߷���/�z@��ַ���o}�[���k�%���q����}�`�`���d�|�A�h�K�8�d1�r����ü)`�N�]��r>��k��+"��ߖ�]@��y�`u	D*��{��8����K��M��!'Y�,G�lC��X�Z=���*�޴��V��A��$:�'ƻ 쀝��G��;4h2����|���c��w��sz����8��K/���$�㏆cPz�&_�lSZ�����CĐ���`*I��;-=@��?}�� A#���â��Fl�������>:�U� ����jE������}�#��7n�̶ke-�e�ir�;%& �Tj
G}-�����0��� `�H�n���풎�'�\��/�r_L�Y��V�%��I%�0�2��^�F��,�Ӳ�m&�`���|aZ�ÛM*0G�ݝ��N��1y0J�\w�����E@e����pC�oؽ�\%� Ȟ~纮����z���`��~0H6�3()�r�г\������R��>�g�'�l������?�E�V���_fd��[������������	��V�^*�$~<J�[Q�|�<���1�,���';�kaE	���R"��~+����~�W���O�sֺ�R�kz��RҗM���(*[0�+U�g/]��nkܲ=�p�B�u�z������壮��m�5���m���l��ԙS ,cnwb�4�_�m��|���c�C����?��Z׭����;��^#vA�����e=3	���5�����s���Ґ�ϰZ���*����@�d�6����t%خ����ل
�;�kT���~N�^���4�����N�Al:��sb^lZ��1���&�;����x��e�~@��[6d�K�m�e?�b��E��=�0��Vz@��NY���lG����d��{�Xݒ�<lU������{��{`$��b�"�P�S�)
�%"ɦa(�` o�C#Oy8���XD��B��@R�����l�Gv7�ݷ�=w>��3��J��j��4�� @�{u�{�a��V���������p�Z�(� ����e��������}g�a�<��$nE�u����NL��vJ�Q$,4`�m�;�-x��5�F�j���,o<�V���{����E�}N6-`*�mW��4��e�Y��Z�Qq1[X\�����n��{���BNX{�A�ښo 0=��]�X����a������������@'�{�	#���b5T��M�^���=w�/�пq���sǲ���1�
�^�5���<���gֱ��/C��,x���@Vi���3*p���6]������P ZSWQ���ӵ^���_�����l.]B4�̥?���.h�I'�t���t �t�I'�t�I'�t�.d @��Ӏt˾)?S/�9���6Up��x��X=^�$�������
����)Sϋ 8.�(��pQt���w�ck��In�w	��s@�s�"�h�:�� P Z%@�;R���\CP� ��P2�͓+W�c�a�wv�s�����Ɠ#h�y������9���OmF�;;;����}���ɔ����I�앇٤�o館J�41��?�^�le�*��¢��D�z�e)>�����.��&����1��ݥZ�V����g����!|��ȁ�����
"�dTQ�P�S� �'X�8�w�>(���=;���/��p�<����˗��_"�/�����:{�}X_[M?�]鳭30O,0�ڕmc�;C�xG�W���@��׮5 l2��w�h�Nu.g:`�r�atN չ�h���9��*1"��O*�A��y~sІQ��0B*��鍙���r�7Nc��n��B�K��d�fA1=�7Mpwt-SY㊠P���s�f�������9-x��Y�yr51�N!�cvy~3��?(u=�a`���t�h?� &<U@D�a2��i��g[�D�\����KO,�8
Ǵ9�Ьs
 )@!��zCQ$! e���
� ����Q`һL�	%��j
�0Tzgc�٬����%��(,b1��g��b͙�'�/:����+�f��s�~���΃a�9p���;�력$bf����JS���33( }����y�w�(��	@�c��`m�X^��p(�*n'���:2,P�@ȶI;D���P�k�y��M�#��7�ѱ�f���I;�Ec&�9`O��/���y�����Q��0d���	N�Ut��`������x��}fĶNu:�~uQ�L^΃2��8(˕�]k4���+՞�R|~ֆ��T'�=��&�4�zy����eT[C�LBO�fbf) �$��X6�G倈�\���E���n�}�;*E��'1�ρ�yO�OԧQ��Y��� �\�F4�i����X��)�;�u�v��sK?R0Ɛ�Հ5@�"ͥ�<��A����~�uϥ������1��$�P���S�k�Xx�A�XlwӾ�)�XjY���,~�1¿���ߐ��c��P�b`;������GG��,d ��܎I�A/mƧ�0Ռ1*�G�����zS�t�������N:餓O� :餓N:餓N:��](u]���#o� t(�`���/k`ݜOݲ� ;��*�h�p�b�iZ�&��U�R:1�s��|~�|����bq����'�d���X F<��8� ~v��CO�I=�(ec� �ܢ�_���#p��I*��
���$�|׌#����(���v`0�A�_�������0�a}A�s����w���K/
�w�s.R&юϘr�?�e�v���{j��)O r�$c^�iF���Q�5�ic��{O~���)�s:���/� .^ ������M��G�ޫ�W����uX\XL��{����eP_�J�F���F(�\��Lv����v?����,-/���!ܼu� ���S��{R{�~Νۂ�{��VS[���իT���sp�������f:�,��٥L1���ܼ9p���
&r���PpZ���8h��?X����ρ� ��V�+`��,�'�ne*r.�4��򓟄G{Ξ=K����Ǳ�v}n޼��m��	�W��P1�9b|��O��Φ3*�@M�q9���<�ꚲ^�Q炋
Q�苹�+���2?��j\>A�g��E�N�ęy@�!�i�&�2��7f�� /�F�e�A�K�+�XN)�}��"gs��#�@#L	<���H�TF	5�G��i
`��5G��/1%pK�O�ht�������{�3���k�5�\�@)�3�S\��@9�ĺhN�/�s�߷�5�� � ��W:��5|їP�S�����N��� �gJ���jC�)��L�m����JS��2��S>g+�Jt9,]Ԏq���ׇ��@�Bc.��-�\f$[��}������S�q�M�u9g���>��D�����"�=�|�!��YV��ʍ� ,p����!r�G����,�l,���HVBL*j��;赣�lB��#D����5sP#�hЅ��<��n�T��,h
�KĖ�ؿ���ٖ��s��kP�
�����G)�ᄝH��^XiH�+.Ձ�c�!
�g�u�GW���9X��̓�w�`����~h�th�a_�s9�_�5X8�d·jwk���F������u,�d�B+u�
 F���gt}X#��R��I�~���	���c%�.p�-�����4��i3�r݊�߈�!r�����=���y��UϨ:��^�Yҿ�hL��?Q�	*�9���8Ɉ��&�w>dۉ�,iϞLuMw�ͦX�~6�(ȎB��N:��'D� �N:餓N:餓N:y�I�>�cѼ\(����cZ�}c���J�椳N�]��t�
���]%�gx�������A����r�T�����g,:f��:���7�I"��٭�_��m��׽�3��ߴ>0��f�F( 'X���K�n�S�i�h5{��[����'5�9�j8<��x�pfk�ǐ>�3z�����`n޼o��Cx��X"g(y��C���L/W��e sȫ�����p��o�D��#ek*@���Spµ�נ�+X\^���uX][���=r�b��KͿ{w������[o�E��p8b�x:%'s������� ���-�C�G�p#�T����1`A6Ϝ�,//\������f���\���1������_�;w����2\8`������0��9c{�~O��ٞA����4�Qg*A8땣OHt\��"
�_S�Fb�靑2z&�P��F�8�0���Ѯi�U1k��~�a���|�l��g>���,c����f
��{	���a{{�XpRay���=x��W`���ܹs���q��M���
�	4���۬��g�A��掖рՏ,�\BA�o	\1�v��6�c�XІٝh�0P`J@��(5p��h��!lad� ʲ���l8�K�~��Z&6�J�=��B�u�� �|���dQ޻�2���%�`��[m�������.��U���Rb���w�ۂs>�����S��8�<��0����5��$I�h	�sk7~�z@vqq��}P�
�c&3���\{��x�L[�G�&�<�ϵD������������2�^uk>@²]�w�z������m��j�;�׍�-���P�����l3�t�-D�� �}�#A���;>.�}��4|�]���5(��yĬ���R2t#4�r,�1��~1 ��:��|ƍ=bT4��	+K���K�_KE�B ��� }��|T�
��7]��⾪ 
�O�'�+�Lb�8h)�A�2b�%@�/�&:�g�t
�*݀V�*��@�k���u=躍$��R,�OkV_F;��lu/W�~����ڟ�>�ؘϟjk;�S�3�OȓZ����צ �ME[���S[�`iE�v���oHL�X{y\�`
ယIZ󎏏�T�������Ӏ6��2�I]*��C׋��m-��SЧs�Y��xY��(�=Gk����݇���RrGK�:�v�~��S���O*�qq6�0���%�#�:餓N:���. ��N:餓N:餓N�u���ἡ������d$�8�<���v�&�.*2��y�F��#��.���d�e�,;��S����v���JP?;�J %�A���Vf�*`U>L�I�9�홸�v-��'�%�̨\/X��O��cp�ڍuz	��Ѡ1�L 3��A�)�ϟ� ?���K��ptt �n߁��NWVW)���� �-��z�x�&��S�#/�A����n��Ǻ`������SYr�|~�F�����^���~��O����|^�u�{�.P�9�`4���� �pv�\�~�3Ӛ�s���PK��<���9�5���G����kp<����Om���p!����ܸ~n߾	�?�$��݅�x��F���_��߼L ��8�L�u��v�'�	Vt�|nc!�g֯`��� ��I�⛮�)���s�WZ_�S0I](���8Ƕc��f�*��z��=�0\�x����/Q����.ܾs����8�cن��a���wwv`gw�t�hee��B����C.* Q���8��?.Nv� �:�:��jf%��WD}��ε�[AIQ�=icr� ��@.f_�5*��y3�[��)�G�f��/�m`��:�8�j�B_,��X*�K��=hE� '��l�� (˰g���T D뇂B�]ϢE^��Rl��Z�Z�m�\À1.1�k�k���&]{��.0�^���,�t�	�PN�H�S�\
@ۙG-p2���m���5q~,//�o����� �W^y%���a(Ϳ�r��/,e`6�Yb�M�)������o�=���6u4ȃ�F�̎58�u�������S��?�Ϣ��(���`!����N���[+%x/h��(����A�,��m���C ��lJA��3�C�ٮG֢:��-r���l�%>p��FE-"@)�Q��|ƾ:	�~��,��5֕%���[M;.C(��a$��6��KKI��O�Р��J��j�߳ȴ�:@%3ݱ��o��J2�Q�]�U�X�]H��n�<@����jfAr�Y,�62��L�����`kD�I+~��2r��N��ȕ���Y��൮蒼o,��ؾ�<cw�i;��Y����Qy�ϩ������>��E�׷a6s_ԕ�"O��0b�GTV

rk2�v-�]����Iq`�b�Z]쟠(oc�.�����Ȯ7Pv��,|�^Q@��v���N���~ш�a�P������a�!Q1��K�t�I'��DH �I'�t�I'�t�I'�N!o�+�<:�3��ˮE�oI �ۗ)���~�.
��D����l��6��}*DB���H���` �X:�����+����M���~��av�! j��]�?~B�@�W�2�b��q[A!�[rRI���Z Y���hjZ�z��*̼���������^O@�sa{�:Q���J�s���}�Gz?�S�r�p��mg�F�\4��A�i� >�u|����<� �_���1����>�̇����������W`o�6,--����t�]���:F���q1�R�t��i��:��sb���߇���c��$]w��� 8v|xãQ���,�t4ImS�/���ܹC�V�L9;3��l��A(�9��� *�a�h���8CV�6�sx��#Ф�j��`��p�������ŋp��y���H}�H�#fשO8c��htLY~�<����C�������[��K�	�	h��nߊ�O�p΄�۷}u�M�\,�P�]����� eJ[��:�%Qt�z4�6R62�`,�ɵ����?Y�B�����,!����u������5PE/�
�5^[$��g
b�涻
���i���@6���<z�Zy��f�A-�<^D���,��?۔2��˭-� �ҿ@��mO���fhpG������_Q����v欂�Y�Jv�ӂ��v�x˘~���%�8Nz�����PP�<��%���� ��~.���+������L��E�E\����U�u����r����#���*Pfc�E���sq��)�81
�T�9x���F��K ��)�	F��F�+��[���Ӣ���X�},pֺ�>�̪b��~*R���]i��Ko�ж�e ��x�i�����Y�c�3���~.��l�qD�VaKD�]�R�X�LZ򽑮cJ%;��V�O���\K�Ԯ)cT�A�mMßW��P0���_���=����=�f��~4��S�B��V~��Pb�u��ż����y���z@�~�5�OW�x���� !9!J9i� (�����+�7I����X��ا��q��#[�X�	T���
@���6� �b.��D�f��@�gW���A�~��-4W- $�=�y���M�gpi�q���>XC��O�(m?�~��Ҕ
i:8����N���X�:餓N:�1�. ��N:餓N:餓N�e�1� p��	���e�$]n�3�0+��2�ʎq\'{>%�<�4d<y\��k9�J�`�1m�u���a
��S'7�~H��2�O E����	e:���	�![�\�S�w�1�^�J@k�	��t� �4ק^7(��ϊ�6P7�o�U
tZ?�H4�(��F�1e�#�a��\ЃT�xm��G��!ӣc��}�J9�)���\�
�:���5Fs�S���M��L���ǎ��TI��/��fSx���'?@lx�ŋ�֭;��Ї�;w��9�&�?w����s}�A�ֹ��#9�S9g �8��5/�OI��kWa�`�akc��w�v�3xx��Bh*X[_�@�g��m��,������i�S��f�v�  ��y���>�|-��Yr���ufa:g§d2yF]YߢP{ᢥ`����9�{X9��?���g?�K��8P��z���D�CÙf+�}667`�����LϿGY��ྲ\��ű��F�c���f:�k��Wu��f �v�� �-e8�u���I:$�e��o$׬wm�Yڬ�g����x�K��y~�{�u�!�+����ZN$8�cN����%p���A2�Qwq�j�d,� �*^	��b����*7.p@�Q���
_{���D�b�����$�J�V�j�C�)��%��e[�����Ve�+�(gv� �b=)�\�!�8*�4.�1���\��-  '�� ����8D��@��	2�<�I0OX�>������X_*
z�r
����2o��c�b�����F����ɶ8 �ܒ�m-�EAx�AI�e ��<��T�#��&;'���@�dw�w����!44�}�!5D���Wpt�'�dЎ4Q�ّV 9(�Nm���g��CM�%@V���_'�/D����U5��1��cݗ�5��!m+�DZ�|U�F&;ޣ�v/����EQlR:��	�e�\�w�E,9^�G$ M����rL��O�u��s(��ӽl�Mi�Q>� �5pSm�ޙ�m����� t�+n(֝�R�WP��7 ���~�'�F��c�S���_��L&�^s�m����̮���}���� k�¦m8M���=t���CV��w@��=������AeL�rp9P%xf�(��Xih�3��P�C �(o�*b^������3�M��Zsʓ��Q��i�����"���?��r��Q�%*�-36�|O�A	���`�&��7�5��邏N:���M� �N:餓N:餓N:y
��U�^@-��B���e���8E�6f>�)71���L�%gh)���~_^�O��C)�
�I`��<*�B'K�@�J�d�3s�;�33wS��:�c�NkDBPP�?˽~���4����P�*�d�p�pr
�����c���63�#�������h�	�#�wv_z�ͽ�s��ao�}����?X"P�j:�ƣ���|�[����]P`�׫`��bٜù�Hȝ��o2>�Q��ByJ�L����dg}�~���\�x��0^�B�H_Q��lmn�Bjs�9��ܹ-8C3����h����� M5�0�sFԳtqV�gǺa����2��G>�Ӱ�ԣ�wv����_�W^�>ԫ�p��X^X��եԟ^z���=�,�0˿J}�#���莧�� �ǎ��f�����MR5��� Q2����u@�3פ�7띪#��2f��.�/�"��@ �7�$�ZX Pݧ���%@g6\���A�*f�N�ڣ1�{�o��|:{�,��( ��h8J}p�GC8:<�+o��}�Ω{=���=�4R�C3ӹ�N� ��դ+G�Og�&���X�������(m 2 ��)*��)c�����C��%z �Z0 ,���|]�1̆�)�ޖ�Ez$��51O�����C�eW��N(�����[�1 ᅚ9��Rq;�A)�H�eP��W
�X��,�E�;��>ɀ����v`0����m`%K���@s��}@'��덎tT�,/�8.İ�kI(���y>j��fԗ�f�~�k�g���^pH�cN�$�t8��7R�&ں�����)!���8?��cyi��_��*ˁ�II gu�Y?���#^�?鱘��J�e�M9˜�G3MsbD}��>H���0ݻ�����8gR{fXC	h<0�M�mx6��qf�����(E=�I�*f����>��*��Q#�d�X�䜜���Ѿ5�. �v���bO�:��8�	Y��i?8���6c�V�l�ӻp�����Ff0ZK�TRb!�?�q��H�o�d��e�)���Ud�癗a���6���K��j�W�z�>_Z\��G��zP��K�'�y'�a(���_8�K�O�s\��	��K�P�X�W��s{��^7*�5�ٹ����3����߁�}�4v��d$�G*������{_�kn���}un��L4G��ZV���Q	�(�>����{Q0A(&9�R4E��<��5P�VXO����~�^�����Vr����9f �|-���������ŎA����ы2ǰD֤1��N:餓N~r� 褓N:餓N:餓w�,�#)���)Ey��9+,��SQ�cO��-/7�����Vǩ�A �d-E�����فn���-g�F�WP4���-͑��8C����` ���Fw>�e�;�����3 ��(=эˣ �&�gҪeуQ���%����v�E}@ ��b�A�o�NG 4��"�F����k/7ٹ�v�@j�Ga��U����_���-������=� E��`� ����Q\s�\� �\_�_x��4̆�+[gH fG�@�R�WQ@�&��m�|vN;A�*'Y�.@��g\��U�nݼ	�k*9�>���:�A3��v�_ ����O>IW/��2�>gd��,�o��ZzN�0�z��(N�1�L�4HAO��8��.m��Q%Bz����O�
x,��,�LCj[��P�t6N�s^S&c ������ب�����{L%
l��ƞh�+i2<��LO��8I�:��������q�:5}�ߜ�ZA/�3~�KzQ��X� �P55��Gv�c�7Qj���޻{ ��g`em����ᑇ��3�E���3�S���O�������K$��0fT��'&����(�Iٛ���%8�#�#o5�Y�������?*�' ��U��n�.+	5:����u�FR�dp|1(b���Q�����@9Ş��&�)�s��>�	SƩ�.�A�:θ�R�;9�"� yҘ3��ni)mǢdP(��9S���I<��S�k\���	o%\
V8U�� 	ܱ�-�>rvv���B����X�]��@�j�݌:Ŕ�Zϙ� ��`���AY�c�pN8��g��#0�s�$3GGp��Հ��+^7h�v���q�� �ˬl�{6W7aeЇ'?�$<���`:�췞����0����H�m����E�˯�������_�{���`ss�^y���_M�KkE�]����Y�5�۵��1<f>�)5~Y70��;����z�����ʕ�w����e^����EfE��8p*0"(�i��"bO�@y=@�@������Q�L�+[�M���H�B�^�}�i^#��e��s���2K�E�_��&��+P�����ZRBK&(�=/�Ŭ`��~��Cζ�N�����0�[X���MN�;(�MY�qz%�VK�8�� ���lQ��͞�lG�ô>����]I�4�>�O��~D�TC��53�b�'��4�A\lk�����qI�JW�z��k��u(t�TD��(�Z�*(�ރ[�	���!��kAVz6�6^���v�=g��Ol�N/�?��+��l���#1x�E��.`�ao��d?,�*{5��9�&����g��l6��]�%�/�}�{�{YK|�GE��5�:���c@vǻ)����B�a�ҤP��&�-�`�^�͐15U ��E��q�@'�t�I'?)� t�I'�t�I'�t�ɻP���zyrIGuV�YS�-�g�/��P\���E]\ Q&�s�����,�i�v����d���Q�M�̟��u4�2v�q�<;	���Ao �9O�����Y������0C���Y�3��~�xY��U��=�s\#3����8�1�#�:R�c�Iu��~� ��N/&�1��2/766șM��ԝ��݁Ã)��K Vp%���Q�zX^]�͍3p�{੟z�������N�W�P���}0�((�3��=nݼ�f�J�� ���u��J��AKFbY@��C���c���ǰ� Z�ݕ��|/����R��ZjN�3P
f0�=����w�W����~u�� ����V�0t�`�u�6�}��A����ԽR������=�^��i�q�դ��Ȱ�����0�����z�of�c{Y/� �:23 ����]���L�-��������������x��$wU�� jl�]�c�`��H%�("ћs8AcӤ�=wn�E9�����w�>-���&�c=��� ��DB]�Z[g����2ܾs;���I/Mj,�@��Y�S�S@H�&����fC`�9��͜�_�+ӱ�g?�ڲ���P�f��$����t�b����p��Z���6~i��V5�bx��b��cS���p2J�QpO%�J�����p'�/=e<C�V�D|�Ѱӽ��	T��,���b�>�p�1���Eh�>s�����S�1 +������8�sb:����Z� � �
]�+���h�뤫 5��~t�c�P@K�r �6Ѭ\+��!�G<gii��>���V�V������}�5��?�3�����ko�$��>�^�\߀���Ʒ��?�/����4� Wwn�����t�|�S��?�g������VU���?�;wv���o�*-]p�`J�hc�����OE����9�Qz���?��Q�(�;�<�r3�}���)���V�f�6�3��f�vяO]���)��ϣy�K��Nl�"���!4�mZk��,�雴2=���eNm��v�Ab���4
�C��7��@ԗ �H�[���#X H���7'��@f��}�2b��Ιq=*�s��)L���,k�+�e#�n"ٹ���! �ȕ>���K?�\ ���\3p��K޶���K:�+�mJã}��.��N�y�b� S�+�Hp5ϸU��r9A�����h�S��&�[������.���As�\�m���+]����+���oiߋ�S~Ol#*�(�k��\���$�9k8��Q�_�'���?x�m�=��}��=Q���� �/�Iɞ�w:�9�?��_?�8�"l΂v8�����R�:餓N:�ɐ. ��N:餓N:餓Nޅ�X�2�Xs�]�Z`9���ݐ��'�p��q�>���a���Ӌ(A6��B7��;q�:㜝�r�9�+v֜i�κޠ�G�F�N�A�E���'?H <f���e����k�|<��s�^�HY�O� ��g����9X��;iL���A����	����ǰ��uo  �dE�c����������܅�dDm\ZZf���ް��*l嫫sZ�j�+���a�Cz=��t�58{�<��௾�-���U�p�"��~����}��������o5e`e
`�?�S���AqrDgђ���I\�^j�4"S�#����9����% ���
x|1�A�^�G��3*��ZXZb�80x�]
�XZ1�T	�=�����Ʉ��%O��P���׿����>���)����V����;w`kcz�NG�$����.����~�����	�`V ��{�Y�X#��N9�wi<�^�9��QT�"��ڋ�q��t̾����C W��'؏^ηz��ݧa��\�F��7��O��O�#��nl�^�o,���ٿ����O�U��7��6���7��,,��s��W>���0�}�1�������ԏS�3w*� ���B��؟\�� �.H J66�mCx�⼘��$x ȹzDh�Aԗ��ktf%5��I��gl/�ᮄ dpϫ��:�zO`��df�#h���;=���"�mfOVZ�D�k��%xB�n�M���9�����5�0��e]�u�Weˠz��+k8��F��ʋ�7=���x��-A|�23@u�:`Е�#�:pr��C�Qo<�������L�Ҁ ?��h�z�ǹ��?p���O�MZS���OQ �mI����3�����_�;PSp���{.�s6�7���p��eػ�g���௾�u��/}	�����}^|����w����*<�SHk�%�ݻ��)7��jNn�ԡ}L�_P�4`���#����\�td+(��zd^��گ�#�m#0��?��cY��E@�0��ɨ�{���&	�
�4ݘ���)(C����������s#u�,��w� 2�i4��
|ʞ$��ro&D�q?�0#�������i:�O�]���Jwc��\�WU�]��Z���Di�$�u-�N�3;��!���U&���3���T��� ��g�a���̤�|F��>��L�9�av��
�k R�1�3��y�K�%3T)L�[��=L?r)g�����-�nq��zq��D���<��R��̦�A��1>��bb�7p٤)�ab�T�i�&S�����<��a%�Q ��؟N�=X�Ȗ�J�� ���
ڳc 	ڃi����SƐgC��,\�@Q�r=J�w^�2�YD�o��D��8��b'�t�I'?�� t�I'�t�I'�t�ɻR8S�������u�A���Xّ�v����K:��S>��+�U��N��ԑ9nԧȈ�4���~�}�uŎY��!WpU���|�?�<�ȿ�_�̚	�)�:�x�=��~�뙧�MfLc;�`�Ύd�10�� �>f I�s_�bF���I�`�GcT�v�8Ak��)�ymm�77$�~Z�<��q���88<$G��`�F��Ԟ�zI*a!$�����8��֭[��0`0���ғ��t2�~B:a������� i�9��3*o,?�������ܺqF�1����������ߘ��>g:g��=@n^<TP ����)��2��F羇!f�K&.p|�S?�}�{�)���>�{��}�|�k_��tɧ�~��nQV���!9}����7�"��� =�˹�ЧTCo��M���)L�c��ݥq'�=��g����;w���o���>Q�#���{��0����n�b}����o��o���0�N�Ѽ��������X]�A�Y)"��%�%솦0�JM�6�g� 3�	���	ſE�Nbs��[��`��[7�=ˋ+BYAi�i�s	��R�$ 3�I�_����2<��p>�[�L鐞�4 �3J��>�GGt�^|	�x��t�)ܸq�ܾ���w`/���ٲ��Jԅ~�=-%�-6A Ĺ3�7�$�*P�`ꓚ.3I
1��b&e 2[	�f鉭a�A�d�pQ�DQ�TV
r�A�)̀�R+�l0C`��tL�x��'�S��$hw�5l��>+�!���98m��s�����\��JY�^~�` �Lu�5�Y��tjϯ)�=*���@n#�Sh���a4���'�@�ٝ�|�t�����Ɛ��_,����'�����ʹVl_�
���1�H
�:�AH�������5X^Z�o~��iN|��o�C
|ھ�Mz���B�F��'�ן�����o�fZ����W�:�D�0��ee4�������[��v,# ���e��r����M��u��K�G��8
|�BI�
�xgeW�FA�Gj�XPx�#��Z']��+6�Qѽ�յ�g��}}���iW+l�F��nQ�X�`=Tg4����vf��/��@�Mʏ8�w�g�_�Dv]��sl݈����,d�Ǹ������<IFt%T�N,���^7�p �%A%��I�'�����Nf�p�10���1 ��c�O{��3+��H����:)E�13[�P�:����А�v��YG���R�[)�S��>���+�")��-��8�v3H L8y���	ԆA��r}�8-���^�/ ��tV5� P����(��0�2�a��Ĕ&\Z���zHA|��"�,� �Q��m<a�d�"�Bt�>��0j�����3��u����є�W!SWC�QS�Zv(Ρ�|K]��*Qh��rP��줓N:��'I� �N:餓N:餓N:y
Ӎ���"7U�G����l;�T�C��p
T��0��k�X����9���7W�@�EK�"T�Avdfz����*��o\��7~㿀�{̀A3VVW�ejwv �3��ԟ���e�c�vM���g�"FP����\���#���2zVi/��B*Py�ޭ�Z2D�K��C@���:�M�f=�"S�� ���3����0N?�� Ȍ���и0;Bv�gV�1q0���y��Y�0syy	�)S�r�k��ۍ��ԺvP8U鹙�Ǥ?X����>x򩧨N+���t��^�l_�J O�e�bY�����4ղf��A�Ne���A��2ّ�`��Ğ���P^�����D�z��c�?F}:�����u�|������ӟ�Ex�8c:&�ׯ~����/�IjC,�0kp�R �#T� =��/����*1`�Z���?o�y��^x�%8H�K U�4��K}����E�v\���gϝ���
P����z�/f�{�u� �  ϭi3��� �@�q���i� ������YYk�i�c0)�8{��Q���{|��l3�|C�|��Gy|B#|�¦��y��sS��.�`ey�tK&�y��S��4?�kf�8�uB��x4���n��� ��p�ڏ�-_��Wy`_nB�ʲm3W -'��ٹ�*^�/C����gS�N)��5�5���)���	�� ��5��0(�lϽ�?���WFg\ �i�ϩ�8�+p����lN�A3��mw��K栯��ݣ8</	.	��@��}���t\w� ��\1�ǂ[z-g0DA`��� �S%M=AqA��}�׽�2%�ʔ��ﳭW:��`1��X__O?kp��d���gKp��X[]�������{w��l����Ƈ��d��+߇+W߆Ǟx����x�l��o���O<N ���1���k�hZ+���� �9H����ൿ����g����i^���{��OV��0N�ŵ���#��Ki8%�J���A�No(�ݴ&�t��_��g P�(D�'��oj����@��(����b�(�|,7�g�zQ,���9�c�y�1ڞ��USq�I�/	��B}ol=z������b�%�	�L�lL$�������x>��${Yu����^�A�,ўQt���L1����$� �~����	�QSQ���(考�<yf�![��!.�upa1�s�].%�O,3a��	B��lne�����5�:�y�8���~k�}s��|����F^���h`���xJǗk��u?���s'�y+,}O��e{˥�r�|w:O%h!j@	m� ��3�s����M\_h��Z^E�>\���6�"�E
4�$��/�$���ɳ*��8�l������ <��C��}2���� ���_�o�[0�q_b����8E�TE�gk��*Fݫ;�ۘ��>�ljt�I'�t�"] @'�t�I'�t�I'��k��J�T�v��v�^j�b�e׋(lr�hQz��>;	̓ܒ6(v~+K�o�����\��pXm�� NLʣf8{��ɔ�Xc�̙-x���O ��$��J]3���ָ�+(�����H�O���@w�i�W�W� ����J`O�\$R(^3���6���>�D�]U�}z����&|�\y!��駞�����+`]A@�hV�	� z��k��q�ܯx�	0�����b��CmqH�_��ԫ��K�c�2Ps� ��b��ot�cK��e��g�LD����T�^�#���x��;���������1��jTk,��Y�dd (8�b�K@�ا�����%�^�I���`	�W����߇>�8�<ll�SƵ�m������=��O �ݻ���q6�棰��7o�L�z^y�e�Z�1o����gv��hL�M���|�GzU\��I� U��ؖɏ��',��lE��!L*S�{��2L&������h�M�e�R}Z)�������~9�����ev�c�Q��s��Ϥ��P��b<���b����qp.{�w���QJL�5!����
�[���}��P9Ϛ"(�Fw��2_ind��9��oVb+���ՙ_�{%&��K��� �C����T:��o~�д�(D��Q|5f[��W�� '�-��T����f��V�К��������
��)����M���AkPA��t�� �xT���ﭾ(E�,�W�vf:p<��弳1�`��z8مK|����K�A��|�3p��9�WVV�- �xn40O��}x�����m�:{��#X�{
 ���y�����d�q>b��h4�s�Y^�R{.��������{�e�̭����O6�b���K/S0# @��W_�����
�'�\S�I#��7�� c�(�#����6�Si�L����d�������p) �leMv��}����A@�<�/�J�x����(�5��*{�5�L$:�\1���<�eWZ%�
e+�y��� 5#
D*����b�N,�S9������x�Lq�¬���Z<O���{:(n�SEl��]�уt�K"*�\�B
3ʗ�kV9��]�We&��L�`NJlEa

��Ӱ}�}�wڃř ��w����^�G�k�Y�}1��(�m/?�N�K#RF��y<��,a�C�hʷ*ƪ�A,�t�v0�s�����������K��x=�ڃ�d�Gq�~�֋��r��y_�%k0���*�!HP��d�����;:n9����{9�)߂{ۅ�Ux��G����i_y��g�h�����=����x�!�
Ş�ư����d�z&v���ȧ>�U֒N:餓N~� 褓N:餓N:餓w��|�Oh���{�N^��^g�� ��K<��������&�rLj[O9v�z�,2�[����L�k�CK��b� @��>���(E�(�	8�\K����3�)�Ɣ�n��������4����R];�P¾l����G�nh�
Pj�	P�u�	�'gt p��g��FUƺ�L[� zf��+��V�3�@�L& DԜ���RF 6B=��1�XYY��(���z��l�����O����W\����>�g�z�'^~�а��V��3ı��o��l ��G�_X�n�'�b��*P�cE��
E��?<�5�+pmy���^].]�iU���4��h��/��	L�|�`qi	�~����+W����{�ç���=��Nχ��䰸��o�P�c����0!r��R�A�! �9�+��E ���4���.��/u�9�}t8CE) H�d��d�3,y1a� �E�YwT1 �&x�/�ĸ}�6���e=$�a-�!��3C�_�Dґ��Gp��n޸Mz��ȓ�2����vv����>1P`a@16x��Y�
��3i���nc(LҗA1e��PrB"@+�N��� �}e���b��3�Z��A�	�,@:S�6�^3Z ��Gєh����Z]A��Q�D1b���"�l�<����l_��6
�E�(?O�Lb����q^���Р���s��������vO^�|~nЬJ<Ӎ���b��*��������5�=`iy}�1f,Du��l��?A�BA_b�Z���z�_����$[9���5�e����G?Fvgfp}���7��`[~���*q��y�R;vwvi�KA�oHc�����Ԛև/}�/�?1�~d�9Ls�Y-!����y�
~�?ɢ�C,h#��n߼
o��<l^�7ݼKg���X�kR�NL���`@.mB�E��7�s� ���q����ʾ�s0 >�ÿ�T�	�n�� �ӂ\k0�bK���D�G�9p�5���uC7jc�������떝)�g ���(�@C�r���	����J����b�{$4f��o����s�a��В&4�v]J 8^�9�P�;�t���g=b*��?�Ԧ ��,��8M�5\OP���}ػ�6l����~��#b^
�����`�Hw��9��0�9�ˎ�6Nl׌9C혦�� F_|nc�י����r&�O�r�BO�|]���rʩ��r�3�n�� �+<g��p��S& ����y����;R�C�znŉ�<�f�3:�K*؅r�@�u��WCA��dt��Yxᥗ�^�a8�y�Gi_%�Z����џ��V��=��TO.u���B���O�]V���餓N:���D� �N:餓N:餓N:y
��v��1ڀ��5u��p��?1�R8�N8��k�"�C�]H��}�4C�,`�Qsu5��Pf�勲C-�-L����8ƽ8���(f��zʮ|�	�uZN@��=��0����y#�}/�FN��8�'j&���T�>�+�+�µɯfR�۞[�t�PR]��]�/��T}y
 E�ű�\E�����u�Eg�ǀ�d��*�@8
4�� ����3=t"���%��sЃf%���{� j�Z~b��v\v�0�	�>��s�dv�R���{#Y����q@�W�ڬ���~��	��M�D�~���4��q� b�݊���B����S����C��ڰk�]zE5�н��lmm��k��~��8���t_,�����)�gum����&��KA.R�Ý�۔�#��g�7������:2=�l`4�P�}�@P��P 铃��x�D�l�b<��l��޽
~���S����$ ��35��PJc�`�^
���4�q��a��Ω�w���|4䢧2 aJu˱�>2 �������M�C�cS�~!zu�R�W9P���;e9[�Tp�e�.�>
h�H}��>���jnuvW�Q�拍����,xn������A�~���8d۪+���YRB;g�:�V0�K���aKT��W۞�)��R�����TF:U�+=~	v	�dzq�>�S�%��q��t����m�m����U�.�=�Q�`x<����4�i��:�sI��dK%�R 7�S�W�=b�0�bԛ[®����4�����0͟����6���g\��_�ʹ�3g6a<���ptx�lɔ�n,j���E�z�:��ai}1��Bx��-8>�v�`��^�ޔY(2Bfz
e+pEI��Ȧ�e��d:�1_�g�}:���w��X
 x�Z��4QD�b��(yx2m;O�&����(�C
62Y�U����h�UU���VZ�����A�������4C� ��d�K?��T�YA1kݬ��ب���]�%��׾�fB�{޷���P��%�X���[�+m�i�r%S�*��y�TѺ��B{��N8�;i��L����*̨�p/�A�ȉ�wSb�@ ���R����X0mdf,��eG�-Pr���c:��^���^�:>���EP������]��쒬9�m.�/��	�P�wb��l�)XFS�9x��~���^��p-]�A\���GP�J�7���5=�~-�D���5Q���o��;��A�����.<������m8Lv���ߤ�c�=�m�ߢ}��G�Q��.�D��؜�&F�l��qt&��;��ة�t�I'���K �I'�t�I'�t�I'�J��%�h�G�y1��p֚׷�r�b�s��G;_�y����d>˟��� �z�����ob��Wd*���(����T����AT�����(ۜ���]�����J�&�)�=,��\q�s�mdc�f��s������NDv�k�(�,�cE5��q��(5�%��ў�N2�9�T��KD�t�@����"M���}#h@��x�A�T̚'jU�k%�����lo�{xf�!pf<H� P�<:ԙ�I�gX;�lZ` (;h=TX��\�7�ӌ~�I?�ZV'3`)A�G�Yv�S�ɜ��f���|f���nD;���8��V��(���L�\~ J)�m��{�����k��p��=D�0�Û�l�JWZ鞔k �B6
��tFu��n_�/�����[W�)�`h��8�R2���\
����sZ�;5Á�!u:����{�I��:��v}�cx����>++��3S,.-Iٵ3.C@�%0�Y�W	`D t<�p<$Ь��������,d	PY\Z$��4�2 �q�+�nY�}2�R���y���������0P�0[D��@ �jl5�8��%ZR@|+�K�42� "~�f��v/m)i�v*�(�h}������0g��;��fA��������y���$�T��|`�ȴ�,���a\�ζ(ޣ�׺���!e�j[���ǌYE��U��m-C�2��ک��=�]U��)Ƞ�0\G��"(�O�2�<8���i�������g�Uc�h�@����e�!,�r4<@ko��6���S�����XB�8I�������nݾΟ�_��^}���׾
���_'���+�ᩧ����8<�%�|���e�h�0�:K��2�q��n����~����m�����M(�ɛNV4�AX[�ƿ@��� �+�L�LY�M�	�^�4|���tZzR���g�
��.c�բ�����|8�`�S�+�y�Rఔ ?-5�	��2E
���`�yZF�����3Z��=�kו׽n/�B�
T�%�M)g�v��*	�s��Ќ:+��2>6�X�'����;�|º������RHT"�m�	����4�jd��xP�(y����5HI˄Z�mH��,���1EO[�lOTWs`�ɾ/��,�S�ʹ[�@y����9���pRt-��((��1SI�YE{톂����=OC�^�/
�th�:��̪��m��Y0.�Y��X�y�FY/��V��o@e����RV1�g�<���+�����LǇ��G隁�ͻ�/�s�֟�^.VΑ�w�>�K ��+�&N��N:餓N~L� 褓N:餓N:餓w��U�i����F0��Tk�T�'�/^f� J��L�L��r��ke� �w�AT��G��ǲ��9��9@U��8wpvR�s�S�{%Խ3����*�;w����`0�sg6�'�q�DM>������;������W�#�iq�D S�@�Wq���c�
���w���d����������zLU� ��F����&#�7��\c}c�������J)n��X�MFS���Ux��{a2���)�'T"���J_��GGGIׂd��Rx�Z�*C�dg(:��~�5�^#�Re'��?U+)r�c'��^�3�|�����!���z�?�:�+ʖu>Ӷ���Lv���k�*�j���:�_l����b���t�xF �(�?,���8�׬�p0c׳�xx4�A��E��Qp	���'���9������G,..�X��Q_p�˫���3�#�D�B3� ��Ց�W �Lǝ��r�����:��+�О��.-`ym�I�p��^uj�p2��T�ّ3)�ψ���i:?=���
��/�k�9�ɔh���S�^�,�G��&6�g��<���W���b�H�Jm�E�$_�8�QF��
���\��Ԓtw&�A��h0��3P<C�9���1�=��b��cҀRk;�XLm����9e&�P���AD8f.ӕT�}Z��祝@s\�3 c�`���@4�Z:k~�P�a�t�1X!�IX(����@�CJvH����"M3лl�\0��*�o}�c/����I�h����%(��Z%�l��@7��[ ��^������8z�����誘ڟ�L��AC��̦0>>�
סل��t���7a8�P��������\��ww�a}}n����5X^YJ�����vvw�����C*�O����/����o݁'��ll\J�?�������������uÐ��5�^�H� ��
8ɬ��l�'7!k�k�,���shN�t(���`��a��-`�i\�B��}g]+�KUUg �82�^���u��+b8�మ��h5A%0��Jy�(��W��h{O��}5'ڌ�7sQ�~l�C,�;Z;����� ?�j�}��h=T�^h�]��
	�UJ �W3���z����͙�4�$�E)�=�'��_��0F��� ��G�]��H��j����4�ΕeR��4��(׬�E�gz+'�y~a��Ay��{�z�����N�H�*��� �F�����a��Ï>��Gi���B��@�����nf���>G�@
ܔס�[e�OJB�R�t=*���z�� uu�q
_V���������G~:J�|��Yf�<���h�Z���XE��I�z�mb;�l7���)(���~6�^97k�.0z8�*w�I'�t�c,] @'�t�I'�t�I'��+�" M}T�eG�:�%sY\DѲ�4����3�%Z>;���^�Yy@���:q������`cu��m�:;/]�<e6����x�t��G����'����3[[���N�6fS�Q&4_��@�s�}p��x�Ї�3�WҊ �[it�������M�Ɍ 4+_{�5�&�	��ؙ�t����l�6�F�����
Հ�F�!e�c6g/���k_E�:�(z���r�ꂂ%X��GGǰ���}j���]ٗ��PU�&����T��Q@�E~� [(�ب8�]�2;kG����]ƓJ8�}nS#�J�d:�;P�^:���i��t������Y�YcJяL�:��gjVaH�|<�#zxp �|�[߀�W_%j�T[H����7o�d�<��q��i��~G3f����` h����Q����6��A�@�c�`�==������Yv�����e�3u�;+���`�0����{���mu����z�����A��F��!��\�q0,,,Q�,o��!6�иO����l_���;��̂5�1P%�8�����3�ds�`*L�\�
gϞ�I�0�������=
K���vh��\�s9����<7N��F���d��G?�S����m}���3�A����~5�A��E!��t] H��և.ZҺ����ء�A�J�{"��g%L�Nh�Ӷ��г�4�U<������vV�z�� ���y�Y��P�k@\T��=z
IB1G��� [g9ի��y	8���nS�#V���(ɡ� � e#v-}sttH����&�^�7nP�W?�E��G�1NkR�߽�OA6�R_���bـ���}�s��F�1��ޅ�{/��;���"���Q����|������W`���t�1�Af�	98#
8�0۔X�˶H��g&]�ؤ�4&26�z΁!�4���*�s**��l�d�K�� H��������
Y���;sV�rP��`�SM1O�~��h9WX���@_*�O���s��s����ȴ��t��9�F�Ǩ/3e�+/"/luVpY�G�Ă�J�Z��RUњ"c�C�w�{4��#
���ܢ�z?��lc-J�+���K�����].��ԉ���K���f�%�9����x	�l�c B�������7��i ����BJ޺���.�^�	�N���3
�Y^[�z�@6o��M3
�<a�~0p���>�����\�&s���nz����h��)����U�y�)yH7�f��%� e�0�T�\4F�[�q��x?�%�XQ�)r�}/c����۪Sd�(���K'�t�I'?� t�I'�t�I'�t�ɻP�J�d��	MF�P�I��`�`�͉�r���E�;@c��;����}��7�� ���d`�8A�5N|�X<n�~a:Te�<�������I4���^]{<g�{_ =�%����>9fOb�?e��=Ѥ��" F�^�ͅ@�����x����H�ĺ���jq*
�I��u���VFg����~x��G`}}��	SmGM8c��#���*
H�qt�Azu|0P������.h)��`p�M�r9;v�F��Zf��D�inm�K��Y\�����h�F;?'U�ը�NGt/��gv��ا*��
0��K+`���f���RYTG��5S
�@:[����6�.R0�����O=����J�t�8s�����1\�~���`gg�ɑ�s�V,./à?���,Y��2���/%�]w����p�VjK?Ξ��s���`���D��6N�mk�Un�o�p�s�z��3�ǝ��G�}�M���}�h���rp ����0��\�6�@��SI��`0��(��ϝ�}ui��^�M}2�Rv �wppD��X��B���4i��b��ln@Hs�Z`p�b:/���&����l�7M�й�6���L�"h�@�x������ux2c��fj�"J�7��2�m#�[���s�0�d�s�H ��.f�(슘�<��S���e9G-�lnF��<9�R�-f�0_�֛���l9�"�9���a�L�	,��d����UV�܁� ��4 , bѱ��?<�N;�A�J��r��E�k�]�'&��TZd�t�kd��χ�c�w5�Z��A��m�������(��"|�ߣ���=��{�/�ٗ���[��sߡ��^������{�3l�=+K��������?���n�������k�h;i�p���$��m��}�l_�m����x�:�s� R�+��at�qyo��e-P��<F.$!d�/���z�b�d�<ʘ�ݺvy���*�6'�� ��%�u�pr�0�ꀨXf��C�ז/B���c���p�H7@u[n���ztY��9����`n����˶H; �o������P/�ۘ�W ��sB�˶Pڪl2�P9��*!�?���/�-�3�5��<E�p0�6;�&�r,��� a�@q1ע�	Xw��E�窟TrD�P9�Y��6fm/�(l��vIw���i��7��'S��J"p��`bJJ{��g�����g�}���P��E���ω� ���lP�r()�,Ip0c�L�˕����]uH�<��;eyi8[_#=q�W�מ	���c�� �X��槡�|9Hʇ$���T�֩�t�I'���K �I'�t�I'�t�I'�J���U���;(�L�Y���)��������\.�vl�N8]N�s
��g(�t�󴥭&ǁ p-/��������=Rkv�z�5�2t g�e��Q=���訫$Kޜ������@�B݃�3<U����{@k�]������*��juP�A��-���H�F��Y0#d�ò�XXX����#a0��B���j�A�]��U�]]�z����;�}��Jk�Z%�#U׫����}��߷�=���=�tD�7.D�ʛ:�=�G�D�8 ǯ��ڃ�A��7	(�:�3�R}�Nk�4l/EqSTTM �6���_�x��5~�QXٳ��k���:u
��{]�э���z��ol�[�v#P�#�Z�q����T��UB�.J��3����������n$-`$+��E yaaD�bʩ��qc�	�ly�9�t&�^ߍ ~���1��N/./��C�\������W$s`T�uǯ�� ��:i޽Hj
M���'S��>E�.4}}���ԇ�Ͽ@�9F��xb?�=P�W����Ӧ�[[���SM�h�&s�s��LB�*�|�(�n�ps��� �e\l�E{�}%d
v�y(M@Q�o��N���:lo)jKC�����h~l�q���,�;�=ʍ�s����_�\3���\@d
�����i,P- �����\s��!".��D`+0�6�H�7�#�
$_|��bo��q`&�C%�A"3��*��wCV�*��3"�R�3�	*�ТD�  �S���t���+�@M�o�k�jP �,�������+�Wx�'
Gg�{��K��8��Yl� �g��7(H��  D�օ������^R$��w,�b�~\��O��#�+8�R���s=(v	EW���,-���s��ߔ�fE R"�rl
�ݱ�����ׯ���&���F�����ߤ=	N[�c� �-�j�Ǚb�>��<y��g��\ں�2���Z�c)Oe��	�	 Z����6��]^(sB� �I{�Xl��S���YI�S�'ɑt����Zz��|��HZg��eg!��z�j̓x����۵���Z+ {>@v�%X�Z�����[ڥq�v|T�d��;��:R[˳��kp�;�q6ߴV�������#�a�g���f�,#�2�h!�ņ�>�s�7zt�0�� �&�w�V�ރ�%<�DJE�����5��'�%�4�������\#����V$3`�02b��2��񌛔ܤ��^�h�� fD�j���^�Z�:���B�մ^�P���p�Cۻ�Q���3�TAJx�7{�6^��c�s*�� ���SA�-�@�ȴi���l����3ك��5����S��gH!�%U���˩���*j�(���6��K��-�ZH9;U&�����x��5��H�;�VW�ҕ�t嫡t��t�+]�JW�ҕ�t�,�~��<;y�8�krҪ_�|�sN����%2�\�����e�y���w�Cs����n�̕/�J��ú����(8C��g�F��}���Y���	���9V=@�r~���p�{=s�aoO�>}��`aҁ#�ׯl���E׿��޿INGN�缱=rV�����Y޹p$h0�� ��ԈV󩊇��Q��[8��H�`���%���н��յ���^5 gkUm�h8$i4\�7�m�0HDjA��(`T&�JǢ���X����s��q��e��Ƈ�Q�C�������'��#�wH�=kT���bv,�s0=�* (���شu��/�p4���{�$�MM��5l���tƤ��G�&�����Y�(k?7uI��/��p]�\���^S�I��Z	���a���8��L���[[(^@c�چ<$p��-ECJ�E���a�u��9[@��L)6�Z�]��G�!� ���sdf`�Ăk�^(�A̆*X�#E-�\�ӄ@D�u���(���'H�T5$��J�s�y.�k���y���d+0bzc}�V��6ya#T(x�`o��a�7�q���PV®1`D~���&��m"���0�@� ��vm��@b)cH^j�,lM�����I�@�Q�XT�͝ s�rǞ�%�{f�e��  
�L��t��] R��ʤ�3�x��#!$Hd}�(\� ��l<$��� j��ҙ:Gu��/`f(ԽLyh���f�.(]��O����d���6\Z�W����3'�/|�z�)R	oo ��H �/�X"����lOB�Cc�I�Q�f�뻆JCr��Nkb�6ﲐ겨��"��(�|��b	*���.��>�5�[�
s�6�w���r���F�~�:��t��$�ښR�u� [є W�
�j���'��2{U���w^���wɡ�e]xy~����F����ީ��V2�/jB6	�Y�-��d�@�����x_Z���B���Z��ƠM>�`��
���n�0{�E@Ҁ�m��*��G🕪+/d�N�)
!��<&`VB�P`<ʳ"�������o�G�4��9݋DRL���K��ݸH�z��N@%��V H-y�m��=Bg`��[gN����A�k���aR���t/�bM�<�F�3QN�<��$ ~�g�����2�<�{��&�h���#�(�Ɗǩy8���X5�I���Nۺ���py��%�,���xr�'|.�r6��zs��6Ҍ	U����.��@퍕]�'GRh�get�+]�JW�jJG �JW�ҕ�t�+]�JW�բ��y�ɥ������r���(�[���̑������w�G����N#��_��� ����-�l�X}��IrW��-�z����'�����p�=w���Gr|�L�51�9�܂g�>	�/\���-x�Kn����k�ǎ�@��	�2�`^q�(R����U��ׯLT��@E	��9�B�lq���O�USt>�蜬�z�C��K��b $����C�O���?7%��Zٳ�+��oy��ɀ�H�	��\���D�I �ɼZY^���EJ�����"+^���A�A�Zt i0�z�9��� N�}�M�4����<f���ӌ�=���{ii�@Q��(J��P���8����c�����	�*Ν?��?}�{��C�,�8f��F��d�v�=�(W7�=�4_ЉK2�"={������a8�haD�����?�����Gmoo�8a׸��u?�\��N�>��������`Q�е�� �˺j��Cx��B���^�
*A�0�(L��u�wu��&�?��H����\����@kMZc�"� 	D��L(Q ���ۍт�[��}�$=�6�"��T4�;�=���{��٭{i ;n*	V�P�P���eNA��S?����]$�/`�ʞ=��x;b�����\��c��f��� ���W��{�/[�}lA�+P��ULr_Ad���H�|$~!&�8rB�����N�!�E�۵�ͿۧR�h�h�P�*0���8��8������;�^��������Qڇ�~L݂cK�^cϑ$�{F���|2�S���y���<�@�<����T3�WI��] ��e��0�jS��96�l=*0I�P���>�$߃N\�sA6iyޮ����|��V0<��f�aْ��+���kZ?���|�����?.rQ�!��d�9�m���n5U�W 7W�0�+�����g{C.�����j���L)����n��	�l*mkM%�:B�hvGN}mT��W��RP5��@�1
�v�JM��+2�ؖ�Ƽ<���?G"�ږ( 3^t�7«^�j���`�,\�����	�}�Q��G>��)��=  ��T���קE��y����7�����欳Bi��<K�5�˫��O<	���g��3'�-U��!�B)��_�zx���
�Ν�O}����SOɞQ1���즃��g�lv'A6A�)"�z�sZ�ub���+)EԂ ���Y��x-g�\���)S��@~7b��$gޙ�!�t�� ��^��.n�qJ]�J+�����f�V��E�:��P.A�'�e�� ���mF��dX��t�+]��WU� ]�JW�ҕ�t�+]�ʵX�O��:�T:[�B��K�����bѓ��Z���A�?�x3��弶ιl�8p����?�Rm��v�H]3�r+O���(�\װ~�
����}�=�ַ�n��f��|��]z��}�G��~��a:e��Oz�O?��š�N5�w���M����<�.��`p���۠ �T+< đ@�H���ok<�զ�
���.�ҁ���5=|fi��Ć:��DY����;�E�{ޱ�$�KH���(-���x��KKDP����Һ�H\�td;�Y���/�#�Ύ�(�;z�? �x�+a�7�$ ��ϫ(ªD$3����x?FEaollQ0uC��u���	��Y\��,R�& y����G�	��v�4��z����
:t�9Dc9n���}{Iɀ+�T8;��'���>��O���g��|��lfc��ͱ2�z�.� 
�fǒ��U��%��E� LA0pJ���y�q"#��n4"7H��މac��	 ����I�^���,� �W�	;�IyV���Iف�u!���m���W ��\��+ɜ�
�{������[����Wyt"�$ �%�&����H�GT��`,{2�fH�خ1y*��~�d9�8�H�&���U����[��ԡ�I���~���ĳ��KK� o�Y"�g�ў={$��|�s�b'��1�ߢ��e���<̏��WQ{�D'�B��)�F�����3�`��I'0��l���e�kX[]�y��0bKy����1݌�0�f������() (X��b���m�!KD��w]��ޠ
1VY�vFi�/!D�0��$�3�"�]Q�p}����c�C���p�r�>������[�r�~�f�s�����@���l7����[k���`u��N-0��{�Y�.���=p�+���Լ��Ε�R@i|�|uC{=맱��p�@G�5����]�:=J@�1�;�� �x�m.�ݺ�.�*�rR�y�m̕tWH.�H��������5�ݷ���w�k_{�s%�cm�<'���{�{�����~�����p��?$%�I�90Ҽߧw���?����Q�5��P/6uXij����)�/��{໾�;��������ϝ�4�6�!�6����;�λ�l�ᦛo�|�}d�8J=��`D�bߔ��F�~'��Y�&��`C��� �'���==R�SEޗ�b��(
�4!٭��̊�K$M��HRTO��/�0�.%�������ݲ��d�S[�uPྠ߅h�K��_r2�b]g�t�+]��WE� ]�JW�ҕ�t�+]��5X*``���X@2�k��@���W~,uΙ��ʭ�
s��P��؃7- g�<�"}�����8�= >�P��̒�9�	�C���9x衇��{_�-o�o���5F���E`�ҥ˰�v�dQ�A��7E��LQ[�%�p%y��K�����K�?���e����k�Oi(�(G�p�n���[�c������կ��-.� �LU��#8rq�R�X�Z�E��jn�d2cp+І��%o��GEg5��L"ШC�s%��\=K̲�2���ּ)�w5����d�(9����2�@#-z��(���&��v@��
�P�K���*�Ə�"���/��!+L����d2�^�dt�~��pANm�u��B0�(<����0#o�ߕ�+p��!��.\���%"h �^o�p�=�Ǽ�g�;C_OH:�����ӎH�8d�ѮQ�hR@D|�j"���0�q)�I7�X�ߜ�_�m̩9@����7�D���{�M��e����IY��L�I���i@�,V��#9��!.�z�"Ơ���� (`}0hJ�H�{[ܵ��A�5#L��@n:��QɼźL�gt}��nA	ERI���2�רF����4 ��;�2��̃,}]H;�s���6'�]��=��$�4c�V�2((bpt{\�rI'ۋ���"J�6�XUm@��wdk(�=QĠXK���|�~1�S(u+�00����V��)��<�L]?����کN(}'I������Z�ѱBY"DTYj�:��*� �ݚT3���j�7"�o��Dr⪴�BH/�P$��s�[m.୮��1ܼ�1 Ҁ?�������u��v�ylco���Ϲ���R�#��Z@���n�Z%݋hɨ�������M�V/�/�u�O���8;�������#[hC��#��;�͑��!��i����ϳ%�]C	V����O�y�@{��E7�z���ʺ܈!���oІ����-��
�y�{���כ�?�[�LߑY	������^��׼n��&x�ϾN�>��B�j@���:��g�����x�Ar!��!�Kt>��<x��w����1�_����S'�8m�FX�����(u����:��$M@(j@������v�eY�Y����/ ���*�R�j�3�,�\^`�Ėf����^��+ѭ��y��Rm��Y;�j�*���bkXIő�����3$Ld�SRm��������x�3ej�FzFl^;�+]�JW��JG �JW�ҕ�t�+]�JW����d�X���N�ԹG]D��(R�C�7��k,����T�]J0��]��W-����r�Đ�5�D�D�7� �R�*����o��z.^�?�c�Ibr�&��G �?���G���,� F�眎�k�,�yOk����G~~���!|�[��y�k`�޽��C�,I�S�zɧ��$	g���}�<������8<{�Y�����9���4����1%vxnl����*,--H3�L�<0j�~$g*��%q��qƌ)$`�g����oVVV`��z��n �.�8R@R�&�R�sP��r0#b���5E�g�|����n����=E?3�5�d��5��NB�X][�(4�����Z͘6��a>s|R3��
F��6����`]�u#9�y>�zJ9]	�EE����6��S�\n�����)����r! ��ѼIT-�lmnS/R~\` ��jR�AA2� J�mP�[�m�D������z�`_�9l> )��`��+��E&�0��)�A�7�+��V�N3���T,
� ;s�S��t�D̯�JW�7h>�}6c���?������Ý�&�Z��_��}m`��F2̕�?��s�q!���@%�+���
* G��Hѝ2 �.Gx���a�#*~��b:�+�pg7�h�]07Gp��?'r���fS�R�]'�U=�V$1�l������d��h��2��F����K���<��#����"�e���[�HQ���V�b"V6"�F��$�?pX"�!^Vs�
�21J&�
ArVK�e^[>}ي��+��ܤ�)�]�eVK5��@>tzI�l����۠7��2��l�9��EOe��ײ����A�{k���6��D9�J�1�1H��T+�e�>Q��_�+��Z_���mŶ�Φ�[��ֶ�P�n�_�NtrJС����Z�=��m���#��˞��\�@���9�<K)<e�r)g����l{m�����������nΉ?EW"Оj��$é��������&�rˋ��J� M5��#G������&��qM���o�{ｗ��@l�Fs^x�����'N4g�E8v�=S�^Ei���g�w�^�ɟ�	�{�������܁iG���{���#J$R5�mhd��bZ�+���M[-����|`bm23�{<+)a����&P�X��0� {J!��9��A�*P����4�E(�
|�J��BHPjb`��o��Pr�� �gY�I�B޲d�S���ar��ʁ�+]�JW��Y:@W�ҕ�t�+]�JW�r���c�U�rĥ�rU���wZR����:3O�Qv�g^*.as�)��ߡ�ܖ��n~f�[�9d�[n	�U�N]n�ީ��A$A3�9e���`DU@�#�7�����|���j30��C8w�E�W>5A=c��$�I>U��܃�-�rA�@-��o�3z��}���W�C����uǮ���ܮ�Ŝ㘻y}}676��K���OS.�$����)dl E���Yf'u��gv=�S0$-��j��O��?��ѣᐟ�� ����>q�cF"��]�<@�$f{��9m :�{���K`.�.�;b�I��䃳9sU2�ttD�Qj6H9���Y.W���d�>;���$�?�(-�LZrz�C���������
�`�:�PCȳ'�%E$�[�#`���^�U���$�g� Lѣ���]ռ{��4>�8ɗ��s����¡�G�����g�>����܀�M#�0�˒�Hd9��9G�c�_��ΨN����h4d������\Q�v_���`�6t}G(��:����#�S�v�|��K�Zd�f�����ܙ�7@Q*���Q�+ `h�s�� ���� ��IA�7
H�0�����M�.���y[=M����0;K�����b���4ʔ����?k�s����b�U�%H�(�T��ZU�kz`ы�?4���8MD�
lK?Sڊ���K�0�u}�#�#��RI�\�H"755�x @������"�X_f��b�x.����@D�f�����[a0���gO����c���!@[���xc�gd�����>����T��l��-䚬6Xs6[{DE�I.��Jҹ!��(2�5�)I q�T2H2og�&D�&(�J�lkgH� ��X)��o٬���A(��F�`䔧4�x�r�����d��Y�{P8��~�[����M�b�D ?g?��t>d��9���p���f���vA{'�9��I������~��	�I�T�D����/
	�����1��]l�|�Kݔ�bk7�v?���N*pf�/uU�V�l����ܶ�;� ��B9�XZyw4{Ҿ��W;���s[�OКS�--b��U��p?��'�'�1"�6���у��?�������ԩ������5��M���L���o����^�*z&�ae�x�۾~���y>�@��~��Kף� x��x�Ͻf��*M������G~����B�ހ��Yc7�����?��?Cj8h��n����Ɔ��}gb�*�]<�D��55�
�?�m��E�FO�JT�zLa��<ɹ�vR�#��5������s�J��(y�N�n�.�I���Tڶ��~$%�%����n�i$��Σ`�E7��P�x�DʷQ��ؤW��(�!��@B�4M��U��3�<���ҕ�t�+_ѥ# t�+]�JW�ҕ�t�+�b�8�3P$���;�	���*����/�4�Q:�8��%�����|�Z�n��b�Y]w^��Nd��]���o>�a�tM�K���/��� ��ib�������Ԁ)ʫ7����ܫQ��R�w����++��rM�5���Q��z(SЇs/��˗/��>&i �DRJ����^�מ�"�j�{� �;D�T�3�@1F��3�����7&�1��l�H� ������(���W�h�ȉ^��x9�s�b|��`H����<���;��.���"�ގ�H��dQO��=gN=������hQ$��j���"y�U�4��By�!`<�&��� G�	�,y��h�D�o���)K��O>J.pq�7�����5����N�_|�A8v���8�{�y?KP����;`��1Z��LN�p���V 1�4����J������_I���%�K�i�*��#W�m��:���u�ӞD��Nh-$J�Ѭ��5K-p-D�(g�&�4���70 /�B�*�zCO�q��# hJNRxWo�U���f�e!xIy��k��O����M��&m�y%d)@	F� �9J�(BMI�5ظ,��D
Q_�`�$�<7룠n!h� ��պ����K�� ��&�EjCӘ��.R
���/኉45�-��*���R��\&���?~=\j�6+
		x�q��W|��c��h�K�,B��N�_�)t/c%�k��׫�DgJO�M����J�����B�L0`�в`��FP[��Se^�^Z��+{��ӑ˽W9L���>s��V<�z[�LF�ځ��U�&��D�*]�B���&��_�\�ڰ��z��(�n��˃���2y;5�>t�MV�\�����}(�%-����q���o|s�#U�z�:e@�l�Wg����= ג��<�W��o���r�7�F�L��E�{����5����r;����/�������O����~��^��{�G�Bx6:z�(n��Q奱��~�	�7�����]6[����_�������"���o���Ξ�!` ���XV��0�U���=w���gճr�>���,��`L'����.����LD�[n��躈eM��E��J�Rc��F�s�4�2���ʜ�2Gl��lw�Y�(�nw>��a�4s�U�������=J��̖��V�_r�w�+]�JW��� �ҕ�t�+]�JW�ҕk���2a�Q�W�9�Bqn	z��M�NH�?�y��{�����2`	�3�Y�ky�������b%���D1��
����$9
�Bt�"`����ϟ}9�ܗ�{��Vנ��Z"w�,N9�G���|�w�
,���T��M�����Kμ:r�8�Me���d}�-�A�Z��9"��Q�~��y��E�� =���h�Nr��%�_3ƽ���
����$�����Q�1�%D��	�%�Hd�yx�y4'{%�3�K@��� @n��o�	m&��c�F2f��z���n��2�uۯX]����uL����$�_4�E
P��X��.e�_]Ц����;��E[F�f� #1�x25�� �����)y{,Ҽ���#��W�Va��<��D���"GQ��| ��@)$0�Ĕ��<9ֱ�����M�W�>0�r���8Y$���x�3��/>\��w49s�'@�����}�}��ABÞf��z�����)���a�����E`F���I�X+%F������~����ѵc7ۣ�HiΕ.Q�8n!(@5�2�c4�5�-S�	{*嵯�"*d��;��y�o�1e ��c�
�I;8ǓFgfI�As7�_@��6�[D�(̿3�/�-Ʈ��q"@�m�37�vc�)�,a��� �d����P�P؞������T�X\\�����sZonn��}�H�e��*ؿ�"�i<�ض(s[H 
��6�"Q[���яM�;���Q8���dQ�F ��sF�q�&�B='��tM�P�(�4��!�3Fh�4ή�UX���B{�J
�P�/��I �(�>�I-
�OܿF�+��Z�݉&Jޱ3��g�C�[󒗋����s cyI3��$�\�m�{��ο�wmiC�׽i߅d�V~�v��F!�ɥ_�kǎ5:W��2_�V����Gj$u��/�a
T�����by��]��GքN��$61:�~���S���Sd����$ǎ__��5{���;|��gN¯�ʿ���鉐�J�H��3�Iϟy��?���w���ko�1Br(�;��$�A�p�<�0<w�9�M&�t"j'��pϜ4���C��<�y8~�8=|���7�Kny	�={�zcZ�Wd+{r�����\����)x2��*%g3�r��z�ʞGDL$����sp��slH�spg2U`Qց�9�!�}�����汝[E1ˮ��n�ff�7'�Y�� ���Ge7g����g���2/[E�m{��X�B���T9�97�f,f���ܖ��JW�ҕ�|��� Е�t�+]�JW�ҕ�\�%�#��Ź�%CA�� /�ι{�8��9�V']���V��F%�s*�$�<��Br<�X��Q�N_o��.����PP/uDk�`�@�)gi�#�����	���7�`�'���� ��"�H�"�s�C0�g�(w?���"�Ǘ�4$��8*����c�3�*.9��)��t���v����<���Qw4��K�Q)� ����0ƺR9;~c����>�� 6�C�*c .}ηnc�}=�D���\grh�I���QZ�k���K7�,Ⳓ;(�G���뮃͍u�nmC/'��^�'��Ƕ+�%P-`�9�#�1���s��kd"`�[V7�L࠾�z'"zD���]�2 �㲼�iƑ�	��g�Qj�':)���̐02�T���g���ۉj@Ϙ���dp#=���C4��m����ps���a�'�i
�-Z�6�?����l?W#{�(��Ur84/r(9՛�---Q$�M7���s>|��[ZX�յ��8O	�?}�4�~�����#?ۓ-���IlIq�k�r2ۢ`��=J�x]�EŁa�Ʋ�<��}�J�L�{�2=y�; �%�Sq��5(w}H�P

�\N��f����ѐ<A�f���I�n��T�l��5ի[��|�6%�ϳ�峳��/m�}�?�3U�8�-�eś@T�]���(�#�G�)>h�
P�v�
�F��؏�W	���$,,��t�D��)Df�b#��v2��̍�ZK!+0�"�+�V2"T�CAg��m��pt
P�YIce+sd){�P��ٹ+s]�K[�Ӗ�4��b�׭!w�,*e>�d��ROI�\�Q��K�c�y�{��j�}�=Àb}f.{�k�N�̽�.��O��ێ�sۇ���U~vmh]�M퓜}��%�9RQ���z�ܪy��J*yT&��fy`���Ή�&KqՇ�ujC�l��\��6����ie��[Q�l|?(�3� �����qi�;o��`3*1�$��)�p㋚��O���C��������N����|���S�4���ŋ��� ���x�73=v^8{���7�����1Q���'�$���6�LDĚm,��jJgZ�uO?qN>�$<p��p�M75{K$�LQ$!�t6R���%g��,�d>�EYk�g� �� ]׼5�:	�@$��X��+o��l�&S��rv��������{ALE0���:)�]�s�B!1�Nmjkd^���Q�3a�e��4Rj����l�F�?z��N���|[�د�96򠕙�+]�JW��]:@W�ҕ�t�+]�JW�r��	��A�E8+�/י;��U'�w��9�[ہ���ݫN���%�ǜ���#��jB>�TvOn��Fc9���ށ-މ��]z9�j��.����!|��{��%��S��ȋ9Oɑ)@���&�[\�<�"Gz���;�F��]��m��S��.�׋�� Q�� ]��ő-��C��?�b��w�	�#v�V=�{T �s� �o��r�]^�(it4#�nY F��ױ���`�t���A�"�!2���纣������G�����I�g����K]�"�+s&j���N<��;���㦯g܎�M.U)*Y�i�B Pׁ^!h�\��v-,.�޽������[���N�L�zk� >}}(B[�97S���q:mƑ�I���2�$��� �s���\�%xu�K=�D�u�$�o�|+�{F$� ~o��Ea�pJq�ak]�
��ؒ����w�+?plx��  *V6G8��"B4������o����r�#������;�]��i�Űׇ��6ES>��S47p��ٻ��^��[��D ��jf ��T<o�;�1��W擷�^�D���E����X���q�y>'o8��`Ҭc��<��<kĝȶu��M�7IA��Fn�5��Z��cGy�Uʸ�eQ�#S����Q^�̪J�	F��J	l߲���@�N	xz�׹�`h���`CC�Is	*G���>�,��R
J��T��[tU�6%�	&�$9��gw��yr�Jv(a�?�x&D&W�:�*�"�|�����$J/I�)���"2��Y��B�`G�m�eQ�ЃA��N���m���6-���1�l:ֻ"H��SW$QL���#�u.��E �<�-�T�h�>&g��b���< ��\���yA���2���W O=q�xd����鸰�AO�Ie*��S��R:(���.���Z��5�����֫[_no�>r�.���;u?�Վ5���q�+]"�K?�[����)�6��h;U�[?�A�m�` %�ɠ�tH9��`�Ǥ��r9�(9�]�F��acwjT1�>^]]��{�����G��& =9����ƶ�����ĉ'�ƛn��V�F���`ڨ
Ν;G�o6K���:H3��~L�.C��0�o���O� ե��Hl��1��KJ(�[�Kֳ��v��(g%�r�x��s"��d����&�6�}�L$�9J�_)�=����DX?Wh/�`��^�E������g�(���w��%�=����l.��+�?� ��e��v���Fv��n��e�TmCѕ�t�+]�
/�+]�JW�ҕ�t�+]��JΣ�;H �|hx�rq��t|
���q,���EjUAMug��c���s���2��8����-�B�(dq�F�W'����0ҟ��`:�3*�S����Xⵞ��Q��3v2E[]�}K}0�:K裓����ʧ��PǓ1�`}�|Q��G ��KȽUT�H�=�Xr���Z�*�jɏ�Q�<.��� �C��B'���*���	@�:��[s�"3P~h�<�ܭ�%�ݜ)7,���y�u��	<i*�t��|mM�OB4��M�EF�i:#�P�?�	������o��[��/]�ӧO��S'ac}���'�	E�甊�XgY�}$v ���G���W���ޕ}�c�\��_^^�:V-�3���ZH@Q�Ԛ�;��9o�8t�lm��g-5]=��锕R6B���6�P� 3<kа�L9���O�Ч1F�޻����M�H \��MEg �e&�w[�e9�7�(T$�����	P�@&��F?��G ��`
&2�I��V�p�����7�t<��3�Rc:MM_o��+k��ɓ�����l:��-���F��U�9� �C@
	9:����<g���p��>��do�<0����
��ڷ����UpI�8�@7����u7\G�� 1@����sP��
��
4�U�(v|7���N��x��!�Q� �9�I�~@u��f% $"���3h	��Q 2�3���|� Y䓡�;�(�׫ ��u�����<5s�������Av����8F���	������'4�@E|?F�"�p4�>bE�D�/���%6� J���L���P�}2{�آ�6Ϳ�54m��5&#>iiV�Ч$�����Qba� 7�|#����RÞ���`s���WJ��<r��Y��_��lnl���@+���fR�KK�ӓH_��9�-����n;>k���J�\�����vg][�3۷d�C����&d�L�~�k7�R/`��K�`���R �z�����`���J�>��N�?� ��+�jk,��7��I(�e3�3خ���m5�����5������x5��x~�U��mW&��7�ꢶ���+�.�υ��HE��({^s�l�m]�wH�YZ���v|������LH�k`�ԬNfnО���@5�?��	x��ga��}D�;r��W0�ߴ�ʕ"�֙e�S���REj[[|���ݳ��0�_�|P������ '����	 � 0�^�C瀦�7r��#^[��N{�ͼ2���6Y:��`m�b|��	n���3�9+%��(	6Ꙓ���N~FUi�/�"R��ʼS
އtZ':�i}��K�	It�ڻjQ��xN1AC��]��i3ק��˺ҕ�t�+_�# t�+]�JW�ҕ�t�+�`�9�b�c6��xтs�Q1`��%��8ɡ� �6��5pcg}Pt��5�_�<�����E��?-����ܓ�7_|��!$���Fq�c�`&����0�ˑ�n�����p�-�4u�Db8�T��%i��@<J���`>i��q�μڤ�e��a����I|�)J�!�t��T),c+9*gN�;����yf�� �E_'�'#0O�� �4	�"��g��(��&0\Xd�x�t���8%2��Lޠ
�`FD|v����"a=�6���[��Vz&�b�DƞM���bIo�rbu�Z�x9�Q*����}͸Mg�g�r�K�|�*�;��YZ��F�b���c���������<^Y[�������F� �g�m���N����Ɏm�>�g1�'�oZ�8��M?aJ�����o�#G��,�+�#�i����5��7@��1�����Z�Y#�`�Gi+FC��($�i��������/�b3�{�QfO�8As�lks�޹0A��dLq���j�f��l�J ��{�5b �8��5�PD�? *�;4�_FF��d������9��VSUlV�26D"j�<{��,-Qq}aI2�4粨G`v�q�=�M�@�����_XX�1�HIlN�44G2���`4 �F��9sZ������
%�A)))�y�hkJ5w����|uo�5�aY3V�8��p��~��董��c���ڣf>a����_�� ���	$e�r
�I%��N��ւ��I��G��0 �lp ���^����3>rZs:�>��쓴o���fL�@�g N��=+K���h�p͜}�"�&3X�ܠ5�fI"Mis���c��8M~��T)U�-��T0B��sH�:�.�2�f&���χ�=+	�����+TIf'��]柽�ʄc�.��n�պg_�s�/Qǿ���E����Ek��-��k��ۄ�R�m�:�|��
L-f������V~~|�f�=#���7;W��]?/D���]�uPRx�@�mrͶ���xF�i�a/.,������瞇G�<����9�z�����VsF��d>c`Z$6�BV�3�[}4��\��2K�f��L�k<�rf־ ����Y����M����m"R�{R�b�sP-�;/�;E�HL�h��+�ؤUR'��dc�J(l�ii��\O�y���5<��-%m����]E"��:�ϵ�9$��"B��ZTsri��D@+P�쒥zd7���R�,���?�5L⓱ľ:m6��p0m��YnV�ҕ�t�+_�# t�+]�JW�ҕ�t�+�ZY �P!�y|�!u�y�\.�:�+ڞ]��
D�v��V�g���?����P���]`��͗��I�)��h��`�|kv��;)�<~�3�(E�j%��μO���^�r�h�����(D�	Ŏ�>P$����w#(�g�F2���q�^ �a/����G�-u���d��?N'3V1i��j=x��31�X���T�E��E�9�Q�KHgΟd.�����C�$ X����F�h{k��]�L<G��Xb*�X'�(���H��Q_��x��U`*� �ڗN�(5�_V@PB���ω�nStx?��0O��L��N'C��'T<��b�׾����GRr	�C6�7
h���j����������0������ѱޯM=ǶC(�oѭ��eU)Y@��+�Q��u�)�l��8x�����������`��=����y0�0�y����`���u���ex��/���>
G���t�p${���0�6�M��2c&��h0r�*���Jbp}G!���a4j^���L�ѡ�)��/Z4�P�8@���o1���-="&�`��)F�'^<Nl�
h.kdL@r���=�F�)}p�?�ie�*P�x�:MB���LX�j�n(��w#B�� ?�_V�D��V�c
�f.�|y晓DF��_ 0\������9/6�?&����lmo	��PK�t�K�@5)�V���7=R�
�)�F��yz�]���и!����E����3��m�4%Hb�0�˗/7���]M�À�%�q�@Y���Im����l����l&u����~E��Ԃ�qʉmR`ș%˥q�g+��) �Y %��#
��W�����%��kM}Tn]9wt)�sO���#T��sv�y�~���;��,�>�6�Bo������C�e^f>���:I�QI��n���g���nק����x� ��#�'A��W#\����՟��m�o��Y9L:��l��4��X����:ú~�^i*?��F��^]]������{~�=Ћ��t��>������{-u�m4�_�tN?{>�����?k�봶Y����u3#72����TN�tvS�ͻ;?�\Tś�j�I�A�Pӹ�Wmw ċ��-!ê�9DED������}��R���\As��3w��kI����2���?��x�?[�+��r����$"<q�N��sISbЯ2�Dx\?�+%Wj����v]I~دܷ��"����dPbG47��YI�~�c�K�ׯs�u}����t�+]��WD� ]�JW�ҕ�t�+]��5VF9�*ƌXj��`U��v��S폝�T���,N'�tQ���s,�'��v���`�\b�8p�8Z	��Ν��Ysy9X�T��9��4�>.W6�!��������-W0;)Jt�ࡇ��}׌�Ǩzr6"@(��3dBu��^����&w��8'C���1�D@r�
D&��_�h�:�0�e�?%���II�O����Z����I�3E��2�D>��u�#�T� o�<�E�S+Lfcr�zǥ� �8;��`\���uQB���[����:?t���j��$p�e���qiO�@N*�ʠةS��g>����Q��>�,=J�3��7�,�YA/rH�h8`(U ���d�(O(u��A  �����)�M���0E�cZ����~�d��:���.��,���"Ut`00�;��x�^���eM�Uh刦5)�J{ő~�gߚ�g�}�lp�]w�JJ
�)ĕ+�ve���Ϟ=K�E.Y	<a�"nT��	2%�\é6�|���� �/I�e�	�����n,�F(��5|���n��\�|��k��Y�,���
8XBR�d�>�I�^e�Y�KI�F����&M0e�QҬ[)���<ϘHQ�t�Ok�� k���l��y҇F���2`����`Ϟ=p�-[��(���!��^��n��>�l�&��޽��]�N��zp�f�TQs��&o'�]�I`�E��\/�0�\ .�~��K�$���AP?��~J1�(���7����Z��D4"���Ԗ(xX7���A���u���;7�t�}�=p��~XXZh�z�y� ��HD
0������������,��L��E=�����弱Kl���w9����Y:���|f���EY�ڗVG���`�<G�_]��b%�d�w��V�l����t-()@�P�j����1]��Un�\'@�*D�Vd�������v��o�6����I�Mn�r=/���r��W
���V]��ݥRE���m��!Z��7I��T@
Ax�L:'�X���u�$~�/�_���	�������{V&���^V��?{��-/����o!"*����5x��g(-^�k��x�E�RE�����:��x��=�.�Yf�B������2�H�)L�9ʑ�������o���Lb��L�V��|��m�ϟf�t	!��H���u�/n�� 	��輎{=��z�j�GĪ*���6U��H��gI�Q��Ɩ�Y�} !�r�8Q��$�eM��
�) bYϲ�+���`;'��PRn�Q�8HQ	��@֫��{uU��ҕ�t�+_U�# t�+]�JW�ҕ�t�+�XA�\U⹃QP ��S��
�[t�\�|�w;˜��o{o�?�37�{B�i[�s3*��kH~D�I`�:kK۲85*9jtfVǭ8:[�N>�T"��	\d�K�=X�g�~>�_�/x�k_q�@�W�Y��8p�P�@���(0��ⰦhHG��`���E�>pܑ�FiV�@���H(�,�c.�g�u)�uH���_/T�/�{T�B���XD�>�)9�3�[�r�"��]Ss:����c��^'�鏴\��*��)E��jMyf� ���	~f:�uP4 �&O"�9=�(��̧�䁤��X%��|!n_�x{B���NT��ؚ����x�KHR ���2R��J�8k}�Ƃ���}_�,T���Kı�q���8���6#p �sjcZOHB�) Wf8���\$�SE��w�#�1����މJ�^E@��-���BH.��q�`N���f����  �~L��f����s�/?�/E�a/�=[�ּ7ϲ(T��� P�����ڦY9r
J+P�9�v�� J�qu-0�c�A	U��f� =x����3
Ne�BL�Ð�ү
*+�@Sq�1rO�v$�����ʁq"C���4bQ�]�.`��Ά�{�K���
@�EI2\���
�q��O=�L�����)� �=����p�
}Μ>S��Shi&��Ga���&2N��d?��*(v����aq�s�ISELfSJ[��ԥNEB�*����F�֬��<Hѳ��Ŋ�$�!��
-�
6�3��λ�[����u/�:XX��))b�M�CR�YY^�~��a{k��Ga[���-^Ғ���s6ʿZ�h���#��/��Cn`?��[���Q.�՜����%�b��p���gflS��pQ��&A���
!%�Bl�F[��R���oȣ=��J��-{��K�$ ���-��T�mmҭ��20Y*ȵ��u˻�D�'0�vRh��b�ܔۧ�|�j&�#�c���c��\����a�������o��)1���K_�u�޿�^����߁��1��j7g�	ߛ9� ��P��@��"V��Il�2�@O�/
2נPt���� ��
6\���gM�1��ܢ��D�]π � <"�2?��!�eV��z��3���JTz��{��y_��$��S������s��k&a����$Q|�d��4s���e��^��u���g� ����r�YY�F� !lن�d�eS��ȅf�+]�JW��Z:@W�ҕ�t�+]�JW�r�� c���N2�/Q�T�R����[�K1�/ƒ�؞�R� �R��4���f�&:-��њ*�]E�UE%�5
U���&���f�xFm�H%���ާI@�Z��" 1�)g'n�/�FNu����K���?ox���o���E��>EQ&)��3��f�9Z/�8�m2�j��F �s���\�3�n��>J�f�$���$��.g�D�=旟l��H���xЫ(M �;��~�@<N��(w��j��/tj&�:C��͍M�z��;9+��	�gY��',�����K(M@�g"��@�W�ٚ�����%��E�+����'G���3@_:W:��e��w������gQ��T
ffi���t�uG���4�):ګ���3�|yFKЛ�M�8�LD��|��A�d�Յ��D爮USi��Dq[]V'�`�s0V�oo`Ri��w�C�\#�Ĭ�w��d��vp��"a���#�$(���>Jd�N�E��x=��y�lG�Ç�Xc���8�;�5�ߣ����?ci.��� $5CVyz^��H^P"s�
{��9H�:*��.�I퉌��_P;���b|P�%i��v��.���))��� �M�j)���&%w�T��A��>�����֠@E%�<�}D���QȰ��k�>�h�*
�i>j�d2,�A�gY�E_��Q �E�Z���v�b��N�j!a���T���䑱q7��u�Nl��%LfQkS�N�l�3�	i;��r"I�أgN�=�򎌥���%bYU�Y������@����O��zZ�i��ˋK������^8���u�Qj��h��D�������Kk�=�/z������)����7�'���Se���X�����W�КO���)$J����Kf�r�{mj��Gtu��I)�&Vg}���QҰ��r��k���&���\�I�k=�^�ۏd��B�l��5Y�L����+{����Bj@�B��ʝ���������N;�y�cB�t�$f�:C�QNYlם�R'3��7��}V� �ץR��n��H͚��'?�	��'?	��s���o��_ߜ-����Ҭ�~_��0�sk{�f�����~����?}�iچ�Ȫ�Jj:�s��w{�֙հ�bI��$�4J?�k�_d�m�DX�GRE��;֋ly'J�Ӽ@��ƚ������l�)��ne�� �U{��8VH[M?�Vع12��F!��J=T2�a���]�R�uA)���(,�b S�yL���g��ΘI��j߄l���N$���sM-���I�#))�)L1eܩ�7U��a�ѹ��U��S4�&0�Џ�p,v7`_�%gϸ�����j��+]�ʵQ:@W�ҕ�t�+]�JW�r��cU��!�9����wLB��Y�rx;��aq��\����փ��ٛ��z��� Q�C�WF�$F0�B*8�<W@z~��y� @������L����)G{�\��J$�9"'JTG�s�d�t�������9�X]��Djs�BH ��C�@_��2�˴����(u߃��=��DM�����fE	p�ɸ*(��I(�<��b :o��ga�V�`��I(5ޣ��(�-��ؠ(~�"�W�1H��$:l�8��(��c�GM;fI����E�Ӕ�����XZX��h��#+PN�m��^q��������ώ}&���#�B��J�E��L� G=��Fo5u���?ا!~��)X\�7}������~�2l�Y��=�X#y~2��Nh�~�<Ϡ��ɺ
�W|쵭�$`N�D�5), �so�o6�[�ح�_���e��Z�QX�1��Nd�_v�F�u=���#��
$�{Í7�&���r��$�K9��5�_����G�I���M�D�)�I (�yޑ�2�L�:�Y% �*]�|�$R��i�d��O|��q����L�1=v�q����VNr��RTV$2��\��`:;H���3:�[�� ��� QɅ�y�[R�U �+��+�\}����*��[Q�e7@�<a@�����8�6h�k�c�����]�@搦~�p��l�F��$�_3�D��J�q@F�.Y�v��%���@�vBȓ������e/fس$���@RՉ�>�IQ�N�Ɲր�H��'��2V$�i�����9����;��_�2"�?�"������Ϳ�k�0h������`ii���'����y<������x�p�]w�_�ko�Qc��}��� [�S�������}����exի^	���4vs*=ߒ�o���MBk>]�\��beWU���J�p WW�ZHT���W�h4���P��A�g���������L�p�u�K�Amh���M���#��o3II�"��K�m[���R��E� �1��g^�«�}���1nL��[�$�L{@�?LR,3,�Y�$ZG^Q
�s ��lGa h�J}��.�uN�P��R(�G�Ŵ�"	ϣ������$�E���K{��%��=�F�������M�=﮻��ڇ��E=�ϟ��x���^�f�.���`5�����K�6���ϯ���*{����z�#�A�߉�˪&%� kC��2�SE�W���#є�+��#WMg�.��TbAβ<63������; �S���H"��l�g`QI���U���l�ft�TE��o�J:�P�e�m��1�6gU�(gC����,"�%"�r�#��Zjl���PZ�%��"�$=V�#P.��M���8m~i8������(��R�R�/��/�/	��3þ�g|�ґ�ҕ��eJG �JW�ҕ�t�+]�JW���c&�2U�V�s��. ������l����\���������\s���kUsq0��;�3��~o@�5����C����,.-���
呯%'�d2���kkk����c��ͻ.�J�Z�`G�M׿�^w>��4\���/�������p��9���9O(:��r`�Z���E 	��>��$��\3�h�E~[\�!X�%�Z7t$���wz�!�۷�����p��O�hx=1�{�}�����)5%�:Kz�X]���ͻF�;퉜7�+&D�3�3r�f"!`t�l2�1C" �0:� A�ꝛ#�eh үQD��T��ކ�I�`����e�k$9�ͭ_��ե�SE�V�;;V���ڢ�4�sr�6M�H}��"�۴��yv77H� ��ؼ���?��h�A�*JzmJ �S�2�H�u-k(kTtn�K������<'{�$��I���l���:�zK�w�[�(F��8:m����-�� � ��٢�I>�9�q�bA�Zk��dɕ��O��ť��W�����8�H�X\Z"������~������%Zo��@$�`�����<y� �cǎ�$�͚�9���O�8Q@� 2ɮ�f'E��/h�Yms6��lS�"��v�z�zM����d��9���TZ9@�=�|m���ĶI�Xj��~R�e�h���78H���g���&��oCs�'���j�
`I���s����2JP�:Db	!�
��HO
2�*�s!�h۴3yo�t��nk����$�e��vf3��2��@Yi�=5�"%��4+Lp����r�l^#DJC��1H�A8�_o~�[�կy�=����^f�^����w�ha@�7��ڕ5���!<�����ӟ�w�	ozӷ�ha�g�</��;`��C�G�'������5��<�֯���O���Q󾘚�����f�Mz����.����'�FZ�������hp�#�в
b3��$�5���� �%�s�H<^��UQ�<�Hh��b�\嬕�D{_`у�Y֭�?��V�9�E�V�F_�M/��3��苭s�y����}�ٕ\��g��S�_�ئ(�X���z.�A9�п\^{Od��	$��"YO�S�`���3�s������S=M��m�@��h˞�����x'�s�]�0���=D�ĂOE 	 x>#��y~(��ݱ�t��@^+ġh��tf(Ҟ�6լj� d!�%��CW
��D�C��x��d�0a-S$B�rG�M��U�&�8#	bZ�����&Re�0��:��jUF�qIL��Ṥ�����97?#y$N8r��*й�����H�#�~fJi����5�� �����yE�d��G��H$f�>��LT~�8��{,H� ��k_�:#���=l���A��-�_)����ܹ�z�y{���/���R�J��}Η�/����/�ݮ��}�^��.X��ʴڱ��=�����_��������t�&7$I��Е�t動� Е�t�+]�JW�ҕ�\c1�D���P"�@�v��Gv���a���/�#3۳�_�E]y*�Z`��OX�(��ot�������o����G��C��p�$�
�׳��������s�O~����M�:��+r��4G|�ZB������w���r��%���V�>@�duu?�(����0�	�I�0qA�)ɆK�YT�(��O-�Κ� A}��s�@>�,,�a�i���&E���vM�Moz�u�]�������4z0s�x.N@������g��~�W�~���:��կ�;o��@���%��g��@r�+jG�f��FB�ŋ�#�<��C��a&�Ѭ�XS�I0�U00���
�Y��8E�l�2�`11�VǱ:��)5Jt28)s7��Å�heC{�|#�E����U�m"t
�H��)�X �
�܃<K�&@��� ��}�e�Ĳ�8�����Nh~N��8�<c:���@g��^4�(�d�,i���A�ܪ���[�����4Ϲ\��˄s}ɦ�҃�[H�-�J
�Q�H��c��A ���-:��q�[�,b��~���XX^"G��"��]L61��Kd?���amm�;v�#F��c�R�s�$�G�~q Q�������5��3�X2� v ��������ҥڇ٫_�\N���^
�V��y(M�+x�` �+��w����x0@n��-`5���@)"�	B! i�u�>��[�\��^��
 hm�*)ܘ��䓨�*]J��ّ�n��h M,#o�$i���׷T�e��F�f�L�A��_<�������x���d�</�����������s�j�^.^�����/�=G6}a��v�m4�1��s<7�|3����?�q���[������E��?�C��௼�[�����g��;g�}��7�@u;|谝9J�"�����8|i^�����떲�g�s��B*�TqP�@�<��e�5�S��������W�H����^��t�sm+�[k͚�#�@���-�Z�>'���G�s��4L�$瞘0�J���\�(@�n+d�����3�!���U��5���d��&���ܣ$��9�kw.��=g���3��R"HvfV�t~�䷏l�2E���L��5�� ���Q}���c�>
�|Ž͹����{�=��Ï�;�k/_�,s7��
�v�馪h6��dK�?���&1q�����m�t&�T�N�;;���`�SN��?'�����u�E+�g�د�w��ZJ��)z��	l�F�F2Ʌ(�%!��E� ���O@��x��VE�p��jQnL� --[�yΤe�Ԗ����zSw�(Jb=:o��٠Tr³��bl��)�(�ޚ��ь��u�>�cW,��in�!O�a����j�l�bA�����i��S F�+Z	;W&6��<��^�C]ׁ�u��*��<=�����9����kjk��T�����u�S�n�Lޗʻ��5���cʆ��Ae�2i����:N&�|�G^���ّ�Z6���W��WŦ{���)0QNZ��͛��J�]Uy��z[��6F��zs���ޛF]�\�a���񝿱�I��ZRK�	M�-`��1&�)8;&k9v�m-�#��VV`!�!+@�����h�Zݭ5R�Ճz����pNUj�U��ג����S�������Nծ������\�d[MG�JW�r�� �ҕ�t�+]�JW�ҕ�a�R�,A�(Ѱ�(E��h<ın�� ̈W�|�w��ktp�6�e\v������_�"���Yf����,5�(�t$�{sf�0�wD`�-/�n������
&���t�d��ћ�L =9`�c��"=q�b����O���ɓ��o}%��[�5<x����J;��=?���W_s5����&|�K�{��=t��vnw��%���{��/�nM�Ɯ��/����W�X]_��}�k^��%9�9�����m5o}��E�G��_K�����������~�G=�F�c?��vQ��c2DC�|U���S����~7��g���R�q���X~VMCb����lA�f�~����(�-g����
4�|l|���Ƙ�KW�o��, dd'8�A\uM�{�NCh�Q3c��Sig����C�	^s�V:&�"�ݲ�ۀg#�Șl4
,��0Z\#�@Qp�R��9�3<��іY�V�t��|�l.p:�RI�i��+|�����97�>s� �X	Cl�"U�E��mrr�c��;�c9"2��\�M$/���LpN����hD�ǫ$�<�� c���`�_�'�L�E�+0B�F֯ #d��:,�F/�V�`�5�A�0� ��r��ZK�1/�)�˻��� P@L!�E��	F2�aHu'�?���"�k������8<4��FZh*��l�(��c8�	+t���}�m�q�*)����jņrN�c��:Ck �a5Vj�ʏ����U'O�t�ɫ�!����8~�$�o���?�|�;��/~1������ِT׸������~�MD�y��_�h��|
�t���.�O>�8�~�K�o氿�7�tS��������|�������0�������o�/=��p��S"��/�E��Á}Q$�u�;�<����E�����u��"��√�[�ώ+�C ����I�y��r��I����J��B��������`Y�y��P���X�h�:�D+�-�?��$e �Ww}G��U��Q�*�˥�P��j�����C���?�(Y�Hik�֞Q�?���U���y�""&޷I�$m�U�����Mb��ߖ��$>E�� g͝����$�1��p,����Q�=��!D���c���t�J6i!���⿆_��IDM�����=|BQErp4���$xV!�"�BJ�TKxN��KK#��"��6X_J���jT�V��}9��p{9UH ]7���&�I���x�뇬���}��/�A�)��/&�DSt��e��-����.G�c�@X�'�@ ����L>�F��r_oc�ڐR�pT>��j=t-�������c��I��3$i$RN'Gh�5�2#1��y��^.�wf��Z��Ѝ�}�W��?����^�ݛL��0�߰��8�M#�\!���S]{�I��N�����L�B�u����сD3��#�z47q�5ǔe�S�}�����v<��8��2��R����'�L#�?�?ҩ�7��<!�l�t��2�"0?�a��(�����R���L�G&�����rs�G��'`�Z6Q�ǆ��!�@��E���y�_������V��GC��$4�����zeme2vV�WwR�m�,�.���/�F���ԽT�ڹCٕ]�JW��KG �JW�ҕ�t�+]�JW���B������"��uю����vɱ��iE��! �Ϡp�����Qx� W8�8�"Gb���o�rAGcOdKAd�I�ىd�D�)K�u1ک���^�
���Qx���I�d�ȱ������?y󛩎��C����f�z�
`X2�g~�g���7��/?B�r�z �_���I"���N�����^���t
��)�}r���2:�}�O�	��[���陮��Z�k�W���c���Fi��c�l��,��؁�{�K�dO��|�>�Fo �јR,���� � 1K�����h�Y]S���'������������I9�)9��8��o5׶Y��9G����zOGϘe��lR1�M^Wؙ�?1iqY=��c�O�Њ/  ��IDAT���Bf`N����!I�;Qaa��a��Nڷ;j� b!���<Fe58'�����u�f�����ႬC.�а���[���Y\�%�� ��ZF�t.�WI� (E2H�Ė&H�=;ϛP�\���18�p@�RD� ����\�\+E���L� Ts~e�h�>����b��3�����q�a��j�<��E^���6��f{\D�K�����#�3xV�%9D�5*߯ �E�k����n�u~)1�+EP�����mU�Y��e� �_��!�V�t��'խ�� ���ْu���9�( e�=��a��-\� ������Y�n����q�d����c}����%�\"����(}?5��� ��rŘ��� 8́��n���<G�#��4����e��v���si]|1�3?���[t%a�p��ӿ��5��yC��;[�t/H�Y�¥��X��>ztn��zxǿ};���S�c�D� 2-�u��9�$�*�HK%�*E�9�1X\7fB���ՖY�C���z#c_�a����%X^���1��uZ/p>��ۇ��}�۟��C�Ikkd?�Q�/9������i�i��ϊbt�l�b68!�ں�6b��Z�㎗%����[[��S��p��4)M���j�\}��8���Ň��Tw&�I�'�&J\h�����h�1"A�|��^s5l$ŏ�͜���T�Mw��ez��h{�A��J��-��4ސ��Ƨ�>C}U�8l~�|ZL�6�#\�H�9n�*�7̮Dq��6�Ś��ŊH��p�1JkU�����6Ҟ�z%���i+���T�W�ډ$��>�)�C�y_.�LGkdnM{�{�n���s~�����/q���	1]\CA�q^թ�st�ק����~	l��u�u/���e����Z:�hze��I���Ѷ7Q���G�B�m�c2@?͉��<Q9l<L}�4N���Ƹo��x^%EL'D�Q*���އ	����xo�CPZ2�N]����I�o?���˗aN�e",#k*dRy��2U��z/J7�OAŮzN���[�jZ�D����=����~:�r��:��~0�M���ƭ;�� ve ���R����R�y���M�(-�M�T�%�Q}�Sa0��|9'��s���V��v������B�'�6�'�)����P�t�q�P��������&lq��v���Y�	�/i@b��G��$� �+d�zi��%�P�߷�q1�#M0��0^w���������l0�F��t������q����_��k>�.����\H���@W�ҕ�� �ҕ�t�+]�JW�ҕ�YA�D�!H|F4��Pidw�3�9���ٱ���C\��v�F�n:q��=��?�Q�Rrp2�)g�)Y3���I�A���萎Ad8���#���{�:|�c�g�z4'�u�^?�s?O� ^����@
��<G��*����NZ�����o�?�g�DN�c'N�O���#���G�8���O�뮃��}����$
	`s{��(�����lo��B�{<�D ��aie�WV�J��%>�Q�N@������`*�A9����t-�@ �xiH��HvT\Y�ؖ>"욝S^�k�Om�8���w��߁�>�i�'֭
��5�`F�;��`/�EK���x!/�+誀A�`��J��� �sw�G
z�ygd��"I��CZAg$G�o�%R��ehRY��8R�r���@S��*��G�s�4�qj'���\��)��D*MB T�@�S��Qt�9r��|�W�(2Q�B�vZ���|z�iA�����F>��p���T�@��$w��qɓ��y�p�׳9"��R�/\�H)2*�W���t���.\<���z�j�b��t>gx}'�y���h�����t.�?�ذ m�|�r���d"���
6�<� �A��e[� S&i���y��9'��ļ�W(z�B�������ޞ��"E�x������Z�Y3�Ed��W`S���Ņk�bݒgt���9%�,�rQ��%Ђ��+�K�i?s�E��7�;9�&�V����Ąs��/y)�u�]�Ms�G?�!������o���G�WE��&A�*��n�:Q�h}��#=c�u������y׷i ��qm�c1��l��Z�E�X@���p��Y"�89�qz��t�&n0��pЇg�y�H�����`��r�h��$���CA��h���!~r�������YW㕯�MUR��_��Ԇ67��Hd�F�a&�9|� �;#�a}c5��fj�)\w�M��v��Wa��r$&��b������Z����U1XHധ}���*<��'i��s�����������@ o��G����7�p��xќNO�Euʗ��
� <��:�j�M�q ����R}�<P��BQ�{��^��sڷ��,��XS ��kN��gN�Ǚ���`�vΣv�-5���1Yӳ�>J�/�,�[��[�y���ǟ��>�Yx�G੧�Jkݔ������Y1�H�9A{͹�P���3ϐ=���K�@�����4�o{�m��qv.m�hz������������7�`�QZ�����E���;IY�ᜀ��J�a<�6�ΫdNM��J�S�S� ��R[?,9��fն�R
«�_td��ú*��AفSX)a���M{yB��{H����*O}������i��j	H4 �)
+���$�U�>�]7�ͦ��+!�\�g�y.]8G�a���J�a�T�4&���T�'մW��v�\4��=�&�����K�&�7s�eׄ��j��ab�I�����#���d�B�d%�I`&�yl��i*�/�K~�T�/�d�w �����ߕ\���&�۷tW4���]@��hr�T@x���hz	Y�Ql�L�35��+*"��)z�[�H�}@Vc��ϊ2���i>�w*�~�ɲ��н���=��[_�G6ֱqy8�iOҌ��Z���s�������G��K�P�!t$��t�+e� ]�JW�ҕ�t�+]���T��<F"H��s�dP�M~ �(b#�y�]	V�6����9C�M`𘣀�T�Յ"��T3��	s�����ŵ7ʉ���=1����25C�Ω>�����W~�_Q%^����#9R�8�g͌��F0���ls��F�a'xOr�[?
?�C�%|��`w֏Im��Oמ�	�?{�z�)hf3x��'�Ʉ��#��!��M�"�3���V���t�|
��>�c���E�UI��2��ً��|�ך"�P����8�*����q@���x�N1�HEBF��d6��埿~���99�)� <I�S��Ay��v�8#��]����t�P`҉cp��#D'N7�
V�.�s�ęM���
;����Ґq�_6�5J^t��aM[��1�
gp)�@z6��ũ��� �o�U� ���_�k��!oOHG`�Sie�紖m�R�i�z�Y��]gO��c�)�]�~'�����88��e~z�d~�4N��GK���M'4�������y8�9�M9�����M�4 'N�|甎�;c�yUB���>9r4����=+�k���{H� !{t��Te��SL�~$�K{Ye�CTH����¤jF��d�E[�wy����3os<�AU���_�H��CǑ;p� �j�:�I��N)�|{�������`� AD�ױ�k 4-����ϫ�����b-�C�៝�J����>�2`(j�m�RV�` #�q���0�Y�����:l^��$��ֿ~ő�L�ᵘsH�Jv����s*���-g}�@h�\J���݂n����Ȯ/\:Ϗ�����.��#��8�y���Y��_7����ΤkQ�;�~׋��>�ax��_�믿
6����Tg�q���Z�z2�	B:���+��K�@�xl�+c<mp��A"�I��uE�G.6��������K��S?S�a�Hk9�:�U��N��pN���� @�r�WU�ynoo�H�<�F�C*4_���Z �V��޴:J	2�^V�!��1�Փ�kww�Ɖ���.���� ��P���tL��E�_���.6F6���R����熒̡�e��ʪsN�!��V��������&�M��:}7I�;l�)��3G����1%�U(��+l��^̃y��hg�1i� �^O���._ځ�#'I���n�W�yu�N�:�ϟ�>����N����\w�up������t:�����W��I��';���O��7���,�G6�G������6�Sz �=��8y���'n��F�"��-gss�ß�{J1r�]�B�a}���4�R��0�%+E�V�p����aa4L �30`>�i>��d��מչ*ק5�@Z�����aДA7&�ƶ3{s�}E�瑁��h5���N��R�/q�<N{�������2�mm����`yuƨ�i�c���=�����܋
 H��S`���ېҁ��
�k�}��mT�8{��?�	gӿ����G;��
 H�"T�
67̍����;�{�x�iTd�	����II���[d�A�#p�LT����k��)�YI���,���l���d��N� ��$UFl���4�Ⱥ��,�$�h&�2���SS<��
%�R[�jFM)>2�� �L���@נtԏ�0�N���:$+TJb��(hG���L$���^�ٌL��s��w���i�ɞ��\���wԸ�`ra4�͎D�n�u�����t���p�,��8�m��ҕ�|��� Е�t�+]�JW�ҕ�<�J�t�ѹ�}���̡�Ȁ+Т^� 9"
G��� ri�$�&����$8j���J�۶VL�����,6ȃ�ӟ#��������0<��i��^]]����e�#?�$y�N�\uM��+�{�_��גLmt���B���3���z��"���ʠ߇o�~����8A�$��t��_���f��~��B�(Xv��w�}��c�:�8 +r~5�#}>��O��"�s��?^��v�� 9��x�i�ݷ�N�9a��j�v���N�H�� ��Q��r�7sjs���$�%;f���.oR�\M�� G���������+����5��}���{;;��oD-�M$�������%T؍ڄ؋�s�N�3.j�o:^�@H#�\�T�͙��I��s���� �H�E]yx�SK�<BᎶ:g���"����:k'����4jX���a�o㍟#��� ���+&�9d�#�2�Qi0Ձ(9�9�)I�c�rJ�!�YHd�qJd�Zc��ݒ���d[x��ώC�	$�|�T�c����G�+�以|վ �$
1}�����
'�G}�c�f���|�J����������^i���c�y�ح�֤��E����9e4�s�N�!�BB�Oѹ�9�+n�uʷaz7����"�+@x����#K��_4��P|�
e
n6��)@�|�Ś�[wpZa��� A�L�/�K�>�D!��	���{NsT;ɯ�`�j�2E��,�򮜌%����hg�%��&��t�aZ��Q���Q�l�˫d���{���!�Գ��^���xN�zv�wagw�� 麫kp��s��C�K�x1�x�Mp�/�~���]��x�K_���i=&������i��1drU����v�q��ƈ|�r3�aW��2��Y�ʫ�k���~A���><��㐦"aN��(�M�?"��B� �y�{���y�&�x g�~�]b���g�A �5r]�QV#rBl"[Qt�\�Iހ�����ϲ����I�oM�R��͍��+b��=c�C�IC�h]�lC�X��	Lqc���:'�tm�N���u"Yo��s_[�$]��9@�K�L�x�������/�}��Uڗ�cq�]���w��OS�bD7����^]Y���"�e���_}+�Q�r�o��߄����������"��_���¥�6��g�?������T����*O��c�<
��ۿ%�-��3�9����,��������lF���>橮�fo�}�t�O䣽�=�wh�I���m�]c?�T>�$�����G���$�/�I���w�su���Y7��Fq�Q���8�����XMl3$� �	S�9�y�ڹL
`�+K0����ժx?xOB
ԧ��gG5�9�+�����} �$&+�B���:��c(��mC�O�g<��F�����֢��fB�s�6���-���#�9H��X���N�NnM#��*{nT�'my�Sd.�ꏗ�QШR�r^%�E} ���o���ƻ*U9I9��>O�ez�%��֢����EM��b�b����@9G���e~s<;q ��� ?�w��������vF�[q�G��kCx��	<�K��l-m�������������Ԏ_L'�I�j�JW�ҕ�t��t�+]�JW�ҕ�t�yX*_E�	�stR)M,��vm`���!M�m;��Q�0(�X�[����:_� u4�Nq��`84@��^�ʿ���"'�l2�8;QQ*�c�9r~��B��e�yh���z��ަ��I(����e��'�;���p���
`;:Qw���.]�{����i�w��q{�9�0Ǧ�i�S�O��8J����F�����DTP�<���_tơ�3�˜��	�ar�ⳓh݈���M�c��i�8@
���Tsl���O����o��w���!�u���h8�'�������z Ë hq�u��3O?��T0̓���L�[���&2a ;p�9j���t��k~��((��%0� �u1P��5 ���Աl�r���T���R������NZl���K{]�������
�9�t���1gi��u*f ��-�3k��8e'f Ŋ��M8r�8�(��'Pe���D�7�^=�I�NԚdikvGmgdǰ���}c��<��?�7��"����>��(���y:ƥzo;/^����1�?���*%} ������@�T dbހ��S�h��7�ҀM�'9_�>���׶��J�PA�NZ��V%w�x��PU�ga�����9��Iʶ��E�D�Ɂ�- Q�����7�6��k�^W�*.�#%DXJ��@��p��fhC�h��tL8�h\T�����Ḡ��^#֥]���C�T
8ϓ
�|[�[v�j��[�+�.�cO|^���	���چ|�p��Y�gM�������Gફ����"|��x#͇W_{L��G��#����>�g�{���{��~ ��[_����X�f4����gͼ�(�����MQ��[�R)���[�^�^U%��j�.ۺJ˞�RJ��b�&
�\����i�;S��ԩ=T���W��Im��✣X]��]F��-K9?AѮ6{�������� �ӽ#�IB4\���os�F0��,�mJR�����%a���֣彁nD��!3X\�� GtS�EŤ �Qj'<��}��QQ��-`l)�bZnׯdi�{R�J�z�����o{�+Am�H�D�L��j�J������ł ������T�gFD��饋3��'>	���P���j�%�����V�Շj���C�1�7�����y��<�~N?�M��;�3�K/#�z>���ɒ#J^1]�p��iX[[J����G##sG�W�'$�RFzǠ<�!�� +�˪��db�1�C��b��U��A0
�T��d� ܣW�+����*�q��ojj��2�5p9Ϳ�[;D|�C�U$MW8����S
(��y���@���Jr��5B&=Ԓ��zW�<����cN���I�ImG:�7�3��*��G@Z�.4wEN��D/�cYԢT �~��\����FDԔ`<�k���(�\էg*����b���=�;J!�_1�!*��N�<y7�L����q/�DO�ce.��Jz��WB`���TFV'��9�������CD���T?��'b
�6���dw�7���ǜ@ ����t�+]�� �ҕ�t�+]�JW�ҕ�a��GAP?�:!C2���G�����m�d���g����#�����4�v>T#�9��7����(S�y�1.:Yޒ�t.b���_���%g!9+8v�L�3r�Rp���� C��g?�98u�4�%�A ^� ��1+:�0�Or�F}��_&�[JE0��k��l^��]��9��e��D9���0��H'G P�@�2t�$����E
۪	�,�&�� t<�vPF�|��b$��3g���<@�C�w���0�sg����}pϽo��!9�(�fj�y=�H� �1���hR'��d@�`㇠��TW���1�6�2z4�������۷��� %���T�G��}�:偌����� A޷!b����z�8O��=�"��.�6��m�1����
e[��\�	8jkkky�+D��8z�r�rN��j&�i�`��(?qxS~ViW�+
ډt,F<S$`_�^�\S��7�N��FG0���:���%p�=�HY�r�6L�:ht]@�G� ���w�p Y�����.�+�
�[g�i�vV�0�ώ[�sԬޑ���>dn�{{o-�n���x�V��Z��¸��K���|B���l�A��R8mo�MѶ:����cr�/�UB<r�tԶqB��9��i�#Wԋ�1�����H�#��zSR�D��o�Qu�K�.��?���ȇ�c�4\�xn��㰻��o�@������Z��&��������F�e�Ͽ�;�O�佴�b�=���Ї�������O��;^ǎ�H߭�K���K���5�}�ِpW�qG�2p2I�K�(��]{NW��0����w	����ƃ6X�O������r$c��ݰ:��3L%���'��S8`/�g��"�E��#y���X8"�\;󚳸~��I�X{mR�SM�Qھ��UA� sW�����{Q�P�o��1�S�)\iB8�1�9�����h"|F���sD��l����&`9no��v��^��[�8V�}�ȱ�zJ�F&~D��ن��꿆��{��5�����R8z���R�^�uW��H8D��W������/|�r��X[�����w����Ỿ���h�c�	"4�T���	������wߖ��˽�܆ҿ��?�[n��_u5�Qq.��:^Z�>��UE:�$.�XY]�3���iώQ�w�u<���D��6V�=(щ��︷�=N��b�p.+�������r� ���S$����diiG66���p"�g����gK�0���B)�H� ���<��b����ޅ�}�4��Vyy�޿��E;�Iz7�Gz�8�<0H_�I{���cc���F�"��@R-�:L "F�A�,]Ou"�����E�癔L�]ϙ�������O���9
�[�}�^4�UD��!�H-�۞��h0iG%�3�J�<ٞ�ݸ#yX��M�dC:�Ȧ-�A�X�J ��Qp���u'��ߵA��濠���Cm�R?讂�	�3��+�#� 3�1��D�;�H$�x���Zz���f�t2 <�چ�+]��7{� ]�JW�ҕ�t�+]���D-.�Jr���A̅��)ݾ|�Q�M�P=V{�y	���:��۪�jٙ��-�ڸ���E��1�ȑI._�Lr��Q�{� 5:���C��`gk�yB�+щW9//�p<6@��l��j8�󫢳i��π=�ׄ�$a�ak{�"x(i8�+8�y�)�}�HQ'���L6<;�5o��x���{��P���t������`��T��|�}�i�)H�D|�s��<r_W�"�vÞxtV�9{�HX?$4���Y�7�S����7]U��d�8��;~��>�� S���h� �˱�����y��ew�+̱�8�k�G�}�7�A	���<O��
�*� �UV��"���?Qq�\���K���'ݧPT g�9�AƐ����(Ƣ�Aܑ6^�Y� �jր 6� B�9�>���}��m_�����hێ	/�D��X����gy�Q�l�Y�W��*_���a$������T�j�;�䀟��n0I]�+��ۃ�/2�1��A�l+LTQ��J��b�_6wv@S��lc.��`r��QālNn>��Hu��}�_z�r�,.+�\�|y@�8D�Ғ���z�\����V3,�r%/�v�s��5�g��N�g�r-k��D����(̈́���F�=�_dme��&'����2\ݵ���ܿ��3��v��LsŒ�A@��ȅ`TZ7�z�i؟�S{ⓟ���.� ]둇��}���SO=��/�RZ'q�GH��'?u|�k������`}�\��C��{;{��7�,ɓ���Qd/��[���0�����g`s�2�y��)O9���)|��FnG��3�DI����ŋ��׳�r�Ҋ =�|Y��ː�>V�䵍��P�v�ύD JQ���� 6�y5�/2��"��s<��{<%s��Y aR_�^�5����o���9�{���>���yT��vj?�9/fE"�?��u�O�sݕ���G��['м뜬����ENs����D�G�K�<��
r}R����R�hkU��~�5뢪��z>��\1%~����~��'?˫kp�m���_~������:+�{Mg5�lo)�#�0<��#������8���gi��a�?������~^����;��i,�J����ۻ�W_�|�O�}Z�v!6,K��N��է~�o�W��u�]�`�4�u��g�U�jD�\��\�����[������9a����λ��4O|���dC8�Q�{��%�0E ��?|^/��ި1�d���cB���8#I
�<����R�`�-�y_1��xy�C&  9v�u�dX�;�3_��<�r���;ۙ~DiJ0�z��&��!�drF}�&r���D�^�h�dO�]�S��b�h��k��^�r�8�L��.�J =nA9���e.�!�� �6�񁆭�1Jui�(G5�<x~_�9G�+) �o��� u!%�� �8��L"j�����$��+�.����y�*�ۙ� $Ii����/d6M�'v[*��ԡ
*�@C��}#��xU����+U���~:���`�����ҕ�|��� Е�t�+]�JW�ҕ�<O�s�j�ӯ�J�D��X((���s!;DK�}}K'^|v���v��R�ގ���-�JTKhN��8�%	������2AgK#�*���A��$ǹ9��i�A����&�"��R�]�܄)J��r�A�����3L����XZY�v��X���MJ!���א��A�@dn(�`)0
���3�Q���P�:4$��z=���H��?v\b�j�gÎ��QE(a�$RJZ��M.��;�]ۂ"�R;�JhHTՔ$�9�/��� %XO`c���%.�)��rP�a�� ��n@G��!ES�%g>,8��)�گ�Ź�G
Ж�TP�,(�L�
N@=�<z=6Z>�=�� 9Z�IT\磁Y��.��E��X���p��e��@����|���؄�7	DwE�����ZGr�b��d�3gs~�h�[����,�M�(J��
J���MNy���/»���d�}�;OcdF����4�]��#bOC�3")1'?��S�>k���-#l�8{ۑ��z��-���2G%\�5�I>��f�����l��T�(�#���l��&���l�mT\m���۶Es�x��qX��!�uN�\^CmNHK�����m���<��
H�gtK� m_�yu:����ri�$r�Ok�<����=��]�[���O`^�
|�=}��ix䑯���R�|��<�h��%�L1��>������>\'1� �&d�|o�/��_����W_u���Ň�Q:wc}�r`�&���&�����Ma:!p���\�pΟ;�јik�?-��c�m��Qp���J&[�C?W�,�4h1�/�\�������'�>{��#��I%àt0p*ۮFf�h������w�5to��b�E}t_U�u�/�Ź\x_�
K΢��DU�8���QR0(Q̐	*)oX9�B�B��H�E���5���mb��Rwz��kMM	�h_F�ھ� bH���6W��1G=��2��&m��h�εl��p�X����M�ϸ�y>����`�r�g���4�F���פ�]S�p�G�?��c�N�I��]x�3���>�I^��ƹ'(��{iYi���)m.���C����_y����W!�Jl�lm�=7�#&h�	�#ҜB�W�ӟ��E���å1�M`�d���A�Eȧ�c;�=�ލ􉭽!��V���`{"������va���¡��<�6�$�53QJ�<�@T/�A�TKs�-��G�hN>s�<)��>��1��	E8b��%Ϳ�����qD1�ƕ�u��FNg��+~~�);�؜����+ �bG
M��C�7����M�����f���K���,�~f��m)��dK<���9U�ɿYX%�bBE/x�J���#	�?��F�}�vtL(uT��b���V�+Q�½+�۽!��Z��WL^eb���p��Q�Zd�B�u�c��*���[U6��[LRG9&�= A;�)s�����߂���xB=�I# �eߏ���^�ҕ�|ӕ� Е�t�+]�JW�ҕ�<Kc���2X�p��Ȃ�Y,�Gq�bPHr��]��mY8�s�w�����`�cԇD��8W�;��%�	#�]��`�H/�����a:����N;S; q���� ���
 G�#���|��,�.����'N¥�]��a�PjoLC��º�Hр���8t��m�gj��ԩ�#�0��K�Q�Nz�u�����r�C���8Ǩ�(�#
n�5IJ�B�;�#�gF�^��0:�5�}NF���Wu��Lk��Y�2h:�t��Á��*Q�x�q1gA�V����f����" ��˘A0 G�a�J�a�.�9 �K��gI�@��5_b>�r���4Լ Ly�(��ٝ������AxP���s�h��9;DQ�+�(�H��F�m@�|��M�ڥ�y�	��H�;���BҘ��mE㱞��2@ `);�]�)L�C"����wJ`K�����>H���[6l�p�k_Iǐ�۾ցsܣ���u����g�\�P���M�YH��_�L�-��~���K�k�ɞ)��^�:Bq��}y�R�\�Ԯ]$�m(�O��?��
b��l..�6$���`�<�4����#�	&r�>����c�>
�Ʉ�U���ww�Ӻ�I�7Pق֣t����馣,?����vv�)�ue�"�c2��� F�F!����R��'}>��O��Q�BG#�H��q���``��� �AD���:'�xʲ���˾Z����0c�c}x`b��l����jw�GA��{Y���t��D��ǒ�����R%hx"+�����9���׆f+�у�*�A���p_���������J|���?�:
���5pU�{��y�vDS#�E{��}��59�X#���b�N�ל�����9��y�=&F��4R�W��M��|Z� ��mpv������҅�V�aʜy�z���Z��>���#���U�x)B;���4�0�� S<)���+��o��sz)�.)�4�����Nas�� ��\&�d9�Eb��� �i�I1�s	�7r��u�{Q3�hr�SOۃrnY��/�3�_�}X�?\��S�EH� V�{r� �k��?�Oa�����K0K��5݁�����0������^52>��*��/���?�ˣ�#�+��� �qJ�R�dV�!��@b���]
`��/R��<΅������*���~Bp8��Dȿ��X���j����މ��g2�#�_�]�J�rj�>�E��SC�/$E��!0�^��y�ۇ�|ӷLw��!�X�$\%�(p]Ŗ�O@��AT�*�9=�W���z�+j�JP�	�&�j�� ����<�t�#{y��|l��T�_�=�7 ����;��F"�����a�Nu�{���R� ]�JW��+]�JW�ҕ�t�+]y^�1����P$1AA�#
�2�qŏձ����\��(VOy�\u����\�����9OQ�>���� �Q.��>��sу��u�.���w@�y8�9�"4.J�;o��!�N�ݍ��U�ysk��k�:�K?r�(�����<Ej����S�G��&�s��Q�R�:�=r�yPn���p뭷����������g���Mx��g(�SO���V��H'i�q�F�9��@��;>��Q��N�0����_"�;��֨fgy3�_��E`�prɕlv�Xu�-�F���z�ʊ*�J`�+�E�~L�Vv���|�A]r8�H!?x�5����d��f�Q��I�+QR
�h��'V��`E��S�K�h% I��r{:&�PDqe@�>�A����\׎@�~�T6�<�r��q�(�D�s��Ձ�Tφ��DBD��soW�F� �9��.�@V��r���)r�C�\�`�R�a�}�
[��6�_�YA��2Ez�M�v�v=m!�Nn����m0L����|f[Z�n�<v�/��0;�]A6[�m@H�a�.�M,���Zϐ/k��:��o��},�O��b.DP���Y��d��l�鄤�5���
�#��A</PNzN�B�KL��H�� ���Yњ�è^l�'0X�w(x>��
��F2���Q��X(�R���g���\}v���~f�/M@L]	Zǭ̋.�=يI�A���@�5+HPz
�9�.�Wp,�%��yM%)��g/����ϸ0f��O��=
Jx�x!�y��)���/�9P���HZ]�M�$�1��]�=&��|��mf$�@MG��?�N#" �y��~Q�E��-9$�8���cca��R�Z[�6����lv���Hty 2�PU�W�C٣���K��ty9��p k/"˸��)w��CD�����8�q��<�6]�oޑ}�%���S>t'
N�P�:����X���e��I�����^���MM
A���}�a�*�I&#sZ� tf{" ٢���A�4�Mf��;`���Ԇ��S��a�� [K۰�~�ZW��`8��1���<P]e�?�˛�aww�j8@3*	��|���#֝�Ut.�R�,�~O�үh�⥟��I�!���]&4��к�Y=ðpT��kA~;H�M���컼������e:V���1Dp��f9�Re�	Q����ơRB��]���c�"B8�QQ-��/�T�>�;h��0�m^�YV�U&�xy\&�q�*&� )�������׻�r�{����$2�&+B�H�F�O}0�Ǟg-��ϱׯ�9hm�3/��7c���+.�\t�+]��.�+]�JW�ҕ�t�+]y���Ya,ʞcY�t^pj.w�Cb	`�"�9{��}X4G֣�#�q�TZ��x8$���9;Y"�IDYI����k^�zrQ䛴���.^�Lm��e��,�t<^���`!��`�jn�lGd�;;��x��A
 �� w�8G�p$-Ċ[ě#	$J�s�
d';�r�ʚ�'�aDK�᪫��#G7��[n��{�8j�#���o���+��E�S�A��g���U �#B1JAPhz$A��d F�`eeE��	�����JNU�[�$������y.�Rs��&s�co"rz���� Kc�Ó�plv��v][�%0�t�=�3���M:0	�K
��J�a�%w�#s'�g��S)�U:^�'��؏"��	�F�I]�`
Й�b!�0q��c�?6b
 / 1�Q4"� ���k���\����q�e�O��P�2M��NA;��+���H���*���en�U��q�>`z�&�v-o^���_/ _d5Ͻm�����5�y=�����"w-�VF�g����N�D���M�5�"Y�{��~z����-��4
@ �B�r�9!u �2E�yL��Q�u2��YQ��;yz���~ޱ0O1�ͮMW�֍^H�ю w�V�#Y�ZH,�qT>lQs�c?��}��d� ���5��5p�j���M	�D��c����d�z�����92����&���5@�����v�r%0�,W"f�c���"�K�����'hF���9k9�G9�)��S9�l��Y_	?$.���ח5@�Q��l���p����3�Xj�|>{���u
:�{0)}�&��Z|YW%Ȕ��3���n y���cZ�E�n�����Ġ!�f��ƅ�%�F�r������~�&�%Ǌk��y&����5ҙ����Q*�E�E	�jg�\�ǣ�����MVc��d�TN�L)G�V��{3�JnN��� 2�٦W�\���,�յ�湞i���,��l��8 ��9@���tSZ����"Dm:~�O�ηxW���uSQ;R��^�У������ ��L˃�6������,�;��#����S��Y���0�y$>�g*���Ț��`@*X�'{D FbL�UI0":�Ց�T8'pT;��	�e�F��c0%�E���4�Os�g�@.��Ȥ�\�30�����黾�5y�v�����`��0Rw��`���W�!�~� ~�~���^X�!�5��`���3�ވd�E!�7�^�eB���t1��a3|*���p����Fd���Р(�������HJ%i0⭽�����U�:ݧ>w��l8���p�$;	MӄA�?�a>ݟ�I����l��L�,Q�,�SW�ҕ�t��t�+]�JW�ҕ�t�yW���c�*� ����X�q��Q�v}��
�(c�ȩ���+�EM	 �,6��=H��U�F=�o���ܣ���Y��α��5���(z̋:�X��;��;���v�R�/?�3�~Ξ{�;��=KA����G8v�8|�}�e*�
z(�4��"�8:�\d�@����#�D���p��=V�s�0	'��'�%2j&�g�$o�ڦN��H�G��)Yg0��u �3��n}�m�xb{@V�8�i#R���eR9�8��sI���R���U������8���^���I�@��{��S=��f6��7�&4_�>SY�%���;[��RF�}|�:�^�g.uX,��]�9gY�T����W_�������V7�1
 ���N���8��B�Jx6�G`G�f���Te *a2�Y��F�QW�,����ҩ����0�͝=ˀ�E{>S\�9��E΍J'�"�8r�YЪ���!;��Z�TAmD"�D7�qH�r��[���I^I�\h�J�|�����ϊgU�2�M�0�p��nio׊�^�" �s���5�o]��S��g�{����Z�<�Ȧj�Ia2�˥�{{�cH�Y��j�_cvP�+�/Dg�Sc��
�ζ�
������ fO�3ɍ
�Z������+��Ik[`v4���8��#	���(��'���!G 7�̜٢��� !-��;�?bϒ3���}A]@���8wQ���ҎD�m@�#Ş#��-u�mwgϢc~Q��) 
{8�ج��72 �G�IPۚl?ھ�	GD�L&tb84�I?��5�ᇜ- ��M��5ź�c;x�u�z�T6��,ǋ�D���	�Y��D1E���i`����L*C�.!�V��5��AxP5
����+�>��\a:��_��Ӽ�>Z*'�ivDJ_����=g	\�|;�Cj/���F*y'Fٿ뤌��VO�����.U]8%B�K� $�h	+����J����hG�3�?��P@�ye/U։o�[v�dݒ���Xi� ���G�@kA�~'�E+J:��oP���~e�g���湫"2���D��ľ
�~Fz�6����?\}{�)�9�	S���\����VN/���2l����%백�[[۰����Ӟy���};����~k׬�Q�8��JJ�G�kVOA ߱4)sՔ"`Fm��Qj��~���^X��C�'�ýJ���}��z�6=߫k��&���b�A�%:Qƈ)L�o�rU�P�%�E��Gy~��*��N�O�v���^ �d�M��h�(�^�)V���D�)6�ϓ;�`� ���9Q�J�΄�w�V�瓤���Rm��{=N)��3��{ڟ�\HQ��SБZN	�=:���}�8�]d�*V}RHӑ��a�����t�y��,��$�G��`،���xi���4M�{.�g�їӅ���S���) t�+]Y(�+]�JW�ҕ�t�+]y�W1�����xw^��m��]<���E$u�

a���`�7֢��:���zOE����Q ?(.�G�l����[Gx���M�ԧ?�/_$�}����ë_�8y�8��Kuix�k�s6�����;��N��`��+��S=����R�D��/�mEA"��������Z�,���+�*��S����UN�$����9�\Vp5G���%�Y���"������xr;ཱ����{#��u���	��������!=~���d9� ��$��ކ�Ob�M"��
�r�(&f&Z� ��(Hآ����lì��6U9J�(���s��y��ul~�(��ãM��%��������1Z�߃�G���pH����9Z{��7��&�l�l/��@  � ڜ�E�ʘFj@ @s���h,���kU c R[�?�@�p�i��k�}� S��)��ULh	- �F9�
���gp_�����U2@rA�V$�I�yl1p,0�_L9��7j�jS�|UچEL*�Ȁ��
8�Q";��P�M�t�.[vخW9�\G����� ���ۮl���}3Xծ�s�ϭ-P�R/���cL�"%��Ib�x�5�Ap2�[�0�� �Av岚����u���`��f����D08r��@)���߸��UZ� �
�\���J�F��u^҈|���e�Y���w���g�y�>
�彆ؓk��:΍��cλW���1�"�l�9�j���z����^]�D���f�WV`ii@d�g�9c{
�$%�k�k����>#��?yS����3-*BY���㬲��u\�rzU%9�#I�G!zQ* �N� �����h�ƙ���7�\��t�*�V<�#�7җ�7<���]���BD�B�PU,�s"hd�V=\��V��,WZ�U����O�{[�>�)�vl-��ExzT-�:�D5TMBRw�~%Ҳ*���������1�8G��Tpy��F��g��1ׅVo�a��r��s0�{�(���!���}-0/�g��C�ʴ���(��<�{2z�e�y\���H��1�����T ��4{��~��Aڟ��i�<��h�D*^�� �G
��>��a�l0��ұ��F<�JǦ���o<���#���t����3&Y����Q&�H�9m�v'��͋�&u�]���;�p)��N��	��xts֖t|��n�>,:��p�iR]}��R��UL�����uF�C#���t��h����^�:�{�H𱇠w�|�	�������jM�:�e�1�=�N�5e����/	R���P��X�Y�@�ɐS��᫢^�aU�y�v.fh��"Ө=m��Xh�<� �k�<H�W���kR��;!T��>Jݡa�.��+]��b� ]�JW�ҕ�t�+]���T��.R�a<�~PF�'�42Сp�N��l�n��Q�g�0s��E�o)�m�`g����ݪ9E6�}��׽��H @��k"0:o8��_�a2�ҳ�'��?~������s�R������8�)�M��Z?�ŷ��È�d$�稛�u:�$�̹��k��'����mɅ̩�X���������@�$3���J�O#Nlv	S����9X�ݝ]"'lom����߿��T/��`A�2����众��>~�8ll%G'�2��@qnQ�O&x����{���`��;[��6�@�e�������7��\����4�
���q��v)A�+���s��7\b�O����z1�:rO�>K������ �� :�9�����@��֏��`Ǐ�����+�0�%zS�/@�f���OȶQn�N���k��g�E�ӽdD����ٳg)���	KJ`�+�@\��弨�4�p\�x�Tˁ-}�D�-lW�F۞ͧ�F��$�	J	�
�;��P�Q��~��������W��}U�0�	etY�� Ȟ߷�=�A+�� �N��u�p�"�{�9@VЦs�%�y|+� �JQ�hu��k.yJ N��e���AB��wIX�L�Z& �@��3(6&��0�ȥCR�S� ��a����W�4{Jlaг�k��M��J� ��W�U�7GWf�r�Wem�D�y[< L!�~��.�m	�.ڛtnϊ�������a����eqͰ�R���\�l�@r�+K#����4'n���cp��9���#���:��7�ӧ�o9T�(�Ա�9p��J�Ӆ�lR�:��m�LD�g�E;;J� ���K^�R�n/��N���'��}�nz�%�o�~��ǿ��#�76��#q����~�y����<³-�}��A���𢌃��P3��P���Gs��2�w��RU��o�!W�;���m~��n�)��	�/s~cɱ�l������B�pC�n�3�,�x�5����9�W����:��?�2���вT�����ڢ#�8�5� f�zh$�ʤ�~���eU�<���P�>N���4���p�b���Ķ�y�f�4"X�7�Z����,HT�jh���;�h�=`���<g�\I)�N�`��P��XJ�GPI ��4�漧a��&�fBL��R�{�4���s��&��A��k�^p���׾r�w��t�_�R��O�v���{'��,]��$Y�����j�GI���Rz��G��x�3�����0G�V==�O�x� _�~��:]��(Z���H>o�����+��cat�C�{�d�+�=�<��^{�w��F^�7���_����5���⫾�W�����ҕ�|�� �ҕ�t�+]�JW�ҕ�a11���w���sb�9;� \2�n��8b�H��Dˑ�م��*��H��|Cb8B��Þ���e��Fσ ��L�G�X��l���G�����W���Ο��S"x_ñcG)r�ꍠ��SRZt4�[�Eo���b�9�������?$�;���*T)ԃ�h̑��q�sBm���I^f�(�<��K����y����K[� �u�Φ�R�h�g�+q�7�&�t�0��
Ha�a�C5���1(�Nq���HL��/|���ߡ����b�v7gn�{Bi�U�� �S�F�˅/�%; k�Jf)A�|��D�����D�U�� ;uvK�s�ﱯ�5�/m��+��d�Hp��7�G�F�IT)�x�]p�����1خ�����#�g0@�'�(J �N�Ł�Ŧ�<G{i���m��?�"��u4�>_Nj'���qĠ����#G��?�ٟ�յu��S��r=��ZY�xMm"N}�~#����bz$�KĆY[�;�~~��ޚ���ŋ��q3���ub�A�2����9΀`�/h�nQZQ�Q��M�Χ���o�b	c����yv< ��I�¹2_[ՋW�1������c>�t6�����|0��N�m5�	�=o		��ϝ����v�0`I��b@�w*����B��9XB�|m~�� 9J;HĪ�01�l[ƪקw9b��H;�DZOWԯ�s�~�uQ%�(9����)p(�J�u��6{(���\\w���P�J�T*(۳��s���g,#t�O]�	%*�xѱ��ٽ��_�R2��4���
Fz��_3�#2��d���m��_^YJ{�]V@�@v�mh�e����1������9�Ž���y�+㴮��Ik=ʞ����`���4N)�v$ r�2�"�M��]�E���-R~���!�> Kqy�@��5R$��v�
�ۜ�2�X	
8M+k4"Ǟ�8�&�g���֌r>��M��U�NW_�)+9�5Y�8����&06~G�� ���
@Z��Xg�l��L���ŜN@��\E���Q�'e	�A(H:_�b�$�JU$�D!,�6��b��*�LoB�j�D�]���&�[I��N�]it�b��k�ZQR�hK��k]��ȵ��D�uLz���<��ն����'W�[�C��A���������ݝV}���8f�~�
3[��^���3	�-9J6�ݝ�ln�����Ï���4��c�O�gP~��ohF�����A����ڍ��ߗ �!�@, ��}D>?/����'�I+�珖Oɛk�4�#%�'��J�ǯs����J�w�+]��-�+]�JW�ҕ�t�+]y����TT���E'����9��}��j�� �����2�tDZ E���SףF)���fL @7��i,�h��1����ц�yD12}��E���������|ՃK�.H���)�9f�H��<6� �\�='����8S pHr�Q��4
�a00P@��$�㼑(��]I�4E���'���~;N�6��왳���gC`+G�5�o�t"�	$V�%��R�ΰ�5�p�*�HR�Z`��"#Q�����D��aG(Hd��kF��+��j�w��/����+�P����g���:���ky�"��r�*8`Nd��|�C��T����h��0�P8"��m�v�(�#����?��N�1U�~������8~F�%515�=��W�����=�"�@��x,SNr����ex�K_��܃0��z�*�� �#��a���KV������V�)<mN%��ޕ����\B:"9M}�jIFJ�1�
h,-/�W��n��F�x�<lmo�����)p&0��G,���B�T~�����` �4"�%4��C<h{%�/� ����oњ�9Z9�/�E�w|g/T�1mX����/3�I���"y�ƢA�W�{=���3Ĩ$(�L�IE�h?̟����E�
�o���W�+9(R���t^��yz�E�]�ƮS�\�Lt,{�D@P�P�C�En�AH����l�Ƙ�O���,��c"h�o����h\8w�#K-���F��B�"@�gfS����W�<�A?νD��u��%�=MR�cR��á�������"�&�S�P,�j�W4i^' rݽ��4&e�Š�F������DTp@2嬦�3Vb���#�"�x"\�<�XtL�<k"��UiT�X�/}.{G�d��KcXZIJ�'!�T*	y����#ѭ�Q%f�<�,��C���y�G&-��G��N�1qic��=q�s��z�_5NHA4�d@a�:Of�J��Q���w%�'�3�S�1+s ?s�����/)F��*������q�6��*�P,�h�e՘�b� �IA�(��{&�����`{6�u(���{F���R���4����\����Q:�j���%H�y>��OQ�i���q?=��b���R��ܦ�ZD�H$���*Ƹz:���.{������i>�q�$}e�]�JW�ҕ��� Е�t�+]�JW�ҕ�<K�blE �8!�wꔏ�Y����N�*ޗ�<����t��#2��n��󍢖�`��G�
o��+}��	��$^b�(�����M��/~��?�����s���>�?w���{���;���׈@�L@gb�h$�O>~��ȷ:#1��y�?�~�G &'K%G��q���懮<�
(�%F໚���F%�Kغ9��z��1rMH �PĶR���0�������G�|$ŋ���I� K��3���	 e7ȹI2�HT �o#��s�R��YJx���\Q�W�<��` B�hP�>�u�/����+ճ|���˧��\y̘�7@!-��B��������<,�s�?��dSW_w^w�=U?/��)�Ȓ��]f��Q}Z}��O>b��A�RS�S>h��FSm���^Z{0zaPU:0��c�(_6)e8��mE�Z^Pz��`8|屽|�<ގ�/~�f�G����G�z���n��8�+!���9��*�u~�����1Y�#�	 :�$7~)��0gFV�NL.�\�����c�V��mY%���K��l�ڵL8R�}�<�љ�����7������ND��_Y�*V���V[bO�F�4�,� �dK<��m�a�ǯC�bm?X�üx<��y,� �4�z�ݛ���d���Xdm�v���Y#2��_${`W3Nw��o���XO��s��N���F<���������Gz0��Z��Ӣ�"�4���]��ʜ,��@�����F�\Y�W��\	f�̑ă1�h��D�{�����9<�P�oQkk�]��C*�i�nF�+�X��iD<8{.G×� ;����:�+:�lT��������s�am=��BeYe���x~���sLK� �����l�h�]3�9��?걖�ĩ�X_�r��'�!?����s�F [#\I�M�?�E��kI��RUf��ti���^89�Kcg�9�M�^�xb
�4I��"�
�;��T8��Q�2:O[S|g�`7�!B�U �,�2�0���U��s�\���!��
�F�_�f�iQr�8��&n�t��#���}��������Q}��/h��3]A���Zee�2�Z����#p>�����q壵j�Dv���Q���E�'�^�E{J����z�;�8R��x��'�9�u(ۂ��W�l]v��Ӟ�������=dF4�cA,EW���7Щ3�\�Vt��(f `g\Wt^��"��:)�y��^é^��ST7�j���v2������U�T��Q�� P�J�*U�T�R�ʃ'dz�J�ٰ��80�����` �l��b��܉�����._�$�Em�����͑�^#c5IǏNN�Ν;p��mx���ޝ�p�ݛp������p��;ً�C�9Ґ��i�]����ܹ{���8|祇�K��pt|Q�j$[K�z���㏧��H%�����%RuU�#P�)o1''��dp&Q��%��Ij&�� ����jA��~C'���2�d��ZOyH�� ���ad8EQ������'ފp��Ll���zݢx���z�)��g?_��8���4j�@`�=X>i��X���m���^F��2����Cs���/�������!���-����D��
�v�A=��<f "�p�v��a�{o����e b:�6����N������D�b��	RꯖE{.�+��ꫯ�Ϝ��IR�@� �]�$����ַ��ô&q��vf}:�L�Zl�1��2�+C@�'oH�����aw:�����:�W���Q��Li�\�|R $�edJi��\G���CPzO���	�K�1d�����V���G �W�<�y��|�����c�غ+-b��:o�� ��r]؁��9���l1z#3M ��Y��G��1M�J�B'L�BX�Ƃ��\�z�u+�"���Æ�H�]�Iu�o�L׺��|n�wE� �3�d�aEʠ��� �v�p�u��5}�I�ٔ*�²�����}�Ed��&,�/�ఎ9��t�Ӟ:�
Z���W����[W̝�n/��x"��ƤP���@�sr �܏���n�6�� �}��֢�Qo�������K/�V�;���2�P��f��o/g�>����֭[�������G���k�/x|u�[n�ЙN�Q�|о�MD#��[Y��c�n:'�9&�ק�ݼy�'�AǪ���t:�+W/���1���� �;����A,��bB�[���b�+5c����D��q:��q������=�g(�NhA��<�����ep�!�#�i���D��bV�#����Z�����z���[��L�;�\�O� ]:�b"�Y 
�W�M���t���>>�� ؛t/Л˽!Z�A�%��pjf)�tV�r�-t!�����5-�8��c]}��.�
���3%�����m�4W�����
NY
ݨ�v,�9��|9?H'�R���N�|�t6��
|��V�"�����L`�DC��lM�7��󑽛<��EJ�J�*U���Hu �R�J�*U�T�R����D�1zK
M�!iԫZSA7�=E��0C��V���y��3{��i4��/S�2hT[����Ǒ����h.)¸�f���߅�|�9��A��b1g'�(��M��lf��ŅZ��7�x>��cFN���W�O>	/��R����[��B�����L���GG���+��/F�q�*��*�(@�Ou�%�����G#!�w��-��C� � ���&���-B*ۉ�����\|/������|tVX��dX����S���_���z}�q���58�ۃ�_PJ�H���1�7�����߆��|��_&� Rݳ�3t����͠�E�o��Q������<��ʳr/�~s{��5��J�:����|�tP@�@O�x��� ���)����ɏ��jڧ������ �ܹw�ޅ�|Ig�4��4�(��A$W5:�X8�8��w���{M"�����Cn0[�n�y�mON*>�矅/~���h9�nKa�h(� �'��q	�p��s�y!�}������?�9=�l(�4�_�TE'd�x���9
��T %jV�ט2�lZ�~���-h�~X��޹s�ܺo��̦���sc��������d���8��������tP�+c� h�7tXh|�����~}N#��P0�F�ago��Ź�l8�z̳��;�{�Ⰴu�\�8��NON�=������(�i]�1�mv�:�6�99�B�,����ˀ����$[�S�� xq��̠��|.Ͽ�a'O�?>��O����|�����{�޻C�o��(M�i��� `$pLC�����cx|85Ƌ(�Y�����a�W�y@۟����d����r�� ���b:�"1��xt��T:6Y�2�H��1Zw��	��D2W�N��\�ˤ����G�5t��=x!��� @�q��C�i�u�P���Q��z(�ֲ��؅�b�E����O�m��m$����"�v��'_��WH��\��D��0��ȸ�A=�f�t�PLݝ�^��Z����J����K� ^uHºk6 �)͟Ё��D��,L
����Rk.�C�-:�:�]Lqx ;;3yě��|t��&�C��.�;>&��cw���_F�yc�Ƶߙ��o8�lp�,�mY��7���iu���י�I.ZMCg]t.Ҕ24..��(�� ���QYTd�B�46��}N�:8�������Z����� �*M��QV�(s��e?� ��U+�9��J/ i7��<�o��]#}��T�w�<�Z��TF��Q�J�*U~ܥ: T�R�J�*U�T�� Jl�!�kt�#�� �/l��l��@>��8UVP$�)��4�d��]�wQU�i��s����E !@�ڋ/C���#�ޭz�.���>#{�*G����zr& ؙM���&�տ�W�94*4nv~��"���8>9J�:#��k������������0p~oI}�����@���	h	 �l|�ww��A<=7�(�@��� X�`?����h94��:����`�O��5�{｛ʚr�Nt]!�p7u�D!�m�y�Ѹڠ�����y=|�����Sx����_�k�˿��0ۙҸv
 P�o��3�T pk� Ђ3����Y����8GU���ǆ����ms{�3��`\��궱> �?u5�9wT��Y�u���ղ�TD��
���ק�zq�I���/��wߣ�Q�g`!��-��G/�/�#�"��؆U�"�Z��\-	�]���i4�..`9��D�+���hh��4��90��7�h�Q���x���IT:熢��c���N����'GG�Z��,;�r�䋖 A�0�F���tKֽM;���C������>9�A�8��޽{0?����@�V<�<�3��b��H�v�F��@�>�.�W������,'�n���V���Шl/��k�t��y����=W�^�O�3����Po����EX,���T�_J:��}<�QG ;:c��i p$���6�_(�.�O���aݐb�>���t`���|S��G�?J�h�N<7��=�4��6�s����L��=��'G4'���~�`����� �T��j���νى@�g�v�������#���d����Z�(�(��S4�(@��#�y�Q�k57��~��~8�����U�$�ɰ �`j����Ioz�)��F�GN��A�r�GٟA��u�0��W����y�k�|�����.�U0��چAjL5��6��.�sY�">�����vf"6	�?��{��ʧ�r��@���hJ�st��t+����%����9�^��/��sp�x�޿V-;w��2D�FƮOk;��h�)
�7۴�;��q��ا��N/`�����r�}8<w|�*%Y��n���_�!80D��t����P�L�,v�mx�Kӌ�y<G���>Lg]t*�~��}�u��]䢮n4�1�X+���˺O��dd�u�B�?��0>�y"J�u�;b��V�!c��Η�N�b$�&q���ɱ�xzK�|�	S�J�*U(� U�T�R�J�*U�<��Z� "��bxʰE	�+����f����Cv����%�'Nm�����0�hҐ�3�{f�������ɠ�����1�-Na�Z]x�h�U�.& _�8RҀz�dk&=|����{'������؝������_���NNN�ݙ�F�
H���h4�!������`yv���_{>��fCxXc�'`��r�÷��]��?�Q�.R[���������?�g��� YpOO���/�l��K�vB������̧&�iA��w�����������`���;��?���Cpv��a<D��U��|�b㳛���3��?�s��_|����ᩧ��t���[z�����x���5�y0�)O� �̎��C��|m�o���W�s]�G�QAo�o\��}����k�r7�=�����y ;R����Ȟ�R00B��ki�)J�R`�;�.�*������>1�8��h���0H?!G���>��^�s���^1@r.Ga�hp-;}c�jR�1pJ��eq44M�
�gJy���4oӭ�c3a/�(||'��.��o�?( �J�S���35p����S� �[��mg0�=H�n�z�QH�ɚ��r?��*�5�$��(é�(���1G�bHi����6���<����Qh�B=�&]&�:RcfSf�@�r IOM���e�,q��C�!��$:x���J:m�
���[pr�.Ю�d�Lx�C*��W���/ֈS��^�AI���ti?������q��\�>�P f�a�v�"���*�"n��5�ņל�}W���C������W�^�6.�1���vJ{ �'�Ѩ��8����{�6�q6�2�Ul��;�Y��سr7��A#=z�u����9=n|�>d����)�����1��g�D�cyG���5�lK2������m%��E�sXWIր�s���=d���i%�u_dP��b9���yۣ�~��2hZ�-*0xb,u��6�k��Y�l����.XJ�4eP�=�=z�`/��/ʌB��E%�0�d�_IF���G$����"�}���ON�I��':�4-��<�I�-P9&����:H6^��y��a`<����,X��J�S���k��^�>jp�	ف
��L0�;|�;�oЩp�&=�:�c;�z)�@t�C����#{6�#���1���q�|a ���4n����(�{$�oI�'g� /�0�Ӟ����fr���T��T,��������h�~|��eQ��q��:���ݷ��R�J�*�T�*U�T�R�J�*U~LD�v9�d�/�"�>[�Y~Ď� �ZK� nVr����P̌᪆-3G�$ǈ����'gg��z�.Q�b�WK��p����t=��������Y9��I�Bs�\z���Y���3��岇�|�[���}�^��5��^}��D�F��M#x�!�믾��?��pv��X4D���;9�?��?�����2=�v�"����vf�T�*ӑ�0��0Օ�X{��&>Es�I�mA�w�/`o.]:����6-R�|z��C�ۑy�
�6�'p�����g��'�1�q6�c�" ���5��14�
=�E+��t��F�ox�"�����Ӌ$X�m������!|P���%jc+� ���{�x�g�⍣t���S?pD�Dw�1���Hzǰ���A�+�9]G�SF���!�ˉ�HWM��q9���[S}(X��+u4��}�X@�H$�Ӭ+`�^d%`�u2A'� y�G2��#3�l��l�M@BTG�8�j���[T#�i���^WW,�w�1�Φ�6��Iy�痓6�8f�}�ԓ��w�{��WN�P��t��OK�ڌ:,J���f=͎ @�C���:>��`���G��w�Niͽ0:�<Q�-
�6�I����9*H�P9�i�Ǿ���y$c�\.�~<�z�ى��=G����ӽ̦;0�~�Hgb����q���q]�.���Ȳ
쨅8^�=}?O.��]G��ZN�B�!Ztu��+��L��{FU[T��>S�۫�v�����S����=�	��aʠ�R�a�{�wd���ˇñ\�|aI��b��=CiTo\nMN�Ed5qzD�Jvs�ȑޏu(���� ��)��%�[ ��B�1W��ܬ+��n`d��g0���E����ٷ��p�Ͻ<����գ\v������:���/_g]�Êm�2Q����D���~�3�����,�����&ᤳ��/�v���yc�'/�k���r�u�.��A��	(5�4�C��a^�{�x��Cp�~����֧�sw5���N�:8:�E�w��r�i�8�B^y:�:P�G{h��yq��ݯz�Pɯ��������&�����]"�� `��l�Y���R����z]G@�a�
��/��4�T�R��%��J�*U�T�R�J�Lb�&�5�I�}� ಉ�4���Mi��ƣl�1V�{�c(�)��m�-� 98���z1�F��`#R"#�3�6Eps�b�+F�3n�xK{�r�0A�3 p5�|��?��ԧ੧�����!��874���E�;8=����?�٤�\�ؖo�C ?=��`b2�����n��*(�>�/�h���"�=>�����{���ΐ"<�z|ʠQ�b@R���l��@�l�cz��FJC�����	݃�g��"R��z�:E�I�����Q�!�jRݮR��'>�,<�«��3k`g��X�/{���hg��jd�,��l�p$�D��oӷ�^�MG�6�{��;ƀ�y�	�"���]��>P��:���%�����4�4J^YA$�DO)08ʛ�H�SELf��u�y�C�0�җu�w��t����8�@�m�
9�2�녾�����֚.C#�IC`�9�3��m�jC� $џ�h����|�q�ĐAiZ���*ۦuT��SE�>q`7Z�y���i
P� ߈��i��Dz��u��Π�=°�� }��
�E
���>���F��
(Ė{����-Wpx�!���N<{��!r�9�{��@��G��Y�5����(J���z�H
	�PO���
�	���Fǣ���S���g��`�Ύ��|����L���"� \
��@��M�`��
0�Jt+��&���=ژe��F#3�����=Ѡ�3���y�[s�ߍ�?�ҥbҒ��ѩ�"��q&�U���U��Ϧv�PF�bVP(�-:Հ�! �	�WpN�?�:��59�)e�����m���q)�j���y{���^�����۪��`��}l(_�hv��=�֯ŸY�� �.�5�_t�ީ�;;l�>"2ٛ����K
A֩��1�9r��8�C�t��2�V���.�s�/�O���������[����p����}!�Q��ș��O��:y:E���D���gY��
�n����hs�dP�{�ܣg�<���@E���STyr����g7<##����9|�
<��HW���_N�����;�΍w`�'��{o�Ž�E������q�'Gr�q�������Єg*����Pg�9��cf q@��_�M$�	�3�����)�8�AT�#��DQ�
�>�s[�Ϛ ��U�˄�@�*U�T��Hu �R�J�*U�T�R�/�jH�����~�.�����+���c�Tw��9�Le�9���SpZA���&1���38;>�g@���/]b�����x2:; 9
�I�(�g�(���n�x��������߆_��_�{��׳Ѭq���@ӗ߽w�������/� �R�����?�;wn���@��@?�/����w���z��dw����?�?���޿���r��n��t�3���{��{�9F�u���B��B׫��b�K'P�g�K�}�6�{l�"]��V�
���������S�L�t]���ܹ}vwwa�XP$�~�}g����{~��~>��?M�z��RL��b0�e��W�7�*6adx���������M�u;zvS��y�_�Akr;?d%F��� �� wR5�,!�홦y���@ϑ�~/W*ٽ�A`�|���']��>����
X��m{i.u��ehZy����3�+�o[�8�#���mZT���Qwɉ���e^��~R�!8����FF��`�C֏Iˠ�ԕ�ht/��*�s����4	��Q��jg��$�AC�#-�r�3M���P_�x����P�
�8CU��3wTE����C�GF zoo��sz�����^������;6d
y���H/XQJG cR�` ���й(m��[Õ(]kS�#�:"�������`:e'�:o����B�Y ��o��E0�E����]ҭ�$}N����>�M��SJi��ؐ�mJ�f>`�וS �B��{��$'*uѱ
�,��^��!�l:���xy����`�ޚ�Ȣ@�>G���ܱIL?藁>-Ĝ�����~W:P��zQ��{߆'?���pj�kꬖu=G��C&����o��CuK���g$U��Y+��m*�����������I�Y�y�A���91�7�o0�/�'78o�zQW�>��Vh�\̬Q��C��������>
�-w�����~�vml�����=���rR�<-��<��uNx�����y]�mrDJ����˒�et6R������*�����A�nq��W���NV1)fLӂ{�ᜭV�g�oY�3�c���.�c��9;��N$)@�r��}#�����i����6H��Q�:�6r�q�B:S��2:2�Ou��M\v�{HVL���A���2@نh�A棨>�.ڻ���U��*U�T�hIu �R�J�*U�T�R�ovB�2ͪ^B[��}���Y�-���(�m���U�Z5`s���AE��Qx�)�/|�7^��܀��"oy��h�{QC�QsG��<�=���"�����=������;�5|�'�$��{���j!�^~����|�_��1:4��-V�������8�r�a�?܇�_��3k����W��T�W��%���|	~�����"P����6�O�R};x�7`>?�)=�5�6�Ӄf'7ûҤI{���N�N��������]ސJ���۰��o��*���r��� �y��W�0���/���.E��L�]��ݙMa��{��8�>�rHop�$� �.�H�MF��갭�W�q��7vP#���L�?h�7�-F�]������{�=�����f��4�s��݁�W�2�#��(��`-塧贞 �U�:�@y��-L�=��r�{�5�
�xg�E?�Y/P�G���ab���:� ���i}9��� �� ò�_G��|��` ۄ�7�.��mzf�3�Hv�Q��$PQi�s��1/������4(�.28��G`:���q����?:�G,(d��9�020x$@#�!!
���=�$ �Őu�so���N[fB��/` 9|>��(��´��ڤyźk2�(���[L��i�Mg3j�
A�a$&]��n��	�|�i��ڄsQ�GG�E.�Â�~�N&<
`с:��s��x��-1p*t��6��4��]��=+dEix-pU�"�ΊS�	��B�y�x��-c�F�O���N�ײ����r��]�w�^Oc�u���ȫN� ��{1�C�o����NDYP]Q��e�/���|��/���k,4K0��HQǑ@���ol����h|ѣNw�<�����/���+1�.fǞ��y��\�U���κOd���t迨+�L�X&3Ԡnt���r�N�Q1/��q��f�Z�s�$a_�(Y"�~)fyyntֆ�ճ�`��B���SFЛ�E��j�V˴�[:������$'7u�G��s�G(�vq8(}���|���3!�ϸ�\��.�1B:��M�x�Y���;��QL]5_������o��3q�kh~�N�|.f 9%7\�ΨA�0�xM�î��SR���x�[��9gg{r�k�AƋ[s�1�%��������L���|�����>I' S?�:��k���Lƪ)�0XPU�T�R��\�@�*U�T�R�J�*��*8��F�
BC��|��=@�(��eԔ�I�P���H��݌,I]��#�Rh�^�d�LZ�����L}�@^����bzV��5��!���(.��ߗ�8�{�j?|�e�o��߅ݽ=��م���V��>9>&�I�85j��,:�h��p������u��y'Ӧ�i5�bk�_1��W��/�׿�eػ~�����s��s�Q����{���D7�;G�Jt����gggp��1N�]Ȩ����	d�@$���ar���h��N�`2��>�'��/�K��󿷞�ez�������
�ԫj�<J��Q���f?���~(�/��������3.o�)����jh7 �9���1��}t��9���hw=����0�¿�����?{{Y	�l�w���~�3���/=D`,1u�-	�����K_��pzr
w�݁�d�'����s�3D�yYz�#�#�'�T�7p��u�Ik�C��4?W�����>,	4aC���|���S,���<_�&�P��q]b䵋��_�M�������Fx�j��c��G}ٶ+��� ϑ��������\��ܼy����x�Q��NK`�)�_�~�6�w煽,��1ۙ�C�i����^G&�W^y��D�K\��'�G��S_"hѳ�j@v�w0��tF�Sg��4��X�N�Y�-Կ��&~�.����" �3:&�3@����N؁��h�:�
�t�d�2�~E4ɑ$�S����q)ON�jEN �+q�|W�3P�\<w�0Sp;iM5^�8*������`ѧxoG��=��)�m�A/l�×/�/�����7n��N�����ӭQ���	P5F,"�K]���k�H�Y*z=S8�5~�3K�{�lR���� ܇|HT�Bе�.d���� 8L���lP����{e���9 �xm ��]���~΀,�X�S�A�(�`N�D��ܨ��������Ђ�i��K�3�/��s,ߜ�8������R��;h<+'g4oNy�;��hK?K���?��'���tߎ(㞅u�kAӱ���QCǷ�2��D��Xw�
�d��������;��!��3_>��u��p��LB@<�GGz�o����W���M����<�L�3�[t�e��������ڊ�S.�4:^�*+�r-�u���Rp��iw�a#�|��H��B4�7���R�Kw����2����eӽ�ȃ�����\f��[)f�8<���'���LG��1U�T�R��\�@�*U�T�R�J�*�Ķ�>bl�F��?�/1@�
/,r��V��V�"�������zj���el�ݗAOs����0pR\�J�
f`���X���"
�gZO5�"�N�B�t�w4ctQ���''��ݻw��P7�ɑ��D;��h�#��~�A�j��0D�С��A���V��VDw* Ah����`����ޑD9�����1
(+�Y��ү��������h�F��R�V�@��2
�bt:t�c�l_��F��N�#��i�Y�cA[A��� ޥ���~5H_D�|��&������v/<��ڳR��'�P�24�"��k�@�c�|�\�Ωs��p$�H;�[�J��O?��f3�v�:��NhZ+Hm�ꫯ�׿�5�{��LՈc��������2��s��Q�����W�W�ҥ�Һ<!�?qPJ���W���'�|�X70e ��۷n�������l� �o2_0��@� �9 (Ҧ���[C�lΫE	6v��~�k�5:���u!�C�*|�ij�#W����<��#���/�S9�8��i��S��a����������ksn�3���������S*��oMà:r��D�����$�����SiN�#��n�����O	XA�2EF�� ���ru�;�#�7�d��ϡ�4=�O���,co������~7@^�H��IMQ���>|h��ԟ���5�����Ld�h�L#�,18��]�@���Lk��}�Ŕ3q�h�c��}�l��7�x��9ڠ#��͸k� o�y�R-dx���?O��!�P_�0r(�6}
�'�b�)�C ���D۳����Z�R���ֶ�:�8w��:v���ʎR�xf��>E֋Ľ�@Tv�A&��ҷ�������8����qn�"�َr�'������(��ZP7xK��OPjǺl�g�4��ns��>�9א8UQ3�~���3
P��f�|-k��s��3�t�w�����j�Q��q?�Ը�yAfǄh�y}�8)p�y-���f)�$�WD'˕�w��gcom�7~��Z\�Z幚�>؝�����C�5Z;ֆ 2�S���~'�/�i����د�����@��������CG���O|<�a�\�F��{��+[��y�<���"����D�ۜ0 ���7��~Ni��>7G��|�:v�@�Gl����!:��I�ղ���@��Z'��t�����rF���-�T>=��X�-Z:!濍@�Đ��J�*U�|�: T�R�J�*U�T��@�"����$���cJt�oc!?68h���N �l���2e��>�9Z��D��P�t�����Ht�.��'Fug-j�Uc�RQ�D �AA� rh�7p�'E�  � z/�8�`�?E���/�`�!,%rMk�D�I�ϫюi�	#*u��\�DU��ra:��{��|�1U�IL9]hT�S䆍��#�4J+�ꖌ���<��z�q�m�g�����,ҵ�-G-���S�H��0��٠�L��!5���M�����@��ޫ��{f�=%��~
�Y�?)l�z��i �b4ӍF(�wD)N��j��#�������i��]�X���D�N4�]+�*���ro���e`��F4�}�9NTf���a�2E�Ogp��U��Ǯ��[w�,������}�=b���م�\�w޽I�sＬ�FRtpzzʑ�Q��y�p�S^��i�Ũվ�
mc��R $ñҺb?P����o�O��jOt ��G��,�#���@@4�1�S{888��1{A`��Ã}�r�J�~L�K�A���ˁ�B
`
e:�qZ�vB��#Y'���sĿ�o�<�ԓĈ⛖�U��^~�Er:��|q$�4�DPrj�3bz������A� 2gzMA�],)�fB,$���8tx�~wRf�	9�pJ���g�'z.���l�ԅ��V��@Ht��h��|��p������S#�������`��=�P-�ʑߍ�1�{��LXȮж�� #T;�7������y�M��T?l������Ou�E�nБ�_�&&�s��2V���R�e�v�rE�m����.��mZCӝ8;9�94Kk�z�Oܷ<�-�������A�czt�RG��=Ʈ�z���х�Q �+���St�:x�!������f�)9��K�`7���.��駞&��7^S�P����ɟ��}�kvf�r�(���~,+V�S={���0p$u��%*[^�#Q8:�����2Z��::=;�
d� _}./�5�K(�^Ͽ��30=K:���v��\R ��� ty��5��f���~w�-�䠓._�����a��@9ɘ��ۭΒ�o�9S�>�&3r������`9A�ך�����^K�u�)�ĉ���p���Q@���جL�R<3�����{c��̥�B�>S8h� �6����	���q#�;8=���B!Z�5���9!:b�q�J�*U�|��: T�R�J�*U�T���
G@ƨ�� �j���8 1��f���r�Ս�f�ʆ������RҶ�V`���(���G�E~�B�&%.�-����C�эs}���2|ކ�6���S<>�	}>�$����$O3�#(��}hg#'	t7�[@{2V�〷��䒊!p'b����f�3�/�9Ӑ�m�܁���ɑe
���S�4�s�f�-9iE�h�$����̟ FN�2�8��Q�:�����h�� ����@���|F)d�9(lsD���q�[�[���8Cv�ޟ�$
�Is<0(L�6��a�����۷ᅗ^�{w��l�ݝ��v����7ɩd�r�6b�ǵ��w��7�|�@��jA�ir�]C��3z?�h�?::&���͓ܻwW�Lh�aZ���S��_&����@���}���j���[p'Օr ���uȑ����.���\W	�A�E���o"~������wݗcX[�<��|�Ѿ�L8u��]i��]\�|޽�.E�S�=R
�RO���DĦ�Sߢ� 3�����j!0w��-�K��F]o������k׈��,ݏN
��[�	�ł����L��v�ܽ{9����+� �'z�S���S�`ۆs�7� B�"��B���R\E��d.4y=E������d0�,f[��ڟ�N�Fր�Ԯ��M���4��$���OOa9���O��@��Q��qX	�	���;�P=p^���]�qA��
��{pr|Fm���LW3�;����
�:�q�p�w��G�Q�9��.i�m���'��u�ۧǺRsQg����QK��_��]�e}�Z�m��}= ����Cx��i. c�K/�{iN~�?A���u�!�=/��9X=�����)�#\{�{�H�����1lB��Bܲ���1��J��N	�b�P����v��;#�����w�t��iiM��Id.y>���*A�{r�Ӣ9H�2�y>�Z���L���%�����?ZG��(D0}� 1��V��	v��l�Տv�њDݕ�n�"J&����`!{��V�p�qlE�ϑ�,�}��H��	hp찮98��yʀj=���������tހh��W���il���EL��u�I�X��iC��f���V?ե����^Ƞ��-���>�\�^��e�د�����<`� {�y,�C��m��H��l����4x���m�y]�� s:�qr�	f�6C�)S�Q(�b�T�R��GL�@�*U�T�R�J�*�I��|��.��Hg9�7Y�Q�j�2Jk����P��}s���zoA�<�&�g.��p�� ?��HW} Bu�z�yg'ZL��L��� �'>�I�z�E�a4یrXO��x{�շ��{��{2m8�v�r{1
�f� 3���li�<����EV��p��̈́jd�Xkdl�x���"��r�]��;J'����3�/`!��M;��^�Q� ӞBအ���b��F
��Ecec�Ji���X�߳)��ÀO�E�o*k��r�ϖ����kE���\��jAU+���B���# Y����CƔK��}����7ߤ���d�;3���}���"����:�����	�y띛��'�-�`ow
��+�Z�E@'�����p�]��� -?����˩�=�����s�"g��ܹ��^x�Eƃ:�xî\�G''DS��g�S��EP��t.s��P')*8�R���0�f��ƈ}'s_B�)o�qXbr�p8[EN��V�t4^�	�Bpe*ή^��\{��O��c���9�-�I��Q����ډ���1�$ũ�ɣ���Za�3�Q��(�u� 3�N(��,c��N}��+i��!co�N��ӿSx�韀'�yv�����3��L��N���b��(8��=��Qt$��8� 6����#�<?=f��q:JA���|�J���%HI�?|�a�?�~rx���47�[�����٫I��N1Ճ�D���r97]Ok���%�&�mj&-����}�������ψ�A�g?󳴆0�{2�Q;&�N_��׈Ee�݅�dF�+H?�i
?�H���5�c��f���H7{uP�:��[c���ǎ%pd��F=;ԕ8����Y�x�y\%K��B�~�g�у{�\���X������i>�ώ�9ť9prr!鳝t����{�r$1�>�qv�q��	x��'{F`�J�5=t鰚�CG ��xuI�^S��tR�\�Ug��_�7��I� ,���d�p�<��p7`kZ����۞��o̂Ya���iOA'���S:�d6%t�住�Z`������{J�$o�|���Y [�A�C�/"�K ��Vx�!����n� ina���8��#IT��?�Yg��}�zvr�泆�NM��q��WƄ�e;�l��%���D����R����3[
�͉�/+����A6���1Ph�)���O��:z�"��2�^�ka�/���)�^.��X�Vبk��D���o7��H6�d.�!�I/�� Y)�����h�7�yB� �R�J���T�*U�T�R�J�*UT�<�b*��b���!{l(�fl�@
#��3� �J�:[�МelĖ R�\�j T�xl��k�6�F5�5/��Q��(}�;߂�yO R�[	�826�y�hUg��v�č$�`�0P'�a>T5@�h ��O���}A3 ,e�;���چu��B�
`��!��+М��[e��.I���Pj�_��9�S���,m���E׷Eڿ_0�<��m`Z���
o��7�w\�n��������XT�,e��eѣ����吮#�{�����홧���+�ק�z�	���MX,��&�أ�����z��g?7߾Ak�S�~
~���=����(����+p��u��u�\-������.\O�=����o|s�����W`2����	\z��U ����Q�ϻ����`֭���ܿs�.|�o�%���q��҉y���g���/2wh.��@[BU�����ԦF��95�-hZx�?���S谁 s���D�Q��HL�#�f�%,�:��-�?�w���, �����[o����`%�/:`T��K���^�vW�"���B�Ge0m&D�O��z;�(W�����RIL�;(�e���6���hK��8��> PU�b�"�g�p��b �����?8Ls��(dQ�Ѡ7G%JY�����,A�4����TR0� �%�1:Q<��'`���Rp`g����3zOGiY�b�#3�	�
��\f�	�Wr��=FF�*�pf��A�G�e�5ԩ�O���/���.\vi���[�6'���i���6����Rv���Ӟ�)Q0-�Б3�)�2�=�n)�9�N^.V�t/u��|P�|T�uT=oMPp6Gn�r�3LMD��˜,�?r���`�@1}	S���;�t��Tvo<�ߏ�N��	�"/+�$��|�� ���}�u��p�G#�;�����K`��5��]c)�r�YC��Gc�W@>p�5�?��j\�,�����}Yv��b�w���(K,�4;��/�]2���:v��I�����U��g�v��g���~Ӹ򬎩tb�!�=���������Rzs�a�AG1�nE��V��o� L6�,���/4]>�]�@�_fPpEE�c��������#��I����ګR�J�*?FR �T�R�J�*U�Ty %"�������AX��E�(��+� Jp���b (8\pK� �]�����r��0Z4_ p-��7�"���{`�fP�>����u�~� �� ?���1j��4n�/�㼢^�����g�^$#������������̊�;��[G�K�׾3s�.�'���~��osF(�.�H�P�f#�F!i�'G�H�V�5�|��&z�m�Ƒ��?
�����Y�g���^����Xk~\���A���^A�2Bӌ@	�8����޽y^x��0�݅ý=x��g��×�F�
擿r�*��h�ǈ=C���S936�ˎ��oÛo�I9����"�_}�U��G��ν;�k��kppp�GGd�o<�.����㏑�H{�<���`:���K��?xNO��'��4(,�:���yx��7���O�Q7?P�v��,�X�;��9�q��O���l<<����A)6�3����f������|�'�H��t��q# �r��! )�W�C�\�m��d]A@I��?8؇�ׯ�[o�E��x��w�0��v��ux��#^�\���xp�dgǧp��=x��W�(�=L�L /�-)%����.�t�{�gا��P�|d�l�^�E|7$��L��Q� ��|�1'�0���+�(
�X��>�!�L��K�f�|n�;��L���
A �cF��s;Gږ���"��+4�<!@, *���N����A����.P*�1p<�5%XT�w�J�A�G�
0*j]�o�&����@z^P�W���W�9I S�k�f8�(�=�mؑ��䄾GdM��r�:��3�P6`� 08�|P�����;OHQ����;f��[���H�X�+bW9�f�/����4H2�@�"w���[�����rfNQݼ�e�,K��?\.	��o��X?�d��������QΝ���A9������Xۚ��wݟ��ź��&��{�e�����ŕ����<�;md��ֽp,�k��tPq�"`�Vi�8����-��6���4��r_�#JO�?Z>����Y�rʘt��{q8�r>BC���<]��<ݻX���
.�[�C
���������V�w���m>Vn~��]п/��#�J�*U���Ku �R�J�*U�T�R�5�G�$�R�� �1�e ]�Fym`�xf+$Eɋ��J� f �g�.�K��#���a�aTA	R �SdS^jה��
�1�s1R4|Ր��z�)	�.�.5f�l�"�:Sk����ț�c�`Ȇ���Ж���N�M�}�;~v�]P)�X*!���k ���B
4����b�v#��n�6EΗ@�&@fx4~��D�����M���ѓhe�798l��m)#GxF�?�1##x�Qol�`k�m�8*.�DŲ-R�ߦ�o�s���www`�\@��oɁ �H�(�-�����������ݻp|rL@�O�Գp�w��3�G�g
�ӳS�/�0��ཛ����=x��'��1���4�Q��or^yl�r��u�e�6*V!s	� ?/�r�ФFz�NJC���/l�z�R� Er
h8���cf�P`��*dV �e�^��=96����:��{�'��I;��r�`W�A�����;���V���x,�#Б�L��T�!]ܝ�R��r:�<���{.���� vt� 
랣iU׸(��xD'�	S�C޳�N���Xl0$Յ����8�Q���W�\���4�[���e���6�j��i�$Gd��k���?��ڠt�����SX��8��?�().��W�X��GJC�ֻI1�2�y�l��^+����}�>���w��Ō��5�����d�oQ�����L�ڧ��.��1j鼂�"����U�{�	,���i��t�t2c
~q"̩t$D�~;��|�(u��(qW�c}�]��9E��iO�;m��S�0~��@u?�">w ���w�gK�lwS#�?���� �K��^�Ct��l��]X-0m�B��4��Vˎ����d�aJ��9pj&qִs�dq�$F�"W�٫�]�K^C�����~P3�mtD<�x'H�G������Y���?���z]{+���L�X�d�� �~��,�2g�_=�:���Ƛ[���:J�ġ7�v`���3���3+��_��(独Cu���V0?����v��G��4�wR�����Q�(r*p�BQD�`78k� U�T��Q�� P�J�*U�T�R�ʃ,�j��k��Q��U��G�ce�b,>2��zdV*l@��Q�D�cQ�_���]��5a-0@]�`��cc�bV�
��2-G�J��<2:v0�fW'�om�����(g24F��o��=[�߸_J�I�W�o,�~���	5p��9K��:L��PD�Q��P��\�����h�+��e�\O�LUc.Ϗ �5����%e�8�_�o�<��"����޹�ٱSCj�m��&plE��qF��2ݶ��(0�(�k��i�57�΋����?w��a������)ܻw���h{���N9a7?;�<�278=<r������}X���������g>�4<�����˕f���D����|�-x�'>A� �v�L�	�H�,"JC{��q=�bX��Š/vExc�uG`�[ ]/���WQ0
�`� |���� ?��s?���s8����G��K�w�j4j�jL1��b�?�GփɄ�fyX��i��*D��@H�Q��}?i�� �18vY�se�X{�Os�%|]�:��B]<�H�u�pi7`:S���L��h�'�g����V�=-/�#��u�fC 'L��|@���u-bJ���A��A�e����	�
�LRz`gKu��%�8�m��AP�p�9�C����`{��3r�s��q�_*u�����zA��&�U��w?�� ��=����Ͻ���=��83E�^�.�WKXMi��a��t:���ֿI���sz���=����O�\Wl��z6˺��4�e�� ��H�RzV�u��?�S\���3;;��
?��茓��v���~���I�s+�r�U��Oo����l� nߺKW�?�8<��3�ܷ��Œt0����o�x��=�����=}� 3�ǉme}�}�@�b���V��E���d���Z=�]��sw��e���H�����B�z�{�Xօ��_��Bŗg"F�Q!C;LIz�Go�ę���H�����wv��D���{y�q?ù��ц;�|�S�[3��������}�{��ɴ/E���L�.��8;[��V�L�Mzav��e:r��R�J�*=� U�T�R�J�*U�<�B���/������	2�� 
���L���(�5rF&Ju�UF
DL�9���l"���U֯�U��\�$5b�4f�0j���Y)����T��ȔJT�Ls��" ���0C�olX�~���!@�&	�T�0��)�R<`�.��R���À
:��(I ��<4��0*3�1S۶֯����97�6���H�m�A�W��}��ݶ��l������&F$0\��t]��{�q�t$û�>!�3 �2���������:i=G���҂j���Z��������×�V���&��\�L��n[�'�y��
����2�M�$޳Z�,�{0��Rux֢�h���S��OgF~g�Kר�r���h�}�M�Xb^`]d<L��z��O�8��z����My��^5؃��Ǚ�ϧ��z#�|+�)�g@8��j��T�ԭ��uN��Y� ;���躀�@A���|��|������W@E�r��W��@�cr<�v�3���E	o����]��vZ 
|J��~�s�D� �yB���z�Ynq�/qxrEJ��w�Js��' H�)υ(�U��ɆG�7�Ж_'�ٻ</�_<�;���v�m���>m��F�Vt?���fM6].�����Ò�c��s���i��N �b�m�_��p�;/���/{�#Ȯ��ϡ��V�^�۝�#��ՊY�%�$
+Q�v�����5;�ޫ$27 ��ռMve���\�L%
.��n���Qz�'���+�։֏��:ϸQ�ޯ���P��ZP�S���'k��9q��߃���/��=�1x��mD�z>#���x�C��;� q[���by�������-���n�B]��=9(���E���3T̿�UI��BK}G��{�{L�L�Ec��s� 9�;+�u3�?f�R=��^G��`�#��qt����/W�@�#��rn��� �Q@I���c���Oӕ9=��Xvk�s1/��U�h�e@�Ye��f��[+����W�R��GQ�@�*U�T�R�J�*�D��	�E5����/�7���\�-�
�e����@6~��t�C,R�`�>��oM�ǝˆ�����5z@��N��j�s�S�(�%ϗF�8苵�E��=��b��`�!S�eê���s�^UV���w�u�ܱ0 �`��9q��$�q��>�V�������Fi�ddZ\3~^���g��?/r���-+����a����~
*Pn㐦G]���#��A@Ac�֊� �]������D�|���䩨�+��D�e�����F���������FVLߋ�����p3Zm�G���d:�2BOѲ|3ؠੂ'����6��n�-;)�j8g4�"�U5!`��0��}�A*� �P1��@SO���f���E���<�i����(�ӿ>�`G)~�ۚ��z�|3`�� N�#ߢ���Lђօ�+�P�H"��U�Gq�uP��əE�>b�cC��2X�:�q�����!���J�{D�ǂK�^u;_�-9��)"n	T
�W��U��~�h�C�l^Xxĉ�u�}S��-N?�	����s ���5��Z7�Z�2r�tʰ�P �}�������P��6��¨��p�zQ����urL�֝'c ������p����݁��]��IQp-t� ��n!�%ڦ@�Q��V�ј�h�t�Z;أ��"1}�9M����쀀���	4���( )k������6R���s5����	����h�
+UCk�'v���X!}<:!J�od`�5���3��v)���X���f��PV:��i�Q���@g��yg���J���|�R��i�([%pϓ���"��+��91 ���I}+}��i��=3��3�@�#<ٞ�{�"�gp~�!�_�g����N=�[ue�G��3~>��1룼ɛs��ϊ��ы�R��iGeZ_= �T�R�#(��J�*U�T�R�J�P�	�;g�-j���`CQ�o�P���")�s�K@�ڻ3�_F�	�UF���F���\b,L_��@'/ˆA+�^/1p�0���z΀nkJi_�Cӛ�/��_3p�1R�.�����	������A˷�I�����(�(�+Z	 x1��Ϲ<�*s �;^�2u�a7G��WA����-��1��L�?�\_�Ľ�i[ٛ���?�
G��O��z�gX?�!@磚v��?-ی�2'�h� d��<'��m��9���An�2��;FO�O��(/#S�O����3�vt@��"�Ry����C�)��R:����ǹ�e���V�41�s�b��kj9'�:02��Jg�2+�m��V �K�7�/�t�h�C����\�b�s��\fp���|��/�[�W��H^4������ 0{ &~�HSJ1���Ⱥ�;����(����WHwH��QDn��Y/�F�c� ʣ���2!���ӻ{�1r�s3��+�4}¤�v'�/�.�>h�q)�����w��/���܆P%�]�;��t����1�O)2[�V����"���8�)�4�#�����Hm�MI����` X��s�P���>��V���v�| p۵m���>�Tϋ��.ҹ��S:uԴ��� �1��������3r�jf{���n��W_�e�O��犃�C��v��7�y�C,�3t8;[���-���ɢ1 G��2�������1 ;�4#ݹMkdr�ZoZI+�oZG=����炱KC^N�h�-\ ���1
)p�88<�+�/��BڧPUQ����$]�l#�d���C��AƑ���s1�1@~�O���ڌ�ƴ1����[{��R�egcfߎ����>J?oy�x-�s�T;����7r\�m�u]���o	q�R�d������(F�'�G[q0p.�C݋��B<��ݒ�8z)?�`ӏP�Z����F���:7���|�묬#�]�2IXS�}m��&h���D�R�J�*� U�T�R�J�*U�<Ȣ��.���`�D��8���O�cӫ~�ϔF/�'��6[��202?�A0�y�Ǣʆ���oC�=����vXq�����0���1Z�z~<�W�+F#sd�$��T�%�������g�F��X��R���C���Y=�����`�J@<�92X����YoE�X�p_*��X]�ka�.��:U��0:������{���͝Ϭ�+�6n���]�ޞ+�j����_ɝ\TA�Y��^�R�r��F� �h�`�@��
��yʐ#���(�4Vh�G&�<,�Z��G@A]���H��tF���޹����Ƶ�v�,���h���:�C�q �;>=��l���w��{�Ӌ���(}�������k�Q֔�c��E�:U��=G��zRg�<��3Ĳ��m޻<4BG����(��pC S6 �ш#�Fn�y&m{j#�=8s��VK����t|�)��3�*�`���;s|`��N����+���Y��N#�z]�.�;��ԁi�� �3�M-�rփܙ��(4��A�5P�k:�����@fP0�Hu�T�c�}����u�@��e�R$i��R]ʠ(���q�(�}�/ډ:���h~�<)�D]����(�X��F:���X�U���>�_G�M�Z4�-�o~��?��{,����ru-[$��3@��h��H�}m�98v4y��X$�V5L��۝Ml�'�p����n'=KQ�I�.��,GXu5�#�Q�u5�&��\-��zF}&��0l��0���|/�#�k���F�$2��|�h�T��(.z�	�Y<���u�/��}���|�&��Ҟ3?>��xvvF��1��)�;�m�+��`���Y�8�����<*N7�a�5J�Ŋv{���=eϮ� ��p&}�N�����	��W'�\�A��FEϭ��q0~�Q�X"�s�s�B��:�^�~���e�{��a�=��ШC��k���;���? <��s�Z�u/8%򛭷S��a�A'��4;���/��sx?(�U��e<���7G�*U�Ty�: T�R�J�*U�T��@�
�	�����j�ʑ3b�*�r,b_:���,+r(N�c6?f|^��z̿����_��ʎL��v���f���R3��3�����f���r���6�_�L�{5D�
�\�}(�)+A�}cF_enpVk�GV�}��Q�2(A�e�h��F�����V�k���ǣ�m4���m��X6E��#�7��?�.w7m���{��X��(�z��d0	��+��]v�*�x���<�u�y�EX-���Q�?E�S�9W,�K�W1�[;w�m&p6_��lN�c������������ �%\�z{�J�C@ j���M4�#H�;��0O?c�LQ�Zv\�t)��Bp<(����E/1��d@)��S�#�A��(�i(`���h�`�Euv�vɚѷGmk/l��"b=����#:�`i8
_�8Y�Q�T�A�ۣ}F| e}@�Qj+'��V(��B�U �1ۆ�lN�(T�E�w�0@�����$1��p��yhB�k��%Mq���#9B03;�5���F����&���*��}�,(�����M���Q�=��y�N-� �s��4�[� �|��t i�ս��@}� ��y�n��OX�|��`r*p#ȟ���u�w�����ipS.�"9O�o���i߁��}��@s�1�Z{@�CVG!�Η�F��1F߻#�9|TG=UW9Y�4Od� P霾H�qt� �]Uy{������s�xmDv�L&�K0�-���6���7�~.]�D�Pd]��"�^�Ĳ"5*Y�c��~���[�Wu^�]2���Ⱥp/�3�����7�q%rjӝ �],�K�Co��KA� 	�:w8�ku
ѯyM�3Pcֶr=�ڈ��3dX/`���~�<W��\U﹌��a�N����I����4=���ܨk0�y(��w��U�I��*�Q����[+�м:@�c��چ�[�	k�����DR� ��Y%*O>�f���ֆ�#�+�2����8���}7vhҾuYig���]K>;���lT� �z��T�R�ʏ�T�*U�T�R�J�*UP!�˨�A�t��f�E�3�ό���>�b.����m�����8�7fDm`�F����l�ʆ�l�BӲRDG1�g._#ۙn,Wha��Քv��D�%���xs�c\�#�LX�F;Bv pe�纒y�4$����1)���]10�� �U64
�Q�GjX,��ύ�[Iѯ�a}�ܚq4?7��nz��g|�|n��OD��8�i�]��}��k9G˛����]�#� F��A�P��<���yܳ��Y@��s�^{����-��GeG@� T�A����W��5��<>>��F0��_�\�:�����g>?�쳰��G�#��\I���
Rٳ��-����:rBiag��Œޏ��
Y
(� �ݲ��|�uk$��& ����$֎�^�aD��B-�S���ޅ�?
�U��Rt>�sg�������� �5�x���G��@�>H�� 	��;eH��1n�^�I����Wp9^��� e+P���ė:��@�����G�7sY��Qpd�#� N� `<:\�<��`
  �i�s�i`�w����Θ_��{��y��1������)G�4�G�1�q���q2�iN���u���f?@:�4W{���{���+f�����UF��{���{��Cv��/k�q��w
N�!0V�*�3�Y�QWnUw��=��&eo.e�oه��c�����ޛۚ]�ak��s�}��{ݭ�54B�Q�nIH�  2��I
I*N!Lq�W%q�E(�R.�b�/���8�I�C�)18�� $�A3-!!�[SK������t�����ƽ�w�s�mD�x�{u�w���=����뷆�c2s��ʘ�D���E�8��S��A�����3�x��,or����I��q�	H�W{�y���'�q5��v���*��G8j`�@*zԓ�N7/m���k�/?�7y�e�-�Fa��<��o�]�&M�������ev��o֟�5FH������fgc��r�){$�Ce��	}vA��k�
e%�z�s��{�g�s��A:��A����p�s��Cy|�1]����;ܱ=��C?��̼-�T���RW��G�9�|�Z�����7���gC2ݷs^K$n������P9�5��'P��ꃁ��뻗-z��#���P�%�K'��N��=�·9k�/w�!��P6jԨQ� 5�F�5jԨQ�F�nA
�a0ų#֌
�RT���&-C��!�y�+uX�:#�F�}֩F�Nm�BQ�k+rd�[�3׾1p�X><j��|w
0�P+�n�ߕG�z�_� ���)G�S��@��N�ʒ2���k��lR[�� (�~I~vR�B.�J2�e|
@c�Ab�C��T9m�7���u�U�J���(
��MU��mQ��k֜\����):-�s���s-#l�w+Ϫ���� ��@�#�m&ё0�z��w�'	�a��eo��<�/�v���9��M^�f���!�� ���Sp�GK�t��G�?�ԧ`gx����?Om|����.�7�o�?���%yLc$X/�~�<�>��/�G�Љ����U/��̢���+ϒ��b�C�ۉ'+��I5�Ď��,	X ��B A$�����d�#9�����a("Z�w���/Fq�b��M��W+�_4�Ib(��L,�y�9]FKX�=���v��ެ�a�f�������	�ulD!��;x�N��a�$#L���	�^�t؆�׸��"��JG��ç.����fP����N�^�ꡈ����9������Aj����� �������,,U��I��"9`8U 8'֣�F^H��`Z��f`���ReNA���87@���A/k�K�fP�UÚ�������s����F��F�lM��x�ݏ�6��g��Z�����mh�a¸�Sߧ��������w���l��Tƀ���R_ w$�1z�.�x����E�q��A�*1�M����u���K��)��vc6<ѴQ�c�9T��n��pm��^G>G㡘�2+��j�T��?�����8�yb�<�,���i���b4�~�J�*{B�m����:|�ue���B�@�J���F���9��`g��iH��硲o�0������N�q�5 `�=�ϓ����S����RZ$[�%Ȅ,r/�*v=���"�4AFXC��Ŏ�|R���Hx�'#���5����i�}1h;���Ҧ���_:�-:���K=��4KW�XO۟V�Z&�~+����uG��7���ߨQ�F/0j �5jԨQ�F�ݪ�8�yu���A�Jz��1�U�yp��;u����xW�W�`�E��Q�-���`{� �����/_��Y�ha�E�HJ77�Ԕg�]v��b�V�b�C>�h��&�X������;��Ku�C��CR���e a5>�h�rU���<���c~ �+j�п��唊�R�nN��xb,}}��UE�Y<צ��mQ��F��T�;���,�j�`�~���m����o�I婔��|���Dtu f�LN� `|tt ׯ_��|��я~��>�5��=S�������_ƶ ���]f`�Q(��ի��)�)lޅÃ㡞CR\�⌀ԫ�^%�v����ptxȞ�r>��ư�ȟ���^֊�ӑ�|Ec�9���$�<0@�ks(�ñ�쉍���ҋp��1}o���5�n>T���hk8we(�Y]��^4�X���2�~��Ay�1_w�y��_����C;��h�1���Q� c�G|Hʞ"��`�4~���03��#^ɜv`�s:�[�C���#'tb���@i���u���X����ɼ,cR�|����A��P������ S��㩀�ؓ<KHvt�Wc� ���E��W�'��s��5���i���mo�����?� >���vMݠ`+�-9�lX��������o�s��eV��e�s��eg��`�����N�o�̆����$i��6�-ul�e��G���|X��a1�@`#>�1BFx�'��?'�(F�;�����Gf!�m�����ޛ��Zʶt�R6���?��pqr�B��{	��ȼ?-��Ȩ%��rX�P�ۏ5GI�6��,�g6�	�)@mq/XK<)�ie�qM&e;m�B��7���	�t��Vv��'��eN�c�r���/i��B�A�P��I���j�L���lS��a���<�3!2]��P#	w6�+�/���{ Ų���D���Ο��i6Ө2X�n�����>!Ȟ �����f	�w�G�-��y�����׃�+@���v}���!� �m(�΢���fN�����5j�薥f ШQ�F�5jԨ�-F�i�$�e�7T��SH��E���>�jO)W��~*E���J�Kɣr�݁�XŠ��j��'�&��$
bփ�!@QZ*���.�֊R0:�Uƕ(	ؓ�'n��埠��2�5�AE~�v�c�4�zOa��PE*+��1��fT�-c�����׳�5��.J�l
��&��s6R2����Sou��-����@�1���(���ORVmQG9������Y�]�y���q$�=ƣk��Ù�R/�z�N��г~��'���A������.z�s�u���ß����G>�}���/e������Ff��O}�S�. ��m�V���F���� w�_B�?����c_�� ʼ O#=���!c��#
 ��j��Zk�m'��@u�BW 7�K�>$W"�rz�ɵA���}%F:wF��d܀�o޼I�����B$�b��1���$�����k=�	�<'�G�p��Uxꩧ�K�S(��Q�r2YS{�8�a ���v�O' z�43}�{*s�#W�0b@���9�g�9�Bެ ;���3ϳ\�-5	������{�8r�pK"���(�:(��Q���[�  � �5�b@C���}��ºq��1TR!�V"���4C�r]|�&�Ll�e
X�@89�eR�7Y<Z��g1�4�{�Q=jS�69�M�U�{��m�|��|�1�k�9���u�p睷S
�A�9��㦽Z�$;0��z5��^2{N6.bC6��tB��%EB;��j���s1D����#�d%YW�H����q]�ҟ}��!� ���K�Ǟ�U\S봖3X6�m�ŸBC��8��r����j��c叶9��4��N�-zd	yek�H*݆} P��a9�&�s�u�*�7@\�f�1����v(F�����3�����'�q���&�ܔ2A�=��ׁR��:Vjjy����I�`��y9���&�[o����?��o�4�sZ{��h4Ȳ�����^di��~�A5���J��f�������B����H�BS�1VA��|ʝz���z~�sY*-_��Q�F��R� 5jԨQ�F�5�)�B��M)暆U�nR��%	j�7O�0����(F��*�+�ߩO��x��;Y�V�j�����
��� Wo�,�$����S��r�5��F5�`F)c��Da���U'�U*�(R�)��x�Q�j'�!A�t�(�N��ǲx�>�x�gū���HڪgΛ��1�  ����9?S�S�=0oM9Aa���vk��m<{V�_��-�l�\`�E_���
�8��9�y�A�B���|og^��W�������C�̞�"�~�E�F8��G��3��{ᮻ^��;����C�������� 㚒�@.�����C[����Pأ�ÿ�n k� hu%,ٳ}�6��V^�x���
ܓ�E.�h�����Eސ���# �޾���1����������)퀂Y�	İA�k'�����"ЌsF`"e�{��W����\!� ���0T�
�RX�����>{��Ŵ���O>��bZ���l���a�3���X�g��J���(R�d�b�ǺѬ |��s�"�����=6@`5�#�)<^I���6�!�c�=f<q��B 3P��m�$����`g�.����]�3F��vc���	%�� #�#B�H +w��>n����pR��	�����)�d�>�2� $�g�~����g����b�٩���.��|m�3���>�L���T<��M${.����j(赯��W��]�?�5����$�|���ׯQYׯ߀���am3@�Z�I6}��_����ʇb�������*S�m���I��;��8�H�\�xq��/���jg�/����P}�A�cZl�C���SfC��R'��,�R
��J��ˀ˱,XI��Y۶wn��ӧS��&T��{�?6>�H�Ӛ�;>Z���\�yP@ao� �-˝V'����g���ƶ�یx��[���|S>6�Trp�8�[����!�lب���b��b��*,K�:L׵k7%�̒���*�o6�e����ɭ�?���ut��[�MS��5�d�A�B�d=�� l��AԿ�������35jԨ���@�F�5jԨQ�F� ��!�DMգ �~.�{��T��Q>VU�U�i�# ?��>��iI��"+�
 �zg�I�W�朸��%u-����L���rmC�l!NW6VN�8��?�0�o'
V�POE���:OJ��P�j�� 
<�P�4�)9��f����ٴ�T�Y�qҴ~�w�K�VLOy�{O��	��O��2(�����&���p:Um�gy���6Q�\B�F�j�0�����4_}�e��s����{��h	.\���^tǝ2?����q ��=^R�~i��~�C����=���޻�._������@^�6I�vm�+���)�?����0��<�=�$I�ؼ�\ߚ��3=ũ@5�$_"嵞I� P=I�|j��п�ae#\]�Z��h����.��fd=��{'��f��x�"hMa�����4~(I�WӚC����	�n�0ﾙ ����M�� a	"�����p���Q �C��os�!��S��=��@`�z��-�r������Ȅ뉲)u87I���S�l
�"b�wl��/��?<�ٙQĉ�b�=#>
d��ȼ��A��������4.>�LW��@����Q��<���n�������x�F8+_rS��/)���\�����8ٞA�'��#"*?H6�=
���7/��F��=̦뫣�����O�q�1���5~��Ӯ�����1.�0��܁�)�g��UjP��R42�K_zb���.��6�؄�@����|gXwнۆux��5Z{�>����OY$քvVs`��҃�龬�ap� <�	�9�����V�#����F��x�p�9"����.^����߃g���y�Ǵ�1�
��I������ZǗ���ߗ��?3��d,k��n��/]��|�kHF�����*�#)I���1KI�F<����<��e�<��t��Y�:�Q��q�k�b(=��x�ɧ��Cz}���L�k�Q����<Qכ9�~)+��lk(�K���|;�I9�	7=�~�9)�s"��a�X����!���6�b5dp'b1|!��1yĘ��g�X;���f��Gqnz���}�4�22����;�.��9�{�:�pߨQ�F��7� 5jԨQ�F�5�E�=KE���׊*��-�`Jw~�Bu��RƃS6�����uI$9,�����z�:�#{���S�ב \{�S\�����P��)R��*�����;E�Uۗ���N�����/�QYq����m�^h;�{��\��}'�����2�S�zeqt^L�˳⛓@�����>���g5|�o˶���)m���씫Ogs܆�l?a��ɢ���I��)�L!�Ӻp���a6�`�f����ä���g��|>����bN@yz�,*#m���/~��	��Y�իW)=ye�-1~V���/4���{Agt��ꡩn�@�Fx T�Ϡ<��� v�f�-���3X+���(݈%�!��X���2�Y� `Ua|���Ԋfd�冞�����8��;��^���^St䕏F ���3�$e�2�q�{�;��Z�����D r�@�z���F��(%���C����>��O?�$�s���H�~Mं�=�5_Q�V�<���xa�SR D_k�q��΀BAo4N�(R ��!8G|س�ȳ�!��Vc�����_���0|�pooo�ʾq�BC�70�%L{P�v3WlȀs��!¡���F�P��a�m�M�9�B��TF��n��]�$ )9hM��/`T1sF��k*� c��<W����Vc/���J���6�^��"�l>;�	C����^��^2і�-�op�����(�m�{�CB�!L���ｴP�����8��J/��A���T-l̅r��͉籜,�!�qO�O�E͛Z5���J_���'Fi����P�@�姞�u���w��x��|M1@�W�e?�!4�x�°��w`1�߸q�@ל�?280ױbt`��H)C���d�z+��$\�re�aǴ�0j�0֔fE�
V�yM��uI{˳E�!��B��<�Z���r�����vu�m;����wT�P�WeB��y= �����We����0���#.�^e���m�T���P�5+Q�em��d{��!r�=�9�n�ށ)�$
�y��	�I����O���F�͑>�E>Wp���<_���\���}16�sy�Q���?�B.�>�4��d�]Ϸ��4ۨQ�F��_� 5jԨQ�F�5�iA��̻$����p5u�i^%Ī�%󆾘�3�`���\k���Y�6e}�φ)��֢�Ӧ:͚F�	
h�6����_NiW�3[�+h
��t"@�L�(E��v�j
>���gU��X�u�O&7_�l�c;Ҟ�ի�ك9G����=�s�&�� SFG������s��_y��1J��6�:\]S��Tӧ�9{� U^s�۞���YZ�\�r��Q�U+��&`���84�]
���!����<ZAD��p�= ͡�W˵ ����A���|�K���	V���I���^����T�q�PɽZ��A�w�
�Ӻ46y��>#�}g>�s�	aƎ�T*�;	��C#FK⅞�L"��L��)�?ȣ����8��<V��`�>�v4�%����C�>y�KBb�C��o��'�����q�R�� � ��A����s�0*�o��}��`���Ȑ$�5租�9�V����r���{�K`9z�+���4Զ12&��Wɰ�@@'nO��y���0fÜ�Dc��݌�ܣ 48�ṡUg�5%w �lyt��>�я�|63>��'��3	$N	pxx8��'C
l�RN��H`,$J��ٞ�����?�U��W�s��C�+��X���7C@�ǩ�N�1�0��a-F4� ��˜sj��N�"h�*2�
@Fa��OД�<��~����4�R���|ft�j]��{y�{\��.�h��M�ײ��;C�(*ܲN�7\�K�_sz�f����k�)�W�|@a�y���[�k�v���=E��9��a.S�8��I���o��Nq�ʳd|�9��2�Ǎ�e4�{�=�������0��M�Q��~z�Z�����jLz�I%U�,�?�v�zc>����^ ���L�?�H��FaUE���㣣Y�|�v�΅��k�" WQ$�)�>�yP��[zz��}QC�{_y;���?tL�멵Pd���E+�u�X��kUZ�˾
{���6˲.��<l'1������PX^M�_)?�~n�eM�K�oj��g��$�r�sz�N�-�/$X���@�����l�d1 ������C���S�?K��SN֍5j���B� �Q�F�5jԨQ�[��Nr:��2�Y wU�)��"%��C%*�8S�ʢ���RmR)F���J
 �SP��P��R�)�)��}�^-�鷂��=��Q�l�J~7��s<�U!� ?�t� �NQ��U먺�h�i��#�kw�����>��(��"�
޺o�-�d����X�ו2�PI�Êת���K��z&�`��4E�fyg��:7cÙ�:*�
��&+[�^���=6�(4@�P���a�	8�u��>�p�ŋp�����s��͛pp��%�e�_"S�"r�1�pU�E=)1�y pUs�'� �	Z8�o2�=���w�>�:foO~/2�`@g�q@�(�������~h�)�M X��(z^��^a����B�Lz��g��-&0�=�����s���]G�	лvv ���x��7����	%_�T�6�,�9�8�m=%Gd]ڍs�����&��<걗_��WL�lM�h�x��������#؎y���=I.m��P���j��F�g�8�%�3�C��I�8�$�^+���#pnt6
�9��vi![������F�h����^����@OF����<�\���A���8d6�:�M�A�0���f�Bc>� 5w��Q�=dR4�ˮ� ö��f�5����Z���g��L���G�"���z�����Q�e{f�Xm����d�r$�J
����*GU��Ĳ��L��^�K�ߟ�r�k����Wߙ� 2��:��1��3���J F ڮjoT�r��Tk.�A|�������~���9T�Ԧ��
8E?K��T
�'2���*��}�"7�����h� �Q��v��nk����q��ڱ���xs����Q����p�g�h������L�_���i�"�O:GE���X�g�\�2��2ؾ򨞵�<���0�m<�s�l�ʄ��M�xٌ\�!�k��zj0���>�(��ϕ�	e�9rXi;A�J��IW�)C�F�5z^Q3 hԨQ�F�5j��#t���>dBϊ����
yp�.��V���| .���{AA(�+e�|�ɽ�*�q�}��a��SНB%����y+Q��*@)7�	�pMaRm��O3X�`wm�,1���<v��\6�2;�BZǻ�FFJA_J�cp:��e�&�1��S�0��FTC��; }m��#���Fc���̓x�,�")/��ß�\B�+p0nk�`���0H#) (,~' /{w�y����s����M)���)������8Z�1���`@*֙�?��p�g��s����Aa���B� &P���m�n4�f�:_�INa[Ѱ Ƶ��^����Ƞ�$�w/b��k]W��u��p��^�Y#л�Cm�p�E�/��؏���x�G�Z6`��etG �r��ݝ]z���`��)F[�Q�D2���?*И�t��� l�	�b�!�AF2'�g�ۆ~.s3L�j�b��m`����G�����Ҭ�1V������9��l�yL��Vf������l!�ر)���)�tƾ-0��H�sz:��Dk��B��2�L|���<1��mo�-�9]�l@��5�n2�����5^Yw*m�7�:�N{f�`,kO���^1J��l=I6��=͐�,�P�e��tC՞������J��8e��_1��6oxPƗu�����ʤ����(�8h���QMd+-g��t%�����dߡZ�c�=�u�}������@�f�P�a��ȡ藣�m����dTY������Ę!@Y_��nt�	�.U6���3G.}���I����R.2�S���{�@����R��=}܏�}��+[Pi�7�V{7��\ڮƺ����*�x:�!�����$���j��=�R������X��c[�U�������)��;�pHnט��֩�x)SS'�A^=:�5j��B� �Q�F�5jԨQ�[���c�#�ﺛ�?Qɽ-�~�DR Z/�T{^}�E�j��i�*JU�E=�{2V$r76��0z�~WB8Q%6~o�
���ZS�2V��S��^���z��HO>}?H�US�gז��S��w�ת{ύ�7�P�>�,��9�kap�g�|��vg��WC�Gl{�$����N)�G�~���&o󎽱�+���u���5����C�� ���1_2y��׫5ݣ������}?88����\�����)4�G ���-�˖(�/���~�_���s�E'`���� ���=�)L5�8.#x�����Ϲ��/~1`h`�#�C�����j�:���J c�����P�z�0�|���l/��_,fp��.��Ã>7�߄ãC���?�k�x^�E�CSs��7��Es[c�_�Ne�׿�+�~X�)p�m���ݜ.�=\��݃`��P����Y���M�����@;������KiN��_��(ʽ���gPH1DX�p�^�5/��G̋�^���AI<��Gd8a �ʇL9�����
���(���[����,kG��#�pH�;{�a��C��q%r�d`�~��^�UASp����<�b��|�h��X��ҁgb�A0����#�Eƨ\���6~^�l��g��SY��'�[�6.�4Y?շ�v�xk<Tc#6�?�#� �=��$ס���H�%���o �e��󙴐ۡ�î�|�s�빬�%pנ��U������ո �X�e��F@�kr�螩i�G
�6���1�p�#>�Ϭ�*�r����������o�a������
�Kue@�)�E�R�FhȰm��wIJ��ո��:��Uʗ�9��s��e�o���,���W��uu��eg�+��n�υ�����X�膋|��f��gw���	k�OK01TA&�a�������d[{�� �ШQ�F�^`� 5jԨQ�F�5���}��ѫ-�1��J�x�-�,5��{9�r�k����J�4- +��HAUy�;�1�+4�
���4��
�1���T�n)L����G^���<��j0 ZD���^�G�Wt�x�l(�����B�w� ��YC�n�>W@	�}��>D��Ȗs���7~o۽���C^g�)o��Ц��h^]��V
��LT�RM�@��P�%P�� 0z��=��6�CܸX۔�xwf��a�1�~R`z����������ӻX���A�G���c�P�/�+���|�[�w�~v	��m�|���:�����r�o��Q��"��<�a�`�m���O)4�vQ����ϒ�Ŋ�(}J ���������s��_"	v�/���Y��&Q�b�x��Nc,2�ViV�L�h p��><��/����������%�q�����˻�?�mg�;�}o��o��z�������;G �&��<C&z����=	�3�º�T#}��	�#��%)�a�\BD���%/d�
�� �5 ���c��?BcE(���*�1�u��� k8�M Ȏ*�#;���~��W~��C��*�$N?�9l1��.���o�����/z���{<�3�f�O�c� %�,��S8���G��kow14bN����b5j��*�x\�'�mֆ��۔,��O{n�{cp~۾}��<	�?��ب��@��� �t�,��2`ֈHv�ÔE�j��,�'���~K���/�,'s��ѷ)�e7�� Fa�����ԍ�#W�f�}�dgf������L	0JWS���u���T�*c�`1��-[{/h*+N ���f�%I���z&М$p�c�8V�F��Ɵ�/�8ݓN3"�փ�92X�0��	tM�}I�27���$l�������ۑ��`�L�c4ip.�.k��Y����:��3��Qǃ�C;Ǘ�ge, �s����3u�Ke(Wel3*���7|�ʙ[��I�,i���Z�F3P�a�����a�O�	�\tQ�Y��fQrw@�F�5z�Q3 hԨQ�F�5j��֣�(�h�jeV�X�|{�s67Ŵ/�dE���^�N	��E灮!q�6D�U�g�4w4�{���+?��V�k��T���I����y���, "���a�2�h;���h[������J�㹞��D�� �6�~�p`t�F� q|[O�C��͓��4�W8�7���省�L+��S�[��K�^S�qhgdҜ"�K^�����g�<���*4׳�m��5O:>����w8��w���T�2��A�ڸ����F���_;|�!�gx�ۜ��s�x�� h`��;���c$yP���q@/��8�B�Z���$�6_�A�����6'��Ǳڌ 0��n��B�@ )�>����
揨���T�\�p�k�Ͻƹ�v�������8�=��cM?O��κ6����_����_`�����6�ӊ�E�ld���\�F��hހ'86����U�a�1�@b/h�����O�"��a�y-"���~m�2�:|^gI����,�4bJ��0�ṣ�Cj�|��r�� � �B�p�ɼ�y�ޡ��n���7�2��aXVd@CQ �ʑs�`4�%�M����李du�2�@c�G��;r٨+Y��:MʣvmʌiY2�\>i�f@��O���z7�M�{� � �s  șIDAT�x�?�<E��!{҃�X����{+�7y��ZC�9ޣp�٫9��~��jǺ5���ֳ���Y5�
eeWB4�5p�f���&�3
�l���<��"�I�mH����ߗ
�	j��}�����C�lr?�=^z�Vn?���lkQ�qm�� ����T�<?>A��4��+[���s�7���fx cU@���q9�h�1縍�K5>w��^�g�컎�[�|O�4��]��|
���B��7����yy��훩�e꾍��u['�����~�\�����+��0��놩lpϨ�S��Bg?�6jԨQ��5�F�5jԨQ�F�nA��H��o
�0��3�f�r�a� ~6o�W��G�R�S�Zq�IچQW��1��H�z{��$O�qY'ՙO��Y�jr`������R2Hnk�*_�'���.�h���k
�P������+ gP4���g}�N����V�᫣ms������ذb���hvj[�ҷ�E z>���
+�!����ہt��r����E)�E�z׆T�E@k���$O���UE���ԃ��
���)���_�����[���5��!H~��s.n%�0�WЛA� kb���+��7a�<���!I?�s>��ǒ?Wƙ\�
����8/��cڅ~����C���牀n�A���"p�B�(�@f��~r�����GG+���|�昽��j)ocɽ�>U����Gy�f穬^�3-}'�j�`b�ԇ���"k6,`äCy/Q����#׮^�Y�?_��
#X�
+��O��E` E"6�bd� z 2? �����pxp�KLE��+�3�4� ]�6<��3�<W�݀�smBf��Q��gcO�L�Re8F��B2p4�@�'dl�����il��
�Vꘒ�^���F��p_˟4���mrn�����m$C�I�mr�,Ɓ��6~O�C���?�/�2��z �\�C5F Y��_u��*k����e�D� :�D�մ<��d��b��8�h"j��}�
�C=�R-(��ݬyH#�����#9�["����k�Go��P?�gwNҳP)2��RS�v���7h ��FZ�"��7�u{�oG�󘎛�76?ۨ>Go[O�9,��N��RNmh��N6����L����գ4�I������_,o���I�˺5X���E�&5HV�{_nY��m7���N��]9�{nH����6��*��J;�[�P0jܰI�/6D��vvK-@�F�� � 4jԨQ�F�5jtR��@R ���B�C�ԝ��d�P^�i��j����`���整t!����F����O�Îk�Nq<M� g��4``mgGC;Վ�뢬�����U���rx^Uz��

R�Fj>[�!��& �<����'����NN��ׅo���:�x�8/���*� ���K��m�O�L���Z����J~�sX<�����K�~�:|�#�~�`��(7���s��<�������Kz*+	������㛍
�ay����C�z�<��3�ZrzMGe��El���������W�?�Sx�ɧ��{�z]?0�l���A=�LVpېד�Aa��E��8&/ul���µg����kp���al�yc-^�2�V����u.�	�ݔ뾇��Cj�o��7�^L:
��}�QZ�{$?���P�
b;:��㈡�	00� ��c��_��{>������I��*8hl&�C��=�������{��~�K_*�[:�8�0�8��$6�4s�P��B�ޑ��)"���?�ԓl 1\{�3�����A2wv1�{sH��x�"�����O�}Z��]���(ѐГ������֜V@�������9�h�r������b���ݽ��8�^��^t�.�Ô�[�C�g?�yW�sFgd����0>�Ļ��9�۹ ׮�S\��f��G�B��L�����ey���7���Eg�3��9�`��=-�O/u}j�O�hp�6O}�� j@Pe;��˥P����Bc���ᗒ��\W�=/[X� ��N=��h~ò.S1h��6pe?�t� ��-k�w�Q_��3X>w~�+�@7<�<�y�\�z� �k��'~�8Z��g�*���5m��d9m��j$�H�N���`�� �Ep�ƂE��Λߖ�����l�t�(`�"�7�*�O��g�~���ψ�^�}v�Z�py�� w�&ܕ�G�LRu&��� ��/��c�6� ��+�	{�>_/��2�Y�S�y�g�^���-�`�����m	�b���G1��]C�5j��H� �Q�F�5jԨQ�[��@���w�1-Y��l����<��<��=�\pM��)`LE�XY��/���� ������>#h?�}^+:�'y��D޸"��l��mj��(T�B(�e7P���E`` 1�`��ul6@��z� ��؝ޔ~��9S?֣*��!���4��q{N���>U϶g�=S�6�Ю��ώ�R������8�s��x�����[��ŜAu�@y���$�hh�,p.{v�GBU�Q��SNuď{ӾZ� ��Hy� ����<��@4���>����/���9���a�8'��&ȗ�'�;����6��J���;�a��p�B��#����쩛tb42,q<cS���P��������C�}�Ø��n�T����B��
ؿ�uD��1��54�X#0k�WK�cZ��q�a(��b2N���(h�p|���+�
��?���8���Hsk���J)!�@�w���"���ptt��7>7Ctn����{����읣��Q!�����:�U!��B �90�ȾE�.r���(dxv1�,	�y���# S��zx�;p��UxϿ�w�裏��0�����Y(��Y&��Ia���Fw�N�(�5`�OI�^�Gq}`��#X�Ԍ��!���Z�y�I1G�3^V��)�!�ϸ�e�8I�z/�jz�8��9�kl��ٯ��{#,6�T�k��Н�q N}A�n��6��9�yDc!�z:���iO�+l�E=��P�9Y���aL�a��V��h�2c�[$���C���� �R^ֳ�����Y�b�������:�0m�iJnC1�(�K�!��Y*�v6QC#�?�:⦐�u�AJa)y~|����,�!������]�A��nyǝ%��3z	݀�bByB�Mi_:��d��j(F�:�a�}�|�C7�灵c�>}?�~��n��11ぐ���s�w��k�6�����3|�E׺��{v\e��D1.D#��j}6�ݨQ�F��W� 5jԨQ�F�5�%�����Eq�+Ȋ��k�lR �R�/HVP%�S<Q�b�p��Ȏ�i�ע�Wu�&�B�R�f���(
,{ԛ%�:���K�M�b�A8����LyhW୻7��w��4�4d��P:��E�];Ti�ir��*��.c�R�}�1��L*��6e�'��`U���m��4�5zA]O2�}��X��c<����޶���)�xN�80�mެSF!��f{{E�e�c^ۚ�)D>{��u/|]^g�Y����:�j @���=����Ÿ@$��H�Sl��6���|O�<F.�8�¿�#9��W]��P :[D��s�� s��g���)���h���4��Y�(,}Zqbw��(��57��W �f�"������&��xn�G����P0��5�.6Y���K:�؎��֡U�B �ulC�؃=%���"^�A�b�I�(pH����f�پ&�ӵ��d�ΰ@#�( ��H\Z�!��#�wb4A�Ŵ 8�]@,��H)Иb�~t�(�BY��\ �0�������ܖ����:�kO=#TD��1�u����P%0h��5�\��,dI��B㍁�_h.e-���r	s`#��"�f�a2(�����i�\2�NC�o�~�K6@�M9XI�-����mFZ���{��)C.�>a_�{���a����{�����9�wԳA�N�̃(_��b���=4ux�#��IDL�����x]�U�5��<�[^��"{t�#� �Xz)�̀U���,"���+� _�<��:���IP�n�3���� �h{��{�S�:S�Y�(`k�����H8\s�� �y�����d.{�Dqycѓft���	8�����$����,%
�E�pe���گ>��+I���4�e>t��5�=���`3n���Ѵ��� {�h�*�횥�8n�S6�F�Mvz-��H�2Ug-�w��)p�c~
T�|�9�N�z>i����y�?:�!�^�F��kt��K����q���v�7ӮjF3R�ぜJ4�,�8�\ϣޑq!����@��eJo�Q�5jԨ��@�F�5jԨQ�F�0��߇�T��s_æ"�.��N<�H@=����H�����^���Q���Z�\���IcPտlG"�-��w����躭|��������]3�hQ%��=W]��j���T͑z���)m�:`V>zem�~1��b��V����>ч�վ��OT��=��+�?e�L�6�ԓ�m+�$�⃩�6�_aN���>��5�x�儁�B��9�oI�O��
�����^���6!�g_�0�r��,�����\%��+�G�P���`��1)m�+�.�I��e/���jg<Ə�[�`�GY����SG�� ���*t̂��7*���C^�"�(�C�7�C�[���D�����%�5Dh�|Ll��=��:�8�L�z�Pi [�9T�\�����C�̓����0ΐ���ٞa�6��8���d�1e�̂0EsC��qM���먞�	�ڃ���QY��32��x��_@5�_Oyq��lij}̟�����4ڋl����������)��$��������}��ֽ�D��������º]�̋�8���A#����*w$o<ɞl#A�F�U��� 3��g$0z�i�:�UJ����WȠ	�����,�< ���yP�B5~bx%�E��H^��OR��v&tU�S��Q ;ƹ�MJi�٤z>��J���r-�]հ@ۡ"X�.�@G�!2��>� ��� �,�RUfp�)HYw��,`5�e� ��~$�g�)��[���=@���]@�jxaY�1�2�B�տQ��$2
�l��{*~�{�m�N]ֈ�5y��n���)~n�,9�I[�FjyT�?�d(c\�M=�W�nU���t��ʟӑ @�u��.�0%��D���h½ K{��ٷl��6��-��b�g�F�5j���f ШQ�F�5jԨ�-LY�l�;�p�&R`A�'芦+{N��^+����M��)�4c����S ��7�0oQ�A�h׸�,`Y���b��F�������q0)^���p���	M�^�f5}^�ʠ�`^m��x�PB�Z���m�m�w���i4��� �q�StH5V���U�p{D�̓���	7�����v��J��C�l��
�:����2���f�~+9��X>�7	�2,IT�ɞ�l7c��r���	�"�5�����^a��j�6آ����w+?P�,^�2��H��zd @���m* T-$pC�>8Pǃ=2c���<|=y�3��Y��B��$l���
�i���2��DEG�Dxc 6��GW�F�x��:�"�h�n�p5:�"�+�	z���1d��}/{�d�F�!7�ﮗ�o=�8��$�X���l|b��Zz��<`k#��s����~5��P�,F['���QV��I'����;ɠa۳������x|ƞ�10��|��-0�ì#^ ���t��'#Y w�93L2�����ۣT*n� _�����_� �}��T�j��Ã#�|�x��e���>�7)�,�!���"m�
�d��|9W�&�AJ�AQ-���j<�(%x���z�w����J���b���1H7|N�:�� Iֹ����#P̓e��u�ؓ��m��X~1���"���Fq��Gkާ��uV�<�n��!�D��y5�� ;��Qn��RD,�/�\�D��]�m�Ԏ��zH��Gg
(���;�p�e�}eOP2C�-�h���)�p���FSl�DƱm��9�U�T�w(�l��8��n"�P�N�g6r[��'���F�`s8*�qv5jԨ��@�F�5jԨQ�F�*IHm�U G0��Y��:����&h���� T�B4�lnG|}D��Ի{
D�֖m�|OaBi�H�,c�X������ RO�S�Ft,-��y�2��9�JQBO���7p�jA�y@ռo��񽆱D9��������x����x���i��E�*�p���hu
X6�����  5h�76�c��ɦo4�čo婙u�U���F!(���[�P�	d}L�%ޣ���ĩ���=�K|��E	�_�b!9dï8�x�V��e�cH��E���(��ԛǏ<�u|4�7�m�@�q ���+�:yo�t��}Mсr�K�x	|.)� �
h��G�"���P����"�H:�\ r6���P��|�h��279K���!@`��AF��ŶC���>�F�LXa�U��,T�\����]�hwc	ENu�6�b���Q��,�����]��A����c�||�4��q9�[e/?`c_�C����:������:nc:�www�o|^��W�����'>�	x�gܟ/<F#�����ϸ�n>�{�������^K� �?=P*	\+(OV����h	7n��>�Qx���װ�:,�!��i�a�ֺ��T�ls�����0�,s��Ub����R�`T�8�s��c�H�-�!�f�9��l�[�Nd4��h:�������I�%��S�;v׷�J���,��J<��`���9D��������8�.��4F8GG��p����?�7H�Ւy+$�O�!�M��C9~�2~v��r��|*�=���:��좎ԧE������B)�[T� ڂQ*7����Ϗ��wt�6#f�b���*b����<>F��|�+��p�p���XP���E����2>���ѽ���^�+a|�:;�!ox�~�Q�F�=ߩ 4jԨQ�F�5jt��M�% ��
��ZIG
��
�<+�6��J��8ȥ4�g�QY�������+�����Si���d����
ox�+�9�gpJ<+7`�m��Q��Qt�� �gQ�9٧ ��Z�|N�ܦ���ʁ�US�t�z��/��/L�������U�N����:��W�;>���'�����:��d�#?o��������yy�>��?��_�7e�*ēx5�8�?0��=���ͪ�V��+���8�w ��,�O����]�EQ��f3�l2j$M��� +�Ǒ����)��� ����Z��x���y�y���!����R
H�sR�G�/r^���6�r͐1�_<���r�9�0�Rgk�zv�w��9]A�(�S*{�+�G~�h
f�R"Ndk���(�w=F@�4
��q 7.������[XH����s�<����u�C�Q��P�]��D(4�x6&��C��u��:!{�N�������Y��-n�&e�Ğ.]2>�-�����{*ii��?�݅�Ï<�Vx�;�	�=p�aF�a�������꿄k�^�n��j��� (� ��/vv`o���������s���Y��e^k]`�{1��|�{��9��o�6��Ew�/��?���^��t`=p��R육D��Y'�΁���1����o��/]" ���P��kשM�j �Z��#�I��1Ü�=�<�����CQ$�g.?��k��7�M����b�D��G�n�����:���Ad	�a�H.qd=��=�kB�_�^L�0�-������䵯�����p�]wsqa�6�2��"�����4��o���� ��J� �_zY��[�e�*�EH{�� �ע/)O�Vd�|�c��|1�4��m���}p*<�7�A~�'���*�<�Ǐ��^~�G�{VA};ÈW~P�
 F\*ܨ��
�]���o�e����Շ�<gm��S�� ��Q���n�A�	�wk���A����<ߨQ�F�^0� 5jԨQ�F�5�)��@3`ޖ��2�U6<���x�J2���k��aB��K����|a+�ZԀU�F�� *�z�C%��>M�c���?��W���4@���N��>Y,͢�V�� ���M?��B����"�+c��SS$X���x+�����͊�����)�Ä
sZ��o�g�?�q��ƞ�e�j^��N�����N}�nS)6����y!�v���������.�P�ox���c�����L��v�_�x�u�Yc��>�Y�. 4����G[=]P��(���H�� ��QWw�o͉�3�1P�&�P���Z�8����Bnur�U����B���S���L�:�
(������}���P���}��f��6�h�y�i�:��mD���A��^&���q�x ?D�P's�䂖q�����uKTy׀��J��-�E��Ŋ�x���&{e��j���mޖU�6��?�F2Ky���4�O�i*b��w���#L�˾ܱ�۸��M�߿	��P���`,��w���_����0�?�ݞ��I7߁o��o�7�����?�3Â�����0z�� v�G����qz|.g�`�.C�F����ë_�:����N��_�W�w��__m��*�+�cJK��7���ܑ1�����/{�푷�[��f��E/��D�~�*|������߃O~�S�:^B��@X�1 ������ï��������*�� � ����ӟ�$pZ�^"�ຈ�����Y*"70���\��9E�������կy�;������g?��O���!t����� $M�����b���G����-𒗼��
vwwh���Q0}úڃ�������{-���(
����1@\S��ٞrJgt�(W�,eǦ%�_��Mo8'�n��n����gSPɝ�)Gܽ�1:���E�����ϗ&�˺5)]�|���w�/'?ʺ��"n�[z~�+}��h<z)g'>�*u?�a��BݟR<��m��/�g������C�gU~�:�''�ҨQ�F���� 5jԨQ�F�5���&\N�|��G��h
0�'�R�P����� V,��i� +����Sۊ���^a(�'�������Kyہՠ�OV�K���$��	Avr]a���@W��@8{�@�c�Z��ۮIY[ꯍ
 n��
k��d����,!�ݜ-��g6�h��
~<0��U9�>(���ъ������!6�s�4�2=��vLވ�g�獻���졬<4�h��o����￳!A�s.�}@`��UVpG{N�MPy���]+D�y�w�Զ�{����գ2/z[��Q�R��LӅDJ���x��-Y���\���~�w���^�&X��1��7ƙ�؛,1�Y�yi��&��\v��p�14�P�>)_�R����MN�H�k���?~�� y�a�q��:7śs�:A )�����6Ԋ��50&�}H�-k��v&�G��V�J�<���"#(s�y���vS^Nɒ���A��Bg�SSm�j�}.4i����I�Ø�|������.����8|���L���\�4��yz�Z�lx��� ��������b�A~],v�U�~5��~�B��Л�_��i[�~I����@Q���.��;;;�-�-o����?O<��nBF�� �7�[��0'c�L�b���w���w���|�.�$������w�s/|����}������_������sH�
����`����������_b�|l�l���2Ýw�5�o>�^�(��P&r�|�B�QbY1�.t�Y�RԄ�?�0�7���}����?�%E���������0�G����0���E�� ��@�=�����]�������h	h��'�4<Xwk�����}������_�7�A|@�	�|$�S�|S7d�G�)g�A�S�Q?���-�no^��_��}��8��lԟ�5i[�;Gz���V�a��9t�o�}%
l���}I���?�' '���$JWe� �Lo��<�z#���������1ؙ&�Ӳ�Sp�4^ʓa&5jԨ��@�F�5jԨQ�F�"�I��Y��B�+�I!ǀ�)ǂW�	�6ҀUP�ꖼa�
��īi�������d=�y�4��OL��`��2�m���_?w����{�0SC�rx[V@���J�_y0uڣ}|Ϸ[�T+۽�����BS�+��pM�,��Q���6.�^�P�C8�]6���f0���W������s����#>ec���o����P��P�Zݾ���J�ڀ׬F.�Ӏ����
e͙@sg�]�� �ƣ~��<�"	� ̙%5�d�z��8�0���C m �uP����07�Z����YA�2*[k�����L=���o��vį���E6ib��[���RyO�9���1<6�'x!�|���!(u�3200^
�0#��஍���[a�qY�diD��R=?frK;��lBlA�����D���oTm��}��k,S��ja�ޭG^VM}��0pr�<*������z�/�'��W����S8��u3�җ�O?�4�랼�绻ЧX���w��߃�޻r�2�/��{�؁�}����F�2��/��s��߇��#2<8wn.^��9��5ɝ��k1�C�9�x�w����'D�W�>�|�#@G���8�{�������z��}���N�D�4 O�V	���o���~��������}y��^��
��G�2����������0���B��DM�"�2#��OBC�w~�;���_%��X�f"g8:���ɟ�{�?��3��4G�jBOc�k�ܹ�p��w����M��A##���� �ဴ	���wN�o|�ۿ��؇���w�b���`C��o�U�jY�'��m��My�d���7o�%��_
z��֞"c�e1}�$�Xrb�4���1�c�n�\���eA�x���`�m�A�(r`��ᖁ�T��m\���HOy��l�����l�\"/e;�x���:6���ظ7A�F�5zaQ3 hԨQ�F�5j���>`
����b`^VU���r�VK)�ۃ�a���n��M�޶c��0�$�P�k��|]��B��g}]�6{��&l�S^�Vz���~�B��rbx[TP���xs�=峭�x��Ӄ������Iߨ �z|�2X�|C�X��(���Gõ����bU�[?nňD<���o����F�NŰ���1�?�V�Q?o)_�w����t����F��l>���k^ȕ���|��J3pQ���
Ml��˥\~V=��,-S5ڮ��]	��)ryO� h��'���<#��G�@��e�~B��Qc�E�!��
Ġ�r|)�����f�� ê��Q@X�	�3`�ms @�݅p�S���8�����p<iӒ����8H�2�yֹ���]hj�9��k�Ρ^����e슇�/s�ȆnzO�[���b4�y�knd����?�Ԉ��')b̈4̷�ft^�2.�o�w-[@~��N���	�1��M�7~�dP��J�y�o��Oy�9�u�p����-��pg�3|��O��/{��h� ���Mx������ ��.����>������Ex�����A �5|�������Zǋ�h�����G}�@�>��O���}��gɀ`ٯ`1����=����_����/%������x�k�>�V��GE3��r)�}�3�O�'��>�Q\d�b=��
�
E @�;�c��~�(���������o�g����U���T�p���+�v���(�ř��T�1h�@�>��Q~�}h�p�ҝ�C?�7����F�et��\��0[�������?�y��G>H}�vvh��z�������\���߼q��3��X-��t�v��� #�'R�sx�[��Ї�����L^��b��(Gk3�,\�(rAd)�P�T*��l]ك�H�R)�a1�ǿnȧ�5��0N���`Q��1�69��Ln�����!$Zڥlg�����k��F��ٚ��Ɏ�G�5JcHp�׽_���󷖣}�85�Jb�����,���h��ue�v���k��4jԨQ�5�F�5jԨQ�F�n1�@�b�R�<�
���8�	H� PO!
)) }�(�����&�)��x]�X���������SBeҚ�YsX�[@zWs� 4P*�zp����0��#�����s����}�3�~�J�M� ���@9h��D��UI���*E}�T@1P���56���žFU�֔G<����qN���*~���xk��L!W��)O�,3#w�+�9$���gA�Ɔ �ژ��s���e�FS�%���=���.+>{�ҾkT�U����r3�2�'�xV�[���?�Jt�jK��h��Jy6i,�+oi!ڏ�V\��z�F[x�ߍ�t��J��@����ei[0����Я-*KY�:��f�^؀��ղ&�l,��RGc�Չ|�;p4���(L�;:������FT ŃD3�K��z��`�R~h������G(hő������[�<>lg���,D�� �\�B��1�PLA��4�xEA���*OzO��KAwk�Px�Lt�xd!��X��R��Yt��媁@��`ᢧ���Eo��}`��"���i_uM~u46�ڨ�9�5�y|mlܧ�2C)���]>�|�~���_?���Y�C�
����8a�o�0��_/���O?�>�#����G�����ğ�9�x���>� ��g>�����(��/��)l����Yf\��$�ß�,�����vt<���� ��s?|2�1��A"I�@�|�n��8#0������W���`d���7������p��+���Ås��׽x�K���zX�"<��7�����G>�v���q�f��\'~\�Z�c8���y��ՊB��ΐ�5���s������p�hA�݁�s�����-���qcY����+8::�s�m�]�#BU��\����?��?�2��17��h�p��M���(
˃Gp��u���Kx�+Oµ�W�:F5�>�vw��Жw|˷��;.�:���;n��O~�	8X/�u1��1�70�kXe���*|��85�ԓ�cg;pk'�+�
��k �9Iw��yj��q��>՟�Z�J�=�5��G��+}��@$π��~]������H&Q�W�8�[[��~��5rC�sh�ד�/�@0G�P����<l?��=�f��*��%�8��o\�\C��8N�gH;xfR˘��y��V��_PZiԨQ�F/j �5jԨQ�F��bt��]s�V`�N���
xŞ���5�bC�Mq��2�&� }���:�1H� ee/q��NMyO�R@�:E��7�9+o�*��~�P8��� ��>Vj���z��
D�9S�+)`(����z��+�[X�R����Zm�4" )!�WP�ʘ*��G_����@?A��h��KPeF&��@�2�<���<hHdU�xl���F��N��Q���h�1|.&t�<�^�\@N��xJ�r�?b�&Z�t�_����`�69��o�Fآ2��NuMŸ�Z�֠Jx��c\�C�g����l�л�rF���W�9�~�;1*x�12��G�ܫQ����p� ��y7&'���h\L�gċб(�6Jd�7����\�!�<c�!�{��A0ovȞ�T&�5b�����5j�t'%hB
V���e����c(s�C�gL�=�*:���"�����M>�3e.�F� OZ���$VF���UW��Ƶm�7i:Z����y>�t��c�P�C�g[${�q@�w4�{��|��/�������\��vx�[��u���x���a���_z���w�^���o|#|�ӏ���`��9�b�9ǟ�����^�`y|��%�8w��;`/�`xw��;Og��Ô�5E+�)\~��~H�}�,���~���<�᳏?��A����?����x��ʗ��{���A�J?������;���� �_~>��O�=��>����׽���Gt�.aF��;_F�W�2~H��&ɹ�c/l��z|�7#��usJЯ���ÿ�1��3��W�Moz#����$)Vp~�������~�B����zx�r��E28<<��}�s�裏���������g1��|��0��_��b v�t&���6��5˞��%��4�N�%B}^�d�T���W���g�<���~Nk$����d���e�g|v�>:�>��a|�?W���Ru��~}{�y��s��l}ֱ���H�o��
���Go7:e�b�6>�궼E�ш�a�	l,ǩK"�S�F�5j�£f ШQ�F�5jԨ�-H9w�3B*�6u����Q5_�gC6M�(ϓ"�$@�s���
�
4,��wP.:��Ǣ�m
�m:���ܻ:�甽�P����/��h �i�#>QN�`ϲR3l(+K?�q�=��	����	��[s���b�?���ߖ'W}خ��so�硙�F#!	=FB�Ò"�X��VXVB�
�?�c����B+��)�X<̛Ā��E��^#�kF�3��}���oU���U���=ĭ�=s���}T��U����콋^���:m1Lz'�0Pj�U� 6�٫�a� �9�q��4�@"���(�k�4�EWA/~����YE@���K�	���9�j���u�� |g�U5Y z5<����� ���n�'{6��0o�M姤Z�R,���Sx���8J0��e�*�#�� ���RS�zu�� �ɰ����,�|+л��93n��A� G��s�ƺ9(F�Е�����{��%���櫓!|��HR}����j�4]M�i7�?�̴_Uw��(��(�0!�@�'��pQMc/���ul���/cѩx���2����A"p_Dt�3~t.g�ҭQ-��?� I�\v�jF'��N�~��,����>-ԮQ������B|�>���������M���V ��=�E���픾r�y��/k����G�Q��o߁�yT����'y��u�{=ڱ���n��K���羂����
[�������7n��I�LC���C8<w ���&�O�)���Nc��8�{ ����>��p�2�>cG�oï��onq���O��?/��'��x�����}�}\}�1L鏚=���������E��%����������W��>����o��͈x�8;�w����Ds5�ȩ�Ⱦd������~�|��#p��M�W���Qf�/����p�[����L
��-���9«��\}ի�g����p�ś�O������� P�l�mw�ǈ��70'�1��¹���s�&�]��n���ۑ�7܏�|we���)��T�>?)*,;�V�5�yP�gh�O�Hl�N�����j���~k����(�rx-��ui�|������w��Yנ��.G's4���j�.�P���:�96um��z˭��kJ��r��eJ֭2~��L�N�:uz�Qw �ԩS�N�:u����K�;��b4�x��V�T�3��o�-�7#�KZCX����XԠfxSU�ǧ��$<.T��tG2,�G�����eA۔*Qz�����%��"y�����Hadî�@���xj)��4�\��.N�g��,�Z42�V���!�;�I����B38�и��@��L�f`1�/��n�ϓw�b���襓�_
H&��-T%�څ�r�t7*�"����w����M��2VS���@R䳣��"Vl~	�+C�G�&��D���āJ@�L��� ���wpp��AM7eJj*31��L�,�\�W�RU����Y�I�0X"8s��E�ӱ� �A`YH��|��WT���UHyA#`=�������x���ݭ�a
HH��zq���mTn�8E�\g��U�\��!C��;;^� �D!Ka��3�J�O����Ҕ����T� �39JU�M��C-�����7�� ��;��}� K���<w=� �����oy?�9F0�
��Cx��kp�9�t3Ë7o�{=��_�%L�)��`�ay0�����իpp�������}ƺk��D����8�8naW��(ϯ&~��DNF%jx������> p~ �j�-m�Ҟ�!d}x O���x,�׮]�o�����^����wb��?�C����� O>�j䩔��&ٛ������&��0�68�N7w���C���:r��о��^St$=�}2��4�Z�`�P�������nx�����i�筣��?�/�S0���ty�#��&9���'?�xϻ�:�'���rvS?�??��?���P֗����$������8�P�I2�L��(�z�}t���o�t�(��i�3�����!%q�} �l�${R7*A��9W=���>�~QE,���8�f�@����f�y�:��͑���sÞ��ئ�['�z-Ǥ�~�9�:���%>�8�Ho�u�+G�ӡ�/��Av���%q��#�${}壇D�e�3D�G�/����Զ�x��ȡF�X�״X��H'u�ԩS��u�N�:u�ԩS�N�@��(��+c�'lN�f�m�2�����ڜ����$�D���:�����MI�)����
��h�veX⊟9�>gx�9mU�ݦT�6
�.ϝ��_��6u���3L��F�Z�u�F	Z�Ľ�o��Sb��� �m�D0-�I�v9tJR�V~'��S���U�Z�g�ּ���_ӽ��:x㶵dn�o�/�6�}Qc4�:����������g�,Þ��(! ડ�����+6E�ۗ��7���Al`1�$c!z!�N'nn�������tJ�X/�� Q|��q����9��ah�@ض�l�I�~;�����Ąb�H$�`�y����D�d�����ث������S�E���N[Y'fÒ�>�RH���@{��@� �c�F>8y0�v��HA��%��� ����N��,k����j���n�ss�~�ar���w���, w�%}^�*W�/`�� �SP��=GG��8 ̩?���7��쓟�q���~����õk��pz~,)�CIy?�nL��(�+]�W=�F����/�l
��Q��|}Б(ad>:�����8�l!N�SV���#�>g�T��0�8Ҿ r6�����Ko��Cq�y������Cx�����g���vz����g>�4|۷~+4ҹ�z�m�[����~ow8�uJ���;7��� 6�<W'�.���K3f�@�wӑfd�ɂG�M<_��|��?8m~|�������$ׁ��;����G?
����_����S89������1 i�飏>.\�۷6p:�I��/����M)��p4ni,+,X��"��}�{᩷>��A�J�=���8>�m��mԴ�������NP�PG!ֽw�G��<��r�T�8�WN�H���s�Pg�0�?�7��ۀ\��-���O�_g����~|�8 �	o����� ��jo��u�~��wW��S_�;S����{��Xj��?���A
��,$7��ܗt�K��v�ԩS���@�N�:u�ԩS�N �a�1���(e���$`4�9��"�$E�C��|(9�F<}����rXUn�����`��3���[�Kɥ\m���.܋aL��5��|-����g'+1���=1nJt�\K]���
kc��ll��u( �m6�,"x+��]R��/k="/�<XR��^�05�{�����t���U/�!�1�V��6��u_6 �>����;�g�������Yٍ�}�����u5���Wx�q!�h��`muA W/_��cֆ�[
]��=�x�F5��֎T���I�Pq4��LwHǲ����)�<�D�gm�K�_A�t�k?Z�4r�nőNNNq/�ɳQ n{4x ���=+̨��'���~���{�,� �q�4��}�S�޲�P�љ�A,�5Q�q%=�y����Mp�Ǡm��E� h�(p�g
��q/_�iK���zv�R�}?��Eg�{���g>�����K��4����_@�W_	.^�k�]��x�#&
���w�k�~	��ܟõ��'?�x����?�Jx��G�ʕ+�f�_����Gy�K��DWs�et�"���4l��y��鈦�����H��.���S;��]���~x����U��2����O��}=���'>��̧��;wn���
��� ���f9N �����y�N�Qp�����<����o~��O܎��_6��HYWl\��X��M����U��GLr�ԧ?�|]�|������������i{w�oã�>�m.�*��������}����K�v�)�?:[��u!�>�8���F<R� ��\��O?��)��X�|�3Oc� 9fŃ�Y4Up:���e�KR�3�t������Ҩ���ܯm~.�M<mM�^k3R�>�K)������eO��0]l���6�~��v�.{gu�R6�9u��cҴ�5I_���o��_��W)�~�7��V%#�p�~E��u����t�#���jŖ��OP��i0-5�S�N�:}�Sw �ԩS�N�:u����2���#�4�݀$�3�M��2��9�7�⨬y�jˏ� `nCk�PDk��z��>\@R5kT��*����6���@��%���;�V���{�d�� 3�ݟኑ�ܧ��wU*iG���=/�< �TUb(uF�(׹lL,�}EƷʊ�i8����J���׊�.��K��{��J��X�����[���h���Ւ�R�7�Z�j��C}}�fх�w�<s��"ۅ�,�Ξ�)�};=��Xb������6��2��Rh��FQ3ĒD:Ё_$���������po�AưB���A�(���W�Y�i��U�W�K��x�Z��*��6}��]f���T!��%��)�;-��:��-ˀ��4�:�I�]�+�7嵭K3��/4KsK���#+�$�c^��72������`z��ݵ�*·�j�C�yw��}2h����v����|ޫsQ��`e��+^��yI�e���	�����k^�Zzq�o|�7�>'#࿢h|�3E"O�>�����s�0b�D� �����X��R>;���3�Z>L�ű����=88d�D �n�e'�� #:�;�kq�d)xի^	�����ѝ;p��x�{���~NO��G"�V�����K�.b;6�y��0S���,|�w}���c0nw4�'~�aV�r�A�;���H��"�xh����}�Q8Xp:���{o���}���pp��^�G���֭�pr������0�B�_%S��������,ވ:_�m@�:&z�8Y�ևt����.����?
W�\F`��I9Z����ӟ�l6%���d�p�� \���`�6�;[E��P���
�]�M�ӷ\��qS��e���c�O˪yW{]�I<i�ԧU������7�s �1�G�:��X��2��*��s����@e��w"����c	���\�� ��(��1��I17�"���x]�3���<�'����6��:u��遣� ЩS�N�:u�ԩ�J��\#U�?��ѥ�TL��
�p�GV����L�&�m{���0?�^���X���D��c�1PR1��5m��!��㲒�ԁ-�y?`�btfc0���[�?�<���p��n1R���2�	�smP����E)�%},� 08cc�Ŵ�3,�;�5K�.<���+���������������wY2h��(a�@�Cm���զ}4���>�NYqФ���]z����9Jd��\�]�P���v"�l: ���؎�AF�4 Y#҅9~��y��Q��`m�`Er
�N���� *��+��E��8@_q�9#e�`LgB�lgv2�}�߽k�DyJf]_D�|!�n *��ڐA�%�c�Y��9^�T[;?�Z�̜��)�I@*�1�LQ�!(K�Sfo�Z8[���~\F7�굄�c��EU����f^������TjG�GU��{��-a��{��3n��/����c�e�93�4�{�q�l6��]dZ�a��[�pL?���B��hL��G���^���TP��A���r4E��柲�Y��g�@�8�5���Kb��B<Ź�dlG�s�I�v�`�oz��v�����v��p} ���B+,S��d/���ٌ
o0p��=X�v�	��pxp6'�<`ف��ΉW�iO���Ï��CEq,r�;��=��k㸅W��*F���o�y\d6m\W�<=�\�xn޼N�,��a,�s���Ib�:ПK����ë�|�j�g�m���;�?�p�Ƌp�9���!.놛���?��y�����!�}+�B�84U�%�: ���6�&m�v��3���l�����=�+߿����a��l��'�!� �]�����U�����YY2ԙ9���+9���?5[��hq�q��G�\�%~'�8�8��\�ׂ�6��:u��鯔�@�N�:u�ԩS�N �# 2���w�q\eW��R���=��F�(x��,wQ�Z�ܦX�vvMmmk��T��|vF?y�}�Rb�K�L1���F�*��@_��t����-˜�$�o���gв^@v������_�^�t�s�hVىQT@���g�/����k�]�?����l�|��Ҝj���c�c�C<o{���ڲ_JYK�D����k	�S����Zb�Om-�3'����Y� �x�[����	
Z(���j�G�6��� c�n|�5邤�D���� ��Pg�")�S�����_I��&�y*����
�ɪ�2ؼ���`���O�Ȩ�J"�X	��4s�!툠�K爎ug�(8��ѿC��q�5*z�?bduȢ�$5����t�)���X-�^%�F7J��:ne�7^�nK���Z��q>�5@�ً���(\�LF{m����%��N�����ƒn�1� ЫL ��}j�wT�kֽE��yp�/��S:�d�@|�`�@���)��n���΋4���n0�|YwiD}�=Q1�~L�+��hq (����!ܾ}��9 �]�N�vG}) ���Y*P���k�+Hf!t�A�)���D��3�SVC��n�g�#C9����''�i����[(�*���8���)�`�C�Z�t��f��p�Lu��sdP�8OPF�-�QV��ģ�ع��}��V��t�B���E^��)���!�>Y���]:6��L�����	�dM��b�) f&XMm*�_����?�0���Ji�8��&���?_��aW��v;�߶(�����b YX�5>;�9�~���vߨkk�9m�^Q�z�xP�8��D���������9���L�ȱN_�=��WaҢ/]$|�u9��Ϻe��jY_*XcCZZ�a��k��Z��t	+eݮ��AVX�g����G�5�����K�~-�7*'��V)�)r���0�N�:u���� ЩS�N�:u�ԩ�H�0d<�1���0�$- O�xؤ���`l�gc���(�<@�5�����5f�ɟN���������z�-�$�?	�C�t�:��/�h%K�����(u�|����H�d4@+3j$��5%��By���mm�<{�}��Ց����}�lBmcUk���a��|$[��{�BJ~Sb�3\93�ɲ=T��1DW�X/��i��t�KYf�n�v��g�U L 0�cu�ü�m]A��m���h#~��R�_���Q�g��t�I�nH<����*�y��T)=*2�`����5��ŋ�Z �������4�e.���-H k�rt��:����@��6�9st~R�H�'��l&�<:Q���d�o�G�ʀQ��-��S���TU�@�k*�LG�)���o�;�]W�*�	f�a��E3H�j@)�����'��.��m���UY;���İ �gy��)7����E~)�M����|O��{��g�V�gz���S��?w�ۤk����xxx�O��)g��`���s��ʕ+p��E�=eH�i�K��S������`�(�Rߥ0��ԛ;J%.�7P�1`�������s��Hz�D֣���K^��j8����ɘ�B�d[�M�~�g�p��s��0�~Ur�Ϲ �%mX�e���W����^e�T?΃����dP�"�# fKXO�Ē�8�q@�9��He]��X��a��t��V"�K[NOOin�i8&^�!j���;�O�+<L�8wx�[�Q�&M�r�����>D'�������൯}��`@%9�o���³�|q��[���&G�2F�d�8D�����v�Se��3�)�����^��"���6�1'�$���S�_{3�.��9{��R��s�FZD�5N��N�J���[%h,{� �|�1T'X�4��+����^zN�_u����3�z��政�'�8�re�,�B��յ�~�C�N�:uz�Pw �ԩS�N�:u������)��q)1,H1�����X�P��.R�g�o�S-
�p^�=9��Y�3VQ8��)�� Q:�aK�m��DWI�I�`�$>�����#]�N~R�{�#]�n����|�f�o�Ƅ�Rl����(��i��\\����'�K�� F۔�fP4��O-F���#R]6�%�*钵��(W��)���?�?}?�"�($�䡸߂��_fj��+{�¾���溼_�-��_'pX�Ft���������%
�o��:h��5���W�(���q�ĖH>�摄��Vݥ��)0��R��Oy>ԃL�s�{N1ʦ\���Wr��|�2��=�%���=D��zQ���[�t��P啉����6� �C~�{�� 딦>��Eߓ�5y��,�aT�<�ه��9��Dƻ�]#ё�馹4�����y��W�E,�81j_�C�ш�W��tU_e� ��\.��	`�/���<,��m6�}�Y��*�f%�u��f�[�Ò#���ⴟZ�4��; �r���ّ��/~���?�o���Ho�Ο�������o���~�T.-蜦>bt���	��^�vg���c���>��v�AGH����K֋2n.^��sS�s�#� B�����l";�PNs�D�Ǽ� ?�S?O�sx��f����i���>@�����?��?
���T��t,:F���a�Z!���qK@�j��;X��8�1	a�o`��]��ʡ�W|	vӠ?������.���_��o���8X�\2���e9�`,�V� �� �"����+����u�0L��������-o�"�P������������# ��c�ܴ7Xn��$�E��a�P���]�˕9n����F�D_�1����a����������t�v{�%}M�yÏn��暍\���aq����sz��F_	��o3�q���/HO�1���@���䚶!ϟ���a~�O@��.�������S���	D��<:u�ԩ��/u�N�:u�ԩS�N�@Z��aw���!r�X6��!�N�1l	X�""��&` !�Ϊ�(C��
,��=� �l�R�Z�P���A;.`=o�(wvI1΅��HdIAn�R��`�e����Co��(Ⱥ]JI4y��D��fL7 /[���vS�x ���鴃� 0��i^g�����r+s"UE6F^p�����}�͸�������͝��|s���-o�,�����*q�زIPx74�gZ�Jo/#g�R�>QA`}���6 *۵&��&✇r�͍�}+��&�����"*By�B|��`�_�����Ok����� n@�'�瀛(����@g�����,td�A��o��Wk�g%2��Y��,�:�oЕ�ת^9�@t���*=�:+U�΀�*S����na&,�=>rT�D�����j��T�}A��:��= ��s���R�h�n[�������w��i��|�5���s8FLq����u��ք�����/�_���Q���Y�;c��� �������o�v�K=���r�<S���9_vr�4O>	��H�lN��Qʞ�h����  ;������G��{���>cN���#����?�����&L�|g��S8ݜ��C�1�8��~W�\�7nM�Qĵ8	Eʹϼ��K�q@�!�;"ӵ�Pb�93I�cJ"�Uz.Dr`��=
�̕r};���s/��~�cp���{�`��[~._~h��	����.8w�<;Z%(�*:���c��.)��j����TN����~���o|c}\�������������v��n�'9n�h j��}F�����H�8���J^!�j����3��e�FK��柝9�[]9�`�ۮ-- _�����3G�=��cl$�Aq�@<v֥�4�V�2ct�0��֫���hmhy�MW��Lg��7(91��s�D�ُB��q���~�S�N�:�<�; t�ԩS�N�:u�� R�	�����i�3�Y5>q���D�����%K�J9r �O��6|m o`����ܾ#�ʯ�`���rܳVX�",�C��
���XE�2P��Z�]�PI��ACA}1jr�������\{삳��1�Ѵ�Z5���wU��~t��b<7Y*���0y )���"��W�H�6r�"{�z�����1���FЗ��<�v��{��/��Vg��oݽ7�� �c7���ë#�V�w�e����Ji��1�9�!���ezď�V?����b��_����`?Y�������^�ɾm�>癶kU���h-Hպ�!����V�u@t������h�<o3�J��Q�21�q)
p8�e��^�`�y	�"Q�\�5���p6����=��:�K�a��N�W:ɭYKYM��y��rV�zB���oX�n��_�˅/�!H�)�i�����{7�v����'�'�\�K�|J[X���=N���7n���֗��e�V�ŗ,;�o�n��d('Me=�����TƦ<���!x�y9�� ���R��je<3�_�җ ���L��e�Qb�:�J���,k��L��c�7%+A�s��0�^��a�K�{"P��S��*Q�-�)Sd( +rn%�~qo(�<���S�ز_����H#�FA2͌�~�a��s����8�s
'��t?���`u ��o���]�w����k_M�e�7!�!��U�5a�>� �s�C���7��M�@!�q��bf�_��_�l�w���t��$���ҧ�%�K��!��W�g��\%U{�cZl\�(z�9��R�ђũ"�g�LاT ?�z�8U�k^۲m	���x kǞ9���ϋ��,�6��� �P"�)+��+����"y�
��9ޙ�xPg]�l_mM��� U�#�t�Q�Y�����c	/I���󡬏{��N�:u���K��S�N�:u�ԩS���9T>��\?s��,��P�I�,��g��YJd��A�QBSnKfhg��$f���{f#4� �� Fl��s3����g 2VF����Ʉޑᵼ$Ŧ�<����7��T�3� ��}v ��2$��'�:L	����@@5����\�SѲ�=�"���I���\�U��u� r�6^<^ҍ��>*�F��9vD�Aj��Z�Ty�ge������.u/_w��8n�h����E.��k4���n� `����]�e���p�1��Y ���_����o�GP�"�sX�]O����*��;�7[#j���T7�U�-�m[����Y�XS��4/Mww�ʰ�P� E �5�$����W��1�*�+���DB�{�l� B�\?���w�>G��!�*gU�1���[�V�}F 7��R[�i���A����\;@K�G�n�ɴ���V.~M4���.� �����^�빎������QeP�X�X|�T�#�e��:}��|w�%<��qO{:���š���	\�r	�-ϗ4�'�-�sc*��ыp����_�J�7|\}�1x��5�%�=냲���c��?�CcI�?�9=�/|��ٞh:~@>�>���^8z������F�,G;J�?=�.�	�d�Jp|��P2h�~�T�����J��hυ���X��\�|	n\��� Rր�mTwan3Ɋ'����iQ�,�I��Y�:��D��]o��g��W=�J(�@(i#t�8 '�I��'M���}�����:�{%v9�u��g~�4��lw��2ջ�mM7�ƎӻC�c��r!]P���5 ��!s�yZ�H�(�uN Y��T��P9TK�y����V0�lVe��kR�^k�� ~�X��KA�ۛ�r�抙G|7��ǲ��^���z���� ��x�J����[���S��&�zd��JV^��� �I���Ǫe�t����n�g�S�N�:}�Qw �ԩS�N�:u���A�P���<t ��Sdd�3#���E�������Knzc��X�d�� �gf�<�Q�AN����m+��m��<c�
���hє58� 7���t/�����I#� �r��N#��k�E%9�!�6$}�Rн���əc��k� j!�.�V�J>>;4"_��Ɍ�bt˩��-��O�T����8S�����BM_+;��υe�-\���³֯2�T��H�"9��Ђp�3^X�ԩ��������^*�E�8l^��j�kTpu�?ӂ��ق�bȧy8r躙��SS>4�1��/�ă�!�,uo'dsb�:{�X�Ӹ�+ x^PvK�``E338 ��}a�0j�Z���a	?������@�A����4��Kk���ˑ��Nu5�T�t�q�IY�ym���$�i�5fcLx����h�X�ѷ7ܝ'�5�O煰,��d�(F�@[���Gp��%� М`�#�~�؆�6�I��8�Z�8�$�[G7�������.���N4�����!�����V�^x����w���
F���bXa���`O��)����L���y�Yx���yp��U	����e����,l��$�"��0m�A`�������gǖ��
Tt�H��j����'�'�%����oW�됹�
Z����	l'ٮ����m�J�q{���iqD��V�x�5��������ROyG�MX��S��I�������[�;���a2��8v��'w��?����� ��I&���H�PM�jT2��(���p�}K%r�+GHdؒ���t<�[ة��{�(Sh��A��꾗�s���ДU�i�V]W�p�e�ciy�,M���K��S�ץ\q"��M�ڌ(���oQ�Nd/*�/�sb�M�o���:4�r��T� y�����t=M��fE�1!�"�2N�w���Z��N�:u��Rw �ԩS�N�:u�����~�j��鼗�r0���! �ٖUG�Y%m�avmf�r��	�� D�6�i��X���칈Io�[��g,h#G� kM���KU��S���b���� �/��À�ڰ,�J�n{'Ȗ�#�i�����D���3P�:� ��s����X� �]̶���*��q��\&���iBՏ�+�����f�g@�w�os}� ��? 
R��W���6�]iI�B*�q�z@�mj@���@�����spŜ&��+�
 �VC��[ 9s���Q�{���<µ��@v��hv��h������!-Xu�t׹�*��%�Z]G�h��­l(~MI���r>�7�~W�Wg��窺{�NG��-���s��#�>���]B���-F�C�}W�8���$���c�Aތ��.��s�(�O}�����Q���#�!�>���������
 ��3aX������������ ����ۿ�۸���`=: �d�aN)�?�SgN1��_�9��*i�����D)��t�Q�����my���0����+GL?/_B'��@��#�ŉGDq*� '@���x��):�%��ԶR�n,�6��7n�$�������͛7)���tU���:��A,)����'`�����~3�fG4�l�2f[�>D�NP�Oq_]�`���#pt�&�9,���el��S�"=`�}A��X����Wǹ��~���Π:ϱ`{�%�*��/g_֢��Uu�O�T�����_W�/Zt��^����S��f�_�}�,�P�jF���P��7p[�8�H�둠S�N�:���; t�ԩS�N�:u�� �u`k#�̀�6�hi��$�� A��`�%�Z��<%���*Z�������^��Y���Y]l�����e�%��Bm�RG��3����lC$p�.�@Κ������(�1ϡ�����u�ԭ�<��� �P�&-RL9f,}kcs�g/��}�Dc���8���a�k�8�<���L��B������T�z�˔9�pЦ�ιō��b��t�g���w�Lke!h5H.�Mߊ�{P��9�zK�^_���^o�u����m3u�d{�v^0�� �P]�hǶM�~^*Q���д[��	�V�Ҁ
�x�?�ቯj˒Vw��r�������;�w�,Xs�@ʎ�^���x�e��k�}�菆�ˤ�=Uf�Vk�̝��Q�8��VM����X����I�g��ȫ�y�[R��2(칷T�^���7�l��n��5�+_y^��7�f�������`cI�?��<�,t#����}|��������� �m�g�y���	x�;ށ���Ï<��ï���	���g��#�{�*����;ppx %�@�0�٧?��G!�l6I��a)��1f��#�F�K�:e+*s2���`��T7�=������GrX�=T$��Q��̑�%@�ѡ�h.\����0��0]CyfȤ���~GGG��T����"������S=P2-���[���nOC�Q��Vd����o�x���C�����C<�)�7�eX���*�w��'�O`5��\lN`7�?�G�u�N,��]�0��Ex��+���|7��o���ix�k^������y���5���M�F��-�n�u/�m@6��:�b�����|b�ȶ({���@Y��]��e���3o��QU��=kո�3/\sM6��Xw���_
�����F���m�u41r���F^=˙u�f�����?O�4W}&��lk����U�� �/���u�ԩ�ˊ���ԩS�N�:u���A%E�)Z�f#����|Nh�)v��j	�
|ve�j��8�J6c��5�Y��{;��"W��o�Z$�+Qv>U��� )g!5�%��Pѥ�+1�q�<'�{��o	i6y������3��sh�F#zP{����)��p���$�sZ~�s�5%w�Ƞ��"{10��S�3�ӄ�!���-VG�?a��e�F1?���[�ר�J�fT��hP=����\�3g�r��V5z m/_��ﭟ���>��E��,����`C���n���:��pt��gY���F�LC4=?NWGYH�d�W`j��R����y���qMo�1�����N�Yv��(��Y��+W =0cs�U��TyBͿ�&w��Mho���ļ?��\m�T�V�N�N��%��Y$,�Vd����f�l�nY*�Ҙ�W�O��C�Z����y� �,�5�g]ծ��o{�ѿ2[�*3~�~�:L��x�Ed��#���ː����i����א��Rx�A��]y��<z� ����iY�ȑ"S?��	��͸�[7oN���p|�F�S�ʌL����੷��D��G�{��{���	�lNa�Zå˗a���(�z� ����%�1Me߆4��ekPҵ$l\*����8�6=�9�P�T�*�3uD�Wd�nݦ���Ƒ�1F���m�5:H���[�
p~.�?����0�#�@G�Ē6��.�(���=��fL���R�usd�}��ś/N2ڠ�A�<T�) ��ʚ�����>���;0�?����'�~��N׆�'�|V��{���� �rlJ��c^�{=������������f���|�#��O��z������o�:ͧ��0%]4��n5�(� �`5ϲN�P]痪Rm�t29�h� ��ۮw��ui�����o{�W�^����2����>�:�δ6��"��{�l���]��������Y]�&���b��I�'���7��#rII��u(�S�N�^NԵ~�N�:u�ԩS�N ����3�~�	 ���@#��*(0+F;���/1�<B2&��(t5r	���U�+���!NA/~3$G��3�Um5㙏��&�\�[�QN
 � +�D�U(�/����M�3���A��O�����t�л�yc����23G�����"�7��4�\|�iՖ�?[����@��Nj����hD>� �6W��,8p��lR�R��p���&�lо:+3@�"��=�޵�3n�K������j�s���<tqR��f^t���w�ܳ3�}��<�k�J��C��~΋шXo`hqA�:'�6S�gMG<�l�
׬�m�Tu<�U��L0'�< P���94�,]��Q����I[�d'�@��ꮥ�K�e�A����JN7mϾ�PͳP�,�2F����e:TI�ܛ�B}��#^4�3f� ��d��pv�nŨ�t)XH
��#"�0����if �}����ʫ/�j��5e�s�|��M"��{ҩ�(��~�k�̗�����}pzr� ���	�|r��d{�!h��/�ח{%{�����n�S��$��L�]������/�/??���~�Uv�=C9�~u)���ed*�z\2����p����i�ϩ�mN12� ��i2�x�X� v[8,)��e<�-F�^�3��� 	�� �vp���xTA�ߔ������<�i|���?t	.^�@GL��/]�"�"��<�*�($�t��ۥ��X�l
$�@8p�;G71�8h쬧:KF�l��9Z�A�x������ptt�\�\�%�n;�sB�饒���'^yu�F�5�ɹc��֧���֧��]����]B�]x��n�x���q��?�ӑ���"��}�7M}��?��?�g�}�x�*��'��s_��,�n���X^�j���Hwi�m�lֳ��L?�`wŁ����������u�[�M���5N��u�T`��q�d�Y����	�--��eO�:��i�W������&g���`��Eb��Q����ǟ�&M���>�����aA>�	O�Z��o���dh~w�ԩS��s� �:u�ԩS�N�:=xB�'��C^�hfo��+�((DFo�3S�g��0��lx��~l�G�D�
�ݺ���@P�&���j��v@�'q���J9Αa/S�϶i�3G��ϑqr.W����uh`��4"p㍵��b뽍ӷ��i�u>��ٞs[=��������UMC�E�5}������9zb_q��T�_=����k����*���jZf�]!��J��Ze����d�~����ۍ��97/z��9#y,ýN�f�A����Z$��,jw-H[������9�)�����Vq���9 4m�*q��u�Au��:�� �`8ݵӝ�Ǯx����3I���C�JK�GXq���Ӈ�W��Jv��᪌�O�3+�M/.���
�q ��*���.�$���"ǋ�Z��f�v�'��!7�[w���A@�,Q���~�0b~L=~���+��Kt_��`58<w�g��%
=�z<�X��E��xh����,�9�''��,��~��ٕ4�������V�w����O��� <t�
�?03@.Q�@Y�
O/\�	������˿�� �?==��0;@B/F��w�h_���xjӋ�+i�KF�����n�D�SD��7� ���Ͽ�YR��/u��.�[��ǌ��<��;<F biE�#<��#��K�<s��c
 ��n�ͷ&^_x�9(�y��8X �'w���0�S+��I�;�w�o߆�w������V��/^���U�������8-�L[��C��N��G,�8JlY���w�ȀYB�r�������� ��E��so|��UW�b�%K�����'�|nߺ.^p[�>�/t��nzE�n8�&
��6�I�f�l��lu����lɱ1��V�����L��9�û>���a�����)[��j�v���� ���,�<j����%8B��$��{�r;�G`n�&���k�U�ԩS�Nu�N�:u�ԩS�N�@�H7��)_����DķT�M	�� j]b �:I�F*�Yk0C�E^*3�l��ހ了j��6�%6�y�$g��Y�k-��g�2��3�YFT ʷ�!mC�S��)6�:��GR�z#�3&3����UY����ߜ1���g����Φ}��kKF酺�!d��a�~��to�ޏ�|�K�dwo���_�K�-����ܻ
��+d�qg�W�[��U�y��:9p�j�gecLƸ+��:�v��:7/�+p'S�!��=2g,�:mjA҅gΜ�&"9Z�#C\L��>{���e:��n-���"	�l%�˻�Z���*SJnu�O/�ސ>ׂ���&f�(N#�H��s�c��p�3�n��cU�¼N�sq�1e�����R�M��!�>�	���
b4�v�� �>�F�KvP=F�l��?�gp��E�h��8��k�l鈒�~X���x��+���K���~�\���:߾}׮]�;�O0�}CIOv��M�Oi�p���J[v�"�>�����|��p��%8XG؞n�k�Aڍ؞�n��qE���Sħ>�'��?��x��j��W_9�r�?�XS���ݒ�`s|
���։�m�8;�l����bwz��	�ố����U,���a��6�����O�}���A��m*�nC��x�I(��z��x<tr���?����{.�� w�����wN`s���i���i(�����Mx���ԦHr�����NY�&í��a3�����S9��x9�S����� n�<�Ͽ _��_LϿ O���U#Y��Κ|�:�Z=d�'7�ax/�ݻ�{���{������ۦ� �#��w�~��u�9zYa>;��j����4�RK��ۊ���纳��%����r-/��@����ԩS�N_�� :u�ԩS�N�:uz@	S����R�GLoJd��m��Ef2�MA&��Hp}�}V� (�0f�5�HQ�j!z���1φ�`�{�V4.%9�td�^nb�������i��o#�Z�d2�k�:01T2o�����[dV��G�@v�ý)�c�^]B���%��j��.]��^E{e��h����L�<�٦�{q�����t�������T��tSS�p?�3{����bp��xm@M_z2�	���y�[�2�����+f��({6�E����h4x�Bݧ�.�n��[9KL�/ǦT'�
MXB�Q�,d�i߂	|,(�Āp��u�8-7zV���d>OFǆͥ�C
aU(r�H��5eI�P��)�0�
H�"|�D�hj�Zoit8�0��k�ό�^%d��A���!�o_�>W',���X��I�N�9�ޝ�܃
��r��w�|���wg��z=����g��6�5�ve���*�]�1�>�f�.�X�z�3���P��������"���o6[���P�s�(����pzr���ҹ�<o˯�Ag��	š ϼ/1`���8�9z�D�pzC�s�f.G�T�۩����� ��>l'�����n�ɿ�����)	3��L�����y���?�/�Cg��!���1F�N?h�@�w*YN�(�Lg `���'ð
�ӣ�ŧ��/�E��7�E�ow��w�_���ӻX�0w�����Ο��Ms�tzW�������s��pz�̏R�W�5@�F�C:�� F�Iɐ�n�xNљa�q�{��޲_��?����0Le��8(ۍ�����T�`(����.��
��,�fe�Ǝ�Ks﬙�rM��9r��d�_�W��������2��҅5ъ��3�t��yp�s0ۖ�c�^�����}-���eAヲC?�4-��e�g�#��1�Ӛ\��,��O��%	\
�Xǭ��v�}Cʔm�S�N�:��; t�ԩS�N�:u�� R�R�ؓ�@!1ˉA,����gR蹀�����`�S��� c��46; ��]��

�����b�gb��/J]Jk`K'� =Z���d��3"�fN"�<�+�Yژ� ���l�s}P�����<Je��ě�IZF`#��ܴσJ�6Rz6�1&��O�fi�kr�����Xn���Y��貳��uv�tuYg�4���g)���%���usgڙ���@�E��fH�3���o��%��OX�H���2g���lt^"�*e�}�P&�=2�9 V��R6���'�Vθ���;T��c�rMp�y���Iڌg�[V����������}Ƣ�ܱ��5���q��7��M��� l��]�`��N�;d �{ �V�&��6�ɨ�W��d���11�]��0�45�U;��X�T���T뉼���΢���{dtV1�zs�ݕ��们���v8^�n����/��#Gn��cĹ�%P>g�H�����Wv�h����%�{����P�QW/�/�$j>eIُe'��둑�]����8�c��8� 9'a����^�S�d3��;���T�fz>F��[��^)2�
���nFt(�G��n�2C�3���f+�t���_":C�]B9������/б@s=dr�*G���"ǐv6�w�TQt�80*�"�J�l���;z������O�W@b9�c꿌Y��������5�k���4��/��$��:�L�˽"{jE����2�ub���1]ݗ7ta��w����s{V����X�U*q��8B��o׊�q_���6��ޫ:fk�w!�;�%�fsqr��2�(��o"�{���PN�,���qW�u�t]�x�-�勃&�d�N:җ:u�ԩ�ˏ�@�N�:u�ԩS�N(p�Ǌa�e�� #ǂŲ��1�#l�����4�"���RW&#q���#˘<@�+��MFq�Ej�3��K>��sV��&M�_��@�%�a_D���lp7����9*�׹ ���(�BZb-��t����|�o�V��ڞ��c�$�+æ�i|i*pg�>/P4;��EQ�#�Kg�YC��R���Z��>1�Ua�a�t,�����4H���	����K��/���z�a�[� n�-U�:�2�*r���������FS�]3��Ԝ�{&�9��9+�O�:�D�
x.�����H���c/����(�GE;�=���2�e�J���Y ���M2�������ܸ�:O���I\<��C��x��@��.�ʯ�ݯs�ӁKZ�t��0+������Ks݃v �T+��Nt���G���p}�ĸ;�Zjq���{�t��G^
�e��u��<SL�8� ��[�vm��Bխ�d(;���\�0�d
�K.�cW�Dq(�ӵ��+ �8�����,%�����{
E�>Ԣ���t?��O��Rr�wps�X�v$)���d9�ިD�G���
���� c&Ny�P�����f���eWP���x��9?p�(�;�1�.����.A�����x�"Yg�v�A۞ƌ�]v��8�_J��}�l�`��ё��-�(s��m��T�9)б
��$��ƞt�8oy��w�'*;�{��a��W��]���%^������6�3��N�-�{�_���-��k�(�����扖���)����r�9�̝4 �V2�@�=QL�Ȏn���:u����E��S�N�:u�ԩS���0�<�UCH�8�)Y�L���#�fv�
ڏ @H2�j*ln4"�#�Q��.�*F�F��W>��b��~�{h!�
XC`�g6 6�6�I�z?����s���Rtt�h=1�Fp(�H S�5kw�Qt'�� `���od'���!KFO5;��"[��`�do*�l/�wnC�R�'����}5 G3�ث�9C=z��$]��1����Q4#�`}&�Hd0�_����r���Wy�ƅ�2֛��J���?W�V���u~���nG��h�ժxg#�Ԥwy��20,�~���4� �����6�`Q�����|�W�Q"c�j��w�J;��j�W�m�����s��������	���q��x�4,�Ug��C0!�9������-�+�bm�\��P���^�@��?�9����{5>���a��[0�%���3+��V�8���
lN�����wʐ���2-�rIS����C���6�z�/!�n�����/��RX��=k($�uD�� �!��N�6;h�T���ʑsꃮi�G;�|�s%����8+~�X�����`�e�'��	HX�g�?U;ܼ�}�:�,�]����T�K�@k�v���0r�}��f��xK��	�w�甈��(r�a=�#���89�_��*��������(���z$v:�� �`�24�(ٛ 2�4rq	�O��k�\�gȔ��.dN��k��E��e���Y2�o{�ӝ������J��^��6`٩hl��I������P�5�}�Ο��C���J0~�}`�~ʵ�����{R�RP�@�� <��B��i��d^���z`iN=��7�r�8e���i}�/N8TDVYVg(�N�:u��uG��S�N�:u�ԩS���D!�<��3XT��h��`^�DB�ͺ'lم�9��R�bT��&
��}�[�p-��Y�o[/�3�լ���H�L���!5�g��� ������ >B� )��cA�-Qnf��Y��LQ�K����k��R-��Fg����6�;9H9&v6\4~e�d���Q�iy���6�>nǊO9;�	�QWe�~<d�g��3�{c� 
"���<��Z|}��z�	o���/���fwLC��^�����=�9yF��r��ɠ:%x���(3XW�C[��7�l�Ǒ���	M*��Q�
�.i�EV��H#� �Է�w��T�W��-юG����k��¾{���L� �tAR���79���E��ܗ��X�6�ˢ�O���W�)��� *ǔ�����0�9aP2�՚�����j�-��
�v�UA�#9�l^�N!~�V<}��(��Y�����:y|jt1G���k3�若L�j���S+���U/j��­����>����F�����A�{���בEI�箆�b�hm��z�� {,��*Y��[߼��z*��G�z_��<f�?�ڵ-���8z�"�m�4 ��V���N�eP�L��\���1t:��5=?R�3�E�#��(��"axw̩ifuv�%�!ߠ㛺:+@��&9Vk�6����8>�=0п��O�~��w1�c 9 �kL������@��)�1M��j��C{/��:��'j�_�*U���k��U�� ��S��׳������&�y����uپ�<Q5��5+�2@>����CY�R9>B�x�1�
]PP&e�뎜*ٴr����hrhزswAu�ԩS��� �:u�ԩS�N�:=`T���8SbB�\���eI��)�Ƥ`A��0�d�`@Y�ј)&Ӑ���u9����I���~�����T-9��X.O@��L[����3G���B,)5B�l�h/1�a-
D��Έ���<�����j�f��Ȗ������#�Co�3cc%S���T-�^M�G�9�|Mb�Od�hBJ�Ij�oZ�qj�GQpy���K�=�ހiH&����U�め׿�`(0P��\r��A�:� ?�/I�+@�*��L��D�Q��9��-�?��E62���Y�m��+�V�ƨ�3ͺP��#������,0���x��2��6�$YpB�u�q�
d1�sz|�(�a}lN$�츋u.(W3]H].@H����RD#�ō�wD�������ED�mk`E�5@�F["�Y�܁
(K�����o�R�c�(x��,LH*��8@G�fW��1�Ftw�|#���@YI��Y����.9+����k���7@���L�L$����#^�������̯
	�O�K]���6�j%.�r�D��Ц<oC�4Ugiٶ��֣�g�N�'�i��;3����Q��({�Ds��lO@�9�%Ʋ'�9y_���mC�sCjOz3�n�~$��~�S�#��\H������4�����
��^��� ��N ��d.&�9~�H���Ɣݚ(�Ӝ��1&kg�= ��	$7���>X��5N�D���1D��({�ȼ���؆�:z�S�ڴhz�j`�IB��g>kUβ����2�����Y��e;��2N�a�����Z�㸩X��̫q~�g��s��`��rS/�gXQg;��${!�w�8Yd7᣶�����u�;��3�H)�?��'��mFgE>��v�Ui��=�m	�)ȟ���F�ֈ�-,�鯻T��&�.��S���4n�jEG_�#`q(�hy�ީS�N��N�; t�ԩS�N�:u�� R^keIy�E$#���r���4��T5���f�UK��DjH��f�l�r��`�`��}1��Q]J�.��a�3��� l�(/e"�cQr�T ��A	v����Ԝ]R}vv>]�����l���(�Z�^F �B���9+�1 z�L���gE��'b���-���}��*d�ա6�ֆ�6�q?�M���i�!޳�!���D$`��lIri���25ո<�����֘fu��l�N�%�a��3�~.�^���g���6���C=6@�<Z˜�S
:�d�Wsǵ���v�bb%_�5��i���}բ�4�R�3�?�  �ͺ���90�!�Hm��``L#�9(�\^m��X����f$�3�0�ljF�,~� ��)"@��$�S��9�IuZT������Xg��\rl�ϙC��jy���\3mr}�Yd%���m:,���2b�\�N�s�U�'}�u`����"7Tk�q0o���ڭ8]&=��u���@�Wè�1���4�;�'������m�Po;�B{I��HS稙��gbU���xM��E�g�W���5%�.��x�.���{ءL�%+Sf�[~�������B�Y��1�l��D:�gk����e� ��1����by7-<��[�n��q4:`^���Ź@���m��
|5SU���V�O!��#�b�uM����eM�Z4������@�}���m	�d�62��e�=���ty}�_�w�y���Pl� ������z��_�w>�=�����H���q�����G���7b�۬�e��`e��]��`r�'���g�m�4-궁�l����8��>�&�{k���9*$�8��>aڟ(����r=�:u�ԩ�˅�@�N�:u�ԩS�N"m#����X4�&4nf�^ڕ&��@�)�&T��b=��`���{J�:����W��w��7W��%����l@KUh1ގV���P��z�3~�љ9ZFo`��l�����M
f4� ~�y�@Թa��K����g��٨]5N-r-|t�25=����%U� ����� �X��
�������Ƴ�������QQ���Z	�O��9K�@fO�Nl�t�� ��j�Up��������3��Q��l���w���)i
W�7���!f���z�h�n 4���傍Վ+���52 E��p5 ��q�f�H<�p��
�W]�r�A囙�(�(*���Yy��(]Ɇ���{j�Ĳ�hq
�)�&"�t�z9�����!�@�C��9�inf�{ �i�� p];��pq`�M���材L�6v-SpfC�4vrfJ��/ǔ���G�X�YAV{��,���U2��˴�/�K�S��3bH���|��,�X����)w%Wu�	S�1W}��<�5N���``, ÓYc4jA�ޣy�,9Gc�[�	��yt��v{�X������ڼr2�Gp��y=6#�&\���j_Ї����s�u���c�({�8G�2��ǭ���#q"����X?&�� ��Q�Ǎ�ڙ.xg��p\_W��E&���%jYYĽ�x�e�����"�~1g7�x.�\��e��:���$����2��,m�� �C�ÔM�Up��OR�>�y���u���) [����l��S.�����jc}�=$�Pe���D�������A>S�����H�yM�F�&jJ��3�^�9�i��"�T�e��X�c(,NN�ޑ�MǓۋ �A��E�����mV�ߍ_Ǳ̛j.:����B��n�.s��h���N�ۍ,��:=$J���~�C�N�:uz�Pw �ԩS�N�:u����ՊOE�H��㎌�i��g��$!��s�����
 ��S�o����g0�7{C����!vY� �fu�yhdn�������`�P��[&�r1�+Ɍ�)Yw2,�QX��hG3��g��6�XA;aH��� +�ȑ�z{�V<�Lj"E6�X�6��[���[+{���wv � ���\,������h9�|:%��3�K��*
ƍ�i3�F8���2=�t�p=V^b ��ؚE����]&Z�4���|6c��%}���z��!��f��n*���F��d zn�!�|Ku��C'���R�C��L�9f��l��[._S	�J�y��WiQ��$#֏	�W����\f��Am����[���KT(h�>���	��.�5hd�|�A��8AEI搠2$�1�����t�; z_�ŨV���ze�`�-�>�t� J�R xj���59]-q���y�~s�h\�+�N��K�%���YF�?�ңk��� κZz���*��دPҬ ��	Y����Kˀ���ʏ�s�לҠo��B�E��ٴ����0�<��
_�s�R����!�?�����ДK�������X@cA�b��G{�R��vc|sV3�є���TJ��t <��FT����qb�Yٷ��qgQ��ݢ�C5X��h˃�qs��Jl�qsGOQ` Tem.���{5�S����(�dw��ˑy&��W� ��ݸq��+�s���0��b�c�x�̎�Ղ.�~�َԒ}�_z��0�����J����ӳ5�x���^v{ �􄌥����e�=K{dC�3p5g��Z�Y"l�g��Q��W�v@`gP�֡r��G�X���}��@w<T�s�m^q|�]��)s'����:���	���}�ևv�N���RD�+��׌�7�7=@�N�:�ܨ; t�ԩS�N�:u��Q����`7DخW�81���R1F�[�3J#�Y�-���D��j�Cs)�\zN��L7�VO�������J�s����܀dZ���Z��o1t	�"��X��7A���q3�Wg���MI�*�b�����1�&���*gl
���f?W�MeA�ݝ20���A�Z�FJ�UN@���� �K����E�e�ɘKb3c&d;w���w��׺km\� �+������d����R�C��� �hhs]E��:nt<��ء�  @��y[j[�?���`�Šn)����}�GW�l��l��L���ұ��12L���`�HNƬF/:p�RKs=QT����R�z��M���y2c}ʭ{FQ,QہѯXoT��[ �*g�N��	wi�W QX0���	,eÑh�`�̳��L�'�i#dl�|��a�y�ۂ��ndYgu_ Q��]�10�#	e�7��`� ���dT/�mu������T��]d�k������;���ʷWC����1T��I��n�V.]繮e�h�G�>{p���g`'���nr��!9���2}Ү'*O���� }��S�{w	8�dS-�L�^���SZ3�m����	��K�N�S#�;�0�ڥ~�W����$�{|�������@G&��I���>��K43;�qd�
��v֍	ӿ���9������MJ�@4���ߑM"��B K�º���/���������W�i��@��%ST��V��z�d9(j=%i;��H�v�D� ���M.�_{w�#��.�Ş�e��'v�(?�/����%H �'H���cM��f}�g$�d;���c�3��7�E�޷��6=�rn�)ak�j�\�et���)�out^��9km�d�%.�ml�}Ԟ������}9�K8�㖱����O�s[�zq,�ϯ�V��;�[K���Z ?�ڤ�oh�ǲ�ؓ��r|�!=�����?�gm�מ�S_�5&�^K <�������^~�e|V�Iq��
K{6��6�Jп������z�ļ��9f؟P�n˼�#i��rRZ�bM�=ip���^ɤm;���n[ָmO�v�����  �qH   �ߙ����w_����OaY�_�O����_|��~yX��{�����<]��a�4ކ��e)��.�4�����f[�=���g�^�[��5�>o|�p-�<6��Ê�Ƹ!x��W���kCg�M:�'�>BQw� H�*�?�=q����u����iδ}q�b[����hWZ�����^Q�;�����{�6_��16>�i�0�w�5�J�x����z	y(����OВ�DzP�n<w���.�G5���ӯ����S�&����[����y^�P�-xt���z[�0,u��7Ze`���cMs�*ĵ�Z�K��ZOq]�]"A���s�ekD�W-,5�Tv,���c��B�A]��{��}��_?1\����@�%��tq�e=���=�{H���kt��u�Zc�֠K������L)xU�u�X�����u���J��X��>�~l�k_ͼ��@ޮ�\>�Yj}��ڣ���n�����+���)�X��|Jۿ��NK+�$�\�P[�cMa7���m��aM���}�ž��õ�;���]��TYGڇ!�2��Չ�(th;q����1�'����@LX/CP3O����kviǮ�1��0�k��>m��aX�%�2�r��U^�1�C}C������H
{��ʺZ�x�����q?s�i�ό��ٴ�9(�y��� o͞{���_��{��@�Y�[�0���2|6��2����Z}Z>:�m�κ���!>���M؇�D@n%����!��K�R.�XF^��k��^�+Koݭ��pĆ����|(���R�?�;�oZ�p�]�{����vN���}a�}��y���~���Z'������qK[�B���ن�_�=�T"B>�C:�Ro��O���r�y
���ɑ���o[^N=�u��\���Q�`��'�:�����i�z�����1l������$��HF�<�z����eo5	�%����xm�YO��ך�\o���X�cu�~����-Q�6'`X��F�g�~m�zc��}�;�x����my��:��R�w�'��׽���o�JK����:)�����ԝ[)�Բ:˔��<ڽx|��R�abK4��&��|��R��F���c5<.�>����l��R��5�G�[���Wo���	��]��zl�C;5 �H   �ߑ#
�����x�q}�|��۷߭���e����X�޿���������)����17D�q��[M�%��dh��Q�|�?o�{՗)������'�(@��ueʴ��-��U/���י�U�����sP���yca(�=�!Q��vc=o����<���>4���P��5��@YL��# r>d��4��m۾����K;m)�U<mh㺨K	R�9 ����RLC	�祝5-'�F�zZ�l���sP�S���-���������e����aՇ^iCD ��bޗ#��?<��9�I�5S��A������~�kС����?����d��릗�#�<&܌�[���$c?qð�{�'��8�ӱ��<�u�bxW.�A�S`�������̫��tK.8Fۈ���A��j�>횷;��ｮ�0��k*��e7�ZbHߟ�O�p�rP ��VOf=G��\��4���<�1�y
 ��҂7�4�H%%�a(�>w���`��z�,��n��zm�ס�/���ݰau�\��c6��>���͵ܽ8H�z�m޷��t��d��`zRN��&JՑz�&�W��4�v�=��5��`L��bh�_:�K���(��\���\z���m���������.yd�-m1���Gj�UC?iպ����$�Op]O=���=���wa�,��kYDm/-���r>ԃ�@��:m���J�l��|�v��˽�3�����{�_���J��Nh��h�l�IU��GZ	���Ї<���S�h�2��R�.��]J1
���Sݪ�P���k�Rl���t<B)S��E��\4�؞�2�~���.��z+���Rꏥ$�E�-7�sV�]����9˲�{{a`m�m%!���Zޕ�\������v�}���e;r�W��^Wž�m9�e{�2��6��ے�0�1%�\�C(ur�����g퐍Ay�o:K����Xni�$��د�|�j2�x�/�␃�|Ժ*�׳���JI��@,��!'D/�n[N���6fD���;ZU_MT�O�������޲<٪޿��4�U��%�����<����5I%��}>����qe�������ƿ������S����ix�`z   �w�����oÏo���e}��o�|����������?��������=�����e�n�轼�Bbz+���=~��MC�@	��H�RB��5V;��F�Sp,�|ܞ�C�d��s�ae�����S�`{�5���e�%�w?�@ߘso�gM_5����Al�e�C��%�u�M,����GG�ڳ.�8T\�")P���R������cZ߾]{���}���([NCn�Ǣ��6N���@A	&<�p^J0��P��CoθA�҄96 ������m��kJ@��p+�=^By}�P�J�h������Ѽ���,ʍ�)PWZ�CiL�m��ڳs_�SP`���v-���rYj��H}�>��S}ia��{L^Ʀ�Pz�!��
�so��z���[����k�r͔�s�1��-���1�~���,����at�%�T[@a9(�����um!�ei�e��{��{O:�>�i�ӻt��ܯ�����wl�49��Z�?�.���/�ġc�c���^h2ϻ�� M�~�{1�������a�a�8�|_�#;�=��/u�����q��=������*�^ʘ)���>Mww?8mV=��0�?�>�4̛
��hK�jJ��)�!��'k^����k*�e��eiw�Z�k��:zE.=�_�#}J�8�V����>M}�y��a=���@Ժ��]�h?�o�^>h[^mأ��!֠�~]χ���!�߿.A�v�3�{��6�R� �|�ݶ!�]������V�=����~��6�N٦��=�����2����`1Q<߼�z����$ʣ����"�Jl�?�����i{>:B��?.�-�`�/��t�~���Z��%�-�@g��&4�}���%��M{�@�S�oڻ#�"^σB����"_ʡ܇�b��=���iH�I����z��5]Rǽ�>g���r%�{��2JB)��AR�^�v���A��%9�)�>g����h\K}�G*9l�ɞ��/GK1�Z��c�m�B)�J�R�kh��چ�xm�밎��<k{�����WýlX�q(���Ӿ�2����a�r�C����W�����"�Q���b��Y�㏔��Y��r{^���\�?�������������?������_^�Y^��0!	   ��s��_���o����?��ÿ�駿�����ޯ��w���Z���{܎�j�<F�G��h�ZCn}
�����F��5�!��ڊ���9ғ��̭Zyx�u�o�;~?^A��A<Ǆzkpc3]�|X?�^z����%h��4uj�{�`�c;����%2�-sa��u�Q}�����^c��_3�Ɣ���K��t�2SL㶬k��������X�,�r�Q�#��;��v����k����n�y�����9Y�����咣�q�C�*��;�C��]+�:��������r�۪y}����_h-^Ch�ϫ4�k�=TV7k-�y��q���ƣ_c>�GI~B�eyL�^����ׇRP�0�a�O�ںl�/��ݻwC9+�*�8�:�����!jV����c�axSmۑ5�~�y8�z��L_A�#ؑ�!~:9�;�Ʊ����>�)'����m_�r1�WVH��k��!� 6�J��#�^��|��9��j^y�����˽P�Q_GR��s�y��F�!i$�򌡎-���bh��}Y��ao{�#���5l��9�6~��V�j�@(�x��#`V_�Q��L�c��0A����[�˭�w�n��1B�zYS�p�o������2dr
�H�#E�l��9�ȶ�WP��^�)�1�Tȉ/�5��LUR�YK@L�d��日��5��������K������$�øƽ��1�~�|lo�s�ǭ�x%�Qy��kK����1S/��i5�5}��WvZ~��g�8��R�X8�y<��vbz��w�܎e�#F�:�!���$�|NSh6��Zn�ŗ�-G�I��c�ZP��s���̝x,��g��y��y�׾����~c^rp-wx�/��7��u���9����^����'��]I��p.K	��a�SU\k�?��u���Z`:䵵ע���>�ܾ��\˰����|a�cu�.�p\�2r+kH��Tβc��Z*cO�y���AL�c봼YKM.�Sݵ=]����ѿ�,/?a�y�=�N�k�;b�eR4=��:I��J4띅C����td�Vʥ���:��7Q�Q�:a�3�����#�}����5��t��|M������\����2jAɯA�J.y$��q]��b�4�A�q��2�H��RD=�qR�뽼�a�Cާ^ַ�:��V���m�خ=��Ԓ0�۠���d)Ě�5$��_�.�{u�t����c�CK�=�~�,y�u���u]K.���k�X�#~�Rwk��s�ޞ�c{��Y��6�My�e*�{J���"s9)���{��m�"ڶ�Гl�y���ݗ��5����u����[�=2�z�!�+j5\ꑸ�~�[��Ǥ5���t�5#�����R��Vr���Ƕ��Z-�!?�ݎs<^����4�E>W��%��p�����].����������z������w?����9���o�������~x||���_��/�����nw�oo�Z$ �!H   �ߙ�v���o�Y��|��w�}��7�?<==��}�&\����	�,K|�[c�ev������5��9���Zc^�%�ǥa�}6�￫�4����������v<�ܷ���}����9���w/�s������ݺ_چ�n�Gĺ%��1����QC�v��0ϰ_����s��N��v��~�}vl?t�?���r��}�,��c����������=�/m�G�?�������Й�����:�Y�\�����i*�5�#� ������?���-�^:��i��o*8ow�̤�v�}���C>8�q"<98���=�OƷ{�������̼����4�gzѿ��Տ!�b������p��{�������g�����ܯ�~��?Ka��a;[���n//m�x�YW�Yj?�?d؞�$�g��~���ܔ���?ߗ�Nޗ>O��ٽ/���Q�{��T��:��Wէi?J������z�JQ���D�)�].�9ɥv����]���k)�-���/�TUǺ�a|�g�!��P맸�ܒ��w�_^F�K�R>�=��cr�3�����/����Ąl˸�W�3���k���qh�����/[z:���K��sZ�Hy	Ҿ�2�Y#��ߏSt�;p>�s
�z��>O�/��m�����e���͛z�����M��1�K�U �G   ��&S矧����������|��ߕ�ޝ���_������m0������C����h�Ŀ�2>������s���~k���g��������E�}�2>u�4����%��Z������_�^�ىa�o}j���n��ܣ>W���>w������������W��5�?������������E]�������%�����cˎ��K��S��ϖ���||�:��_���~���?�� �zMŏ��~�:,�14��۟c����W��?	   �;Up���O    ��&        &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &� E[:#�^�    IEND�B`�PK
     !M[��P�#  �#  /   images/62b25533-4940-4036-93a8-d94b028d26e9.png�PNG

   IHDR   d   H    �P   	pHYs  �  ��+  #�IDATx��|i�d�u�w�R�����޷��Y��q��!E��˱)�'FDĂ���aB��(��@8�,&6IS�djHS�����9K��{O��]{�����^ի��a�$��w���{߹��s�9߹���i��ҧ��ҧ�Œv�o?�.#����
�n�B��8p�!�qda[�
y���&�|��7_;2W��B��I��˲Y�q�煛Ǐ�<�����ꂬG��g���8n;��Կ�U����m;���X�^�(|������}T^sb��O�'�h���0���눪�_��x{�����s���$�Z4�l����N�Ɲ��ZX�GQq�%����3j<���#�Q�m�5����D�{f9.{U���Eu� �!�d�W ��k�2��<�(.-�:�ELQ��(��*Lm`��n�����.ʰ��	W ���|-�G�R�|-���G����f[,j�J��V���YĨw������栍���vc����	�+�#)gê���ͺ����4Wy���N@Yd����n����n��&�T�@]�<!��^]~V���X�!~���;�����u�W��;[ZW��)�M�ا��_��*k�|y}�d��r>[DI��B��v׳����у/�m���8w�Й�*�.���a�ڪ����i{��ߒ�:7/�x�4xxf7�`fc�N��]W��Ԭ!	�_1�¾'��F�9r����oL��/���hk�@;� k���R3����ַ��}�ȩ�L:]Zu�v��Y�"5����G��S����" ��%�8�Ȉ��T4�'��a=*��s��zgqe��V�:�ޘrF�c�yҎ��z���١�_���Z�.�_(,�R4Vn��6[�	6�M�F@��)���h���ǩT\��+E�@��Y	�+�&�)m�k���ԋ7�<�5�5:����j� *�O&͂���ˮ.<�����\�0���>L�_D;I[��҅���$��⣛����h��4Gv��Į���pz�Z�L�:f��U놱�[M^�qE� ��-NÕ�_O�B�|�'H�S���d�yҳB��@,IL����WKF�PD}�6��Z}���]s
��ݱ�fO�k�X�TX���UC��j����@�SK����*���o�ݗ48e�H�¹;ҍ���B�&���,��n�I�5����������r,��,��򪦖�
R�
����-(p_!��X��>��"vI���0/��.nr��S��P^��*ؖ�1@���
�-U�44�@*����N���+�(_�}��%��Z�i�Y�`���C�*�u���b��䝼Zk�� 6Y!���)�2�=w�βY��J��K��iV�M�j4ݖu�Ը\�V%�BWLD�GTx�^Zm�]Ҭ#��� ht��eTM�Y�`������깣$������.�iW��h�V�� �9[�I��D�pH�l�#�o'i^TQgr����0��`mK���8v���?��-�p�z?�r����s7�e�U���GGx����Y�͸p���a'�HS���ܪ17W�F��I��o
W���MU7kCٵ>[;���P���\)����mYUѦV���R(�B���jH�Y�Ǧ���r�t���l{�lj���a4KG��nn�f���y���s�zܤ����!��I��Q�n�'L��DM�G�\���H�������V��f�l7�j�Ae�c,��'/9�Lێ�T:^|ӈ�M�ih'i�'�����q+ef�m8B2x�QcY��.|_�l<�j�����c��q��v�˹&ҽ�L[��g��iz�FW��� /���h��i˲e�|�'@��m{���v�������/����U�|�W
nw(��e�:7�sc\�C�%8_EߪSSf�G���s�L���T��1���E�&2�a��DN�����$�4[�Ϧ{}c墅��q�v(%��+�EL�~a�nO�ވ����.�ڐ���?���BOd����=�'Zg\s{��&��9f��d�]�����2�3�3�\7q��5)�=w'���'�$�G��0v �w�{��i�������1qb=CQ����E}�oWW�Z9�׼�d9h״j�z<ޛ�U����֫T��Q�ճ���%n��<(�x
=Wq��r�'�D�:��R��%fr@a\�;�~.G�J�<f�����4��!��ǳ�w_�ig�[�01з��Ŋ29��c��K�U� p��p烝Hs�w�B������GO��7D��S���)�K��� �f��ӗr��V�#d��$��"�H��t�7+�P�$d���a��m�,��/��D�̢���4��q?~u]! �ߕ���"��Đʄ�z�L���
���}�!�/(QY�����"��-Ұ̀�D��pT���,�%n4/wd�����R�{�F4�I�,0n˹�똻�'za�;t�/V�W����afS�~���F#�wo��I�4:�T�c7�z����oU	���I�-�}�@�ED�aJe͊���u$!�{��n�X!�3�؄-���`.�������0��Ꚛ-�*6I�*ު"H�%��h͎g��0"���JeŽ�=����p�|�E�m�W�X�H3����
�ܸ9��]:�|(-�R��3ټ��2*ʣz�.wd�Ud-���\��C�FY�ķ-"x�FE�4��ƾ�M��ZE2�m�=�uS򘾜�Ѥ`�J�����"�ua5P$sq��e���#1�~�&������.��J�D�i��Y��G��Z�Fo%R��֥	�w_J�=�H��E���̠�u��SY9bҽa�I�(�xJǮ��?.�h���Ų��Eh'y>�U�X���Qb�=���R�=�An��t�w<��L��	�����5M�}+.�q�:a��s�p�d$�?��;��ljx��%'�8S���'S�w�a+��%5���ɯ����1�F���-��3!�P~�|`��x�S�RV#���g�P�0	ª���=��ό���6�v���Im������j{HK�74�
�~Ԙ˂玧�g'Yl�y�k���О������:Pp$ZIe��gd�ǽg<�!��Y�ڮ ��rM�}D7� -�:X0l&؁���v�q���U�>u�Eh���MSܟT�}`�7�eR�wS�m��.2k#i����x���R�:,?��6 x�v�A���������햓�fx�α�����G�R��h`Z�4�nL�!e�'�Q��Gp,(�X���c����]3
����������e��cƛ�����>��F"=��l]Fm#T��2s˨(�����C��fŒx_��]W)�,M�U4�o�|�W�l�ڹM�l
sl3q,K>�L�)���67�l���MK^�y��7��M.��a�kn��5v����A�����9hsI/�:r��N}^hقV;p���b[�2�� �Y<ԉ���]��^G�]w���;�'1S�h�߂�j�ܱ��cV�1d_�A�9���'�d|r��wջf���!��0��wA&60���oἻ=��b{�����Tw!;�h�[:��1�3=�l*��v��~�͐wp<�m�� !��cg0���EcIU�<6u���v�v���k����u�f ;�v���!��D�r4�1$����b(Ҿ|}�$XIs[������&��>³Ϫ��w7_x���������X�k[�R��Bch��Y�C���<�Z,o���!Q���j�����3��nq�2ȏ�6�N����8N�#�����蓇��Ll"t�_��p ,�WТ����{�>�z^�Uj�?@C^�Q=KҶ�)��I}^TW��uh7��sj���u0�>�𝸼��HT4Ly�@����t�'��vR�tX�U�ׂ:9�DMw%PS(oo�����[h����Q�����JF\`
��n�lh@�^�2P����DD=�y���r��n�D�vms��P�p��X:<�i�dy��j�w����:�����k����;�C	0��̀]>��d4��jC���ˋ��"m�B��d��j�!g����9��-#�����Z�F�~�/M�;�Ztdq�o�����|�z'�5?%Z��Vk��T����쒐��)	�-�n�TE.��A���<5a6hٚ;������J'��i��ZD˻��=���
�uLN�D�0i���}��i�����7jt���tL�8��Ͷ+x��=�a�}Y���J�#��Ui�ǚ"���(��%yڢR�O��U[;Vsp�*`����������}m�#�s7��i�o1�r�F$vV��V��I�����(��84�Ԇ�^�j��+��dPc��p�*Z8���RB�x��!0Zf-6	�}M�Z,�q��X�Խ� <�����6�XO�ơ�� 2j��kPL���0Spg*<ĩ)�wl�I�[�z
K�(i�AƴR�ខ؟�e�u�zB��S"�̬-�s7.)�P�ﴖ���.u�ƿB��'w��j#��>:y��M���7P�;�����#i�҃��o��_��Y�\��sP&�Y��PNQP-OT�Jn9&�����`:�����r9�#b
�V��r��h�ʜ^l��h��pM#[����3�{�D�/�3F��~�����Ey���7�Q睰TJ�#���l����C��9���G�?\4��� K��f;�W�5e�'�\���mD��H?�&z���u\�l
%�M�ϓ�H wI�P~y�^����nn~�bd�o�Gr��5�rcJ�
��	���m>�����4Ymy�GB&d�`�(�h�ȗ�T��PbZK>BB�ڔ'��E���;�;�,�P5iZ�+%t��(ZL�D7�]�{:���Z+��x&%gV�m0�2�JY*�2��<Z+L���e��C�֨l�F��Z����p߃���W�+���w�[s#iG	QE%�7�d$W�HT�iI̷�-�]��	$���wA�"�2�b���.L�ʘU�x�����5�:!�.�𺱈�*�(R3Oj�x6���p4^�B
�/�n3�d5��BK�\��:�*೹~YE���\/GL��F���1m�'Zg�V����N�^V)��fhϔ2�U1���t��F�q���B$,-!���-o�k7R/;����/'�c�O~;�\����h��\c##Km/����W��<>DDќ�3�PM ��p�'�~�յ<�]Y@�c,���!9���!�馠����?ك���6Lt��̇�QI ֣��~�X�c��:�a�<�
�H���;�ޛ!Z6&�^@��^�gא_)������!jW/Ѣ|�n�*�Xe���9��|�-_���=5�wV��@jѮ�o�չ&�U�3$���Y���;b����:N����Ä�Ow�*�л4s�P���%��U�n�$Qf���:_<�x�ry�;�����ʛ?@G��<9����>��b	W�>��O}�=�r���?����"�!���đ#x��'p}n���x��g�����Lc��X��A��&M��#?����N]����x��E�a��c8���p���Jtbvi��Àw������9�T�W֦���b8=���b�x$ٞ@�V��*�j+Ο���-�[ˑ}��U+����ǽ̆����9)&��FA�h�ro���`��ލeu�H
�P
10��>���t�{�����`hpff恬���1��M�e���p��
��j��
���Y��JS�(��q�hH��E�\�d��
�,�2<��Q@9;5�lT��9�겉��'���P����"��G\�R�����1��f	%��*�%��m	��~�����k�~�;%��;j���� 6��c��Q�T����Ɯxʀ!���4 !	)`[�i����1��"�]>��~�71������K��/��
���%���0:>��/!�+�t�<�,�݈��o"���k2�߇�'OɃ5�ã8u�z���u��GЕ����Y�ol`���8u���5�±�'������GgN���rd�VN ��s�O,��Qu�Ӌ���f4���A�I��g7n�4}�*�a�:5=cW���X�k+��Cx U�t�k.IP�&�������73xk��t*���,))
�~�o���M�u6���Z��Lm����H��^����|HS1��Z�n����?��ypK�|�T,�s�P�[f����Mk���I�mcx�ӳ�M��aHFՏq���l$�I�V]3*lD"!���ىp3�(���!e���;59;��U���ŭr���WP�I�D�j;����k0}"�����Q�X�L�<ًӧ�cue�j����{nGOO(�}��^� �≅�,�F�݀�̥���l�T������2A�YW>dVy�#�qU#!EB!<������뗾�B��Br�P.�:��d�T���@&�4���S�?O�ç�����"U����EFH*J"�k�~���?�c�|"y��/P��dO"�Ç-..������*�7n`dd������CH�;q�=wcrz�P�2=��e��F�%0=5Iv�8������|^k�θ��gwz���
�
e69�,�>��(<���,<5��Ihd.������o�ɯY�_\��c��@Ac�HG�po6��P�|l9LdrD�Z���D�G��?�%�m���_�җ�_��	GB_��AƸr�Y�rI.�-/a}�LW����Ittv""D��C�������e2�A�)*�;�H��=��2-Er@�P���
šev�@��+7CiPu��,a��y,MM��6�I�DE!���d+��¿���D<NL�O�'�{��9;:XO��@ht d�Եյ!�v�P���3�L�M��8�z��[�7����}{0u}?��x�CC��$�`�FA�&)�ߤ(Yw�{;.��@����[wG�5�{��=Ln�5��JC�K�\���w�H�<e+0?;I(.,W;:{Q%����g�ah�#T�Z��Y�\�Pt��'��śOD ��W��W_���=��!��c�'�'������L\��Y��*�����I�'q�℄��O���(��M�	������5���ߴ�A`7 ��Al�oHHvt�'��fA��]�"�r?"���o�q;E��F:�A�x?x�F�W�92{�w���ZEGG�S��S�(U�Xf(�L�Qկ ��ÛOD /��Lf�ў�ѧ��IbSFԐ��d,J����E��)��aU�6��H8�ɼ"g�,��q��V5-oGot��[�m��x>R$V����DB��E�r��.,,,�c��4	OCww�1#Ҵ)�&��'~;I�r7��º�3B:���E�+��R��q&�;y�쯸0R����c���d��Ar���o��wc��2]��!Ցt_�c�{zO?*��+z�T^�"z2�`���p�Cb����6�V��TM�� ����1VB".�0�r��\繉�TɈ��a#�f,��RH��[9��}_>�ԙJ�P��F��F|ʕ˕�J��^JHSF�^����SS*1��ip�×��U��s�7,�9���Q궻r'�|���&ĥ�0X���qd���-d`I>��˻,�E+���a]�#J��Y�	4�b�ݕ� f�hpP���>����_�Cwg�]	=FJ�X�{�-�L���)�-�����1f���g|�\*K�c�e6c�*^(r�t>KqJ����t�����p��y���!£�7�~��\�"!��&riR�Fm���*�w>R�1	�a5�';�T�"��V$�
y�����K�t�f�3���}V?u�LW�h��Lw�b�l8Bnu���HV��d����[�Qg�_�"38L�U��t��#x�'q��E<��%���3����I��M���L\��L��&��Rś"at$��)�3�U�.FN���_P~��r>�͗�>U��U�38Ї�=�E�X �]C�LS��}�@Ϸ�J����/r��~��"����u{~jK�m�r��vS_���E�l������b��;�S\�	,,�� ��M�1k8o&c�'Й����Lu#�Q�S#�T���u���#N�4/(�!ᲠH<����!E��F.�F/CX��Y�nʷ#�:���2�����"���7~�k��Mn�^-r�3�7����XLokA䖚���vX ����+&'����L���5�"�1��'��Hx�>�.]<OAa�/��BD/&�� E���+ٯHP\S���+͕k�ti֌pb�D`A���G湍u�:����ёq�~���~L�����o����׿}��w�Hoz����H+y�}i��n-��Ɔcl�`me+ˋ��:�-��2 �ƪrvב��Kd�Y���R��K�=	)ʣ&��$�2�:E��F�x�a���)�N��YQX�9FcE�ٍ�|�2�kY�\�rA
�$�6x��0�����ޑlG
�-����|�s�m���3W�uA���˘�=����w���|�Ě�B���^���˗��g�1]�rEB,�z��~]:~M�՚)��Sļ={o��kW0�G���U��^ʳ��?��✻��[xc����`�~�~�g�n�d�����Hؘ*F�����������[��mK�Z����
o�C8m98d�ůK�?��K��f�>qBL�y$?�\�p�|�&f�'�H$�[�9B����hw!O2���"�>?�tK	d��.$��k��,䋄�-9��q�|M�w���"��`���ߗ��cM���CQ�����6~�d�$@a���v�q�l��Z]Y��6%��%����kh�����l�BY]���}���b���g��-%���������͜w��A �9y���ȱM���H�1�����ށQ�?�oC(�{����V���*�$�fa���m��ͰYh.(H�#~.<����~�[��=�R�4}*�[.}*�[,}*�[,}*�[,}*�[,�@����    IEND�B`�PK
     !M[	��} } /   images/bbfae99c-8036-4c5e-89fd-a87441410720.png�PNG

   IHDR  �  �   ��ߊ   gAMA  ���a    cHRM  z&  ��  �   ��  u0  �`  :�  p��Q<   bKGD      �C�   	pHYs     ��   tIME�#Պ�  � IDATx���{�m[���Ƙs����8��GսU���袍�i�4��A�("�q�6'9�Dq��E�HEVd��HX�d���&�Н��g=��n�}����ךs��?Ɯs����{����f�J������k�5�x��p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8��}�𵂪 ʳwQʄRZ����k��{�Lǁ�%O�h	*T�J�`011@��#�QD
*B)�@ FI�"4"L�Db4��L[�>T	
4AU0����11��*��J���N�L� ��m��l@�(`\m.@aW��7W�G�|������%���<�Ç?���p8��h��@K�J���s�H��K���EFi��_j��R�kh�,A	P@	`   �jQb���!f(PA�U{�B8��W? � �FE}E��z�T�0b��P�t�>��1�yPr�P)[��7���I�����>P�+��T�hT ��ۻL���J��ui� ��5%Nd?#��z�vH
U�w�[��}��rV)R�""�%' ��f�v�U!�bs�!lJ���x�/.��Σ�~�S�����G����7 xD������%b~�]  A�=��~l�,!	"bz���
�*�E �
$S�
t�Nb�Z�L�WaEM����DՀ�Ĭ
�h�AU���!7�(���?��˯���1(��a��%�۽�����]���$���}i8���U�5�ժ��T�[T�GE�C-�J��eC�����	d�VE�RM��F���dQ�liO~M�?'0�w^d^�b�Op�x<��L�$����3x� T"��q���/@%B���w���w��ڄ����k��3o������k�q����:Eӯӳ� e�n|�Z��	U�M"�7h�Yr��((W���� D��@U�����y��䟽��� �6� ���X��D%"H�T�(�R��0+���	|KLO�x��8L����m.��>��m.@aa�]�%����P��/  �Sm/�J��eM�7h.�SD��J�$_+t�RM��
 ن^X�f��@�aJ��QS�t��k��纽o>c8y�l�BqĻx<������{MH��sF����J�v�������U�v�+��K�������]^\��^��������ԟ��|�^�/�-�p����; t�0�>]=����_.���FD�[%���P�)	R
b�K)PUÀq� ̦���2���_�+t�;������2{��W�~N�D�DF���k��q( �fB8�g���90��2�d�����q��o}a�X	�@�>�G�ᗍ�VU����n�./��'�����/%�n���Z�K*%��Pɦ�T d�ά��H��Du�Z�9��yeӕ�����}N�]�v�W-�~��;?��c|���	s)(���QJA�fB�C`036�`6q��F��,��j�@�.�q�}�_o��v�y�~���g��W~Ƌ��Ǉ��q�`ڿ�_�o~��-������<�Β�o�o��V�|����D2��\!���!F\]_#�(Q�W�Y7ƽ˧3]oqǕ�\`S���"ZM"�� J�jTM1+���y����M`��P���ϙ�gƟ��~�Ke�q�1^\!��1��,���;�������/b�]�����U��HI�Z2 ��"	���`^yۨ�j���l&��mH:��@��l�
^P]���u�{	@��9��s��{<��s�7��.���L@��i��%c��؍6���1b�<b�#��E�0�+l����U�_�������b|�_n���7^^���, "���~����g~�G_�2��W����O�����%�v��7�i��|8n��[���R@*��PJC��`�!9���E��^z�U쮯�(��RU����� p� )�z�5���5ki_2����&�5���5�Ye.1WEO�����9
�'����e~������3������1ݾ��}�������o����!����?��9�.��T��9���I�"')�
�慢�B{�g�Z{�^IU��mt�Y�8��ieٮ����$��qԮ�0Q���.~a�9|*���ÌL���9�((#cF�P��BDĆFly����.�<`Ѐ�p��Kx��|}��[����/�~���T�O@)������W�������~�ǿ��y��/a�yʘ��b�]���o�Ͼ��2r�~��p��3,����4�P) ./v�$ bLsƓ�^z��x�ʫ��
� "���ӅA<�t����<���])U��kH��Wy��P��]��� �r��G��C�U�/J?�!�(��#���,o�M���#���#��p}�����u�П���|�G�|���������e��_�|+��*�Z��BHU��(t�ͧg}	yK���*3
�U](y%@hM߯��@���a�y��`��s����N_�8�@IAA���`F �!�b�
��1�6<"P t�J@���p�勏��W�`xTv���8?I<��ƿ�H���4��.��C   �7��+��4�i�p�x�xx<D
�:�ߖ�߭i��A��8o���� � �3��Md�H���#��9g�./����g�N	�^~��������Č@=Q�z�I��;:_���LV6�^�l��H���_׾6	�<vQ q�P��@���Y���q�� �o�D7x�c����@�P���/�*��A_�����폐����_�^�����Ayz�� � �J�h�V���c��S�w�Vν~I5!�)t�j�/%]š� 뤸��P���x=@B"��%Ct��@Q2��j�H1�Z��JI#2fd8!% `@�� 	!d��������F��:��?����R/�t�{C�o���6=~��v��o�~�qw����AU�RP��Bd�p�:s)�ó�?V4��9�ߍi���p��·m)�I��{H:@JB �%�'H�(iF>�Q�H4(�>�@cA�	�M7�i��;()D �%oz����q�9t�:W�dg�o�;��#����u��I�%�X�a���|����(�߮y�#!���@o}���8~vs���[_�N
��~$�}�y��޲,� �Q*��9�%��kXӀ2A҄��4�z�P���oYY����aJ�E�*��j_�*�cYXk�PN��l-(/4;��.�S*7����S�����	��IZ
� H�H�.� K-��"
5�d0�6؅+\�x�W.���xix	�0"`Ѡa��4���g���e��2���x��p����-!����n��K�u����9��3 �����͗���o�*2��O�\~_��o���O�i��N��y"�3Ho�Z 2!�#JN`"��9!��r�0�nn )!��8D��r��E@q���5~�۰���FFV3#R0Yc���Q�.DW��ޛĉ�~��P3	j��6��*s{ͪ���O�u�y�T�����UM�0(�X
�'a:��C�i�ݏ�{|����Ȓp������/	_W��/}�!l>���(�Z��-��D'@Dg�(D$��I�\��%�-h�Ӿ_|�U�v7Zy��1o��B������״}��;��"�ܴMȋ�iT�b B$�j�,�JBT�[J�A�X���B� �غ �H ��`@)B�6(��3o��4��4 �	�kL�c�O��g���8�0��s�Ͱ�~i������w1lw��t-����@��m�$�9���M<|囯5��۫W?6�~�j���K���U��n�O!�-�dYfhI�r��-E��	I,^.9!oq�y
��0n�u����3�4�c��ͣ�-bܘ�#��a�K�J��J�S���$�U�ng9��޳�R_T�9�h�EƂ�@�����OՒ�J�I9D����)㯕0��D�ߺ�<�����~������������O|�ʬ����O�ւ�Z��!�㿡e�(�)G�r�j2[���T�<s��qن�R�T;�Ψ*t���F��9��z�Z&'銢jT�4*���-���9��ւ�Y�]D@PD
�H%�&����Q�VC��H*�b�#Ka�]"�Lϰ��pF��~ʀ(
�y�&��M��7s���Y���t��1�� ~!����g_�t�3�C ¸�Ї��43�3���/�ٳ=��
WWeh���u0����#��̀�rP@b-}�j%A���BH�L@mX����D���Iָ���Z�X�K���jZ����1�}��p�b��`@IJ�A��AT0� Ί�2f�vD���q����Q��0E�t�c���
����v���}����;�y�%��j`���A����o��I_�"��>z=ݾ��*�E�'E��Z�5D8���h�C��	�@��|DIGS� H.ȹ@0�	ДQ�#�t � C���05���uw��"_? �&[T$K||�7�ӄ@������u�{��KoΏ9\����%/D��=����f_tN��;EJ�֛R7J_#�@uF)�e��{�O�����~����~�w~�w�����V���u��o��|���W�|��K�H���"G�L�2�lJ�%ͫn��1F��Ϊ
��w�yL��M����E)��z�ž6^O�:��׾�aU �Z"@�lB��;��,O�@����z!�$(J��ށ ���l���p0R�Ť���3bQ\L��-�����A� ��RB�v������5���������3S��8��"z�oso!�o�?�O?���q(1��%��f�tv"�w��T�Բk�a � J�s�a�q���	L#�iF�G�M3�:Z2r���<�������}��ʟ���G�q���D��2LE��FG�b�c`��B���L��	, )�M��`bb��Y��I ��H�tr��7�>½�
�����_R�U�Fji����P��
U"����V!�K��R]
E� n�b#��:�Ah�t�����p!P �����^������ 8>y��h
n�S� xh+�Q
�60C�~a�.�J�s�JB��g�o��}�f�g��]4b��� )�����/�9^
�Hy@�!��H�q���7��oW�߂r|]U^*%_�f�P�W�Vb�%��@�y�e>"�(ǣy���-e���'@b��%c:� D�4�e����!�@nn��gL9B9X)Z) ��oN��%�T��G�ÛR&��!��Xe�$��nғ�A+��.R�m�e���Ξ-�K��%�i3 c)lT�D@��H��)�''�o.����nz���O��#���a_+|���f-�a�0o����5_)�R�Ũ'�H-+SA˃T]�oQ�a���g�8M�X�jU�X�6ֹ-���s��2�kѩ
Z)�wR��G�؅["D�Ь(�0A� 6A�(g(B��g��#B�dU*`Q����)^C�
�hA��43��A�!��A�^�^"���{�BxF����D�%����ox� �q����ՌF��� r�0��N����N3�W��z���y `_��"����.
D>����d�"ø9��IidC�qP�AJ� �1�C��n�	1��R؍X�S�4A ��(TsE��*7�\5s���C��L꒮oZP�7�7T�/IAbJ]�i*UΩ�Y�(DETUE��Q��q��THJ	�E��,Y@9�EU���PJ�&*��"���T�\��-�˂�-Ƃq,�~�_�9�B�R����٫Z��*���l��r�^�3=��C�<�������`�hH�޽P�E�#��HyՇy��\i�;���9�ΐ־Y�'ת
J� �(%[-�<��#��M	�fS�R ()4%d�ӌ4O��0#猔R�P#�b�R��0����f�� sg8툩9�M�5[���Kύ& ���K�{}��$ԭ����ԍ�ƪ��ηváv�_=]��p�b� �d�I�oU%��w�VDE�n��2��ܼ�i\����zV��*�ӻ�'{�q�M���/i�sH�G(gh��V�V2���>���@��L�QSƴl�N�t^~��۷}JQ{]/1��Q�&�v���^N� ���M^[�f��FR�`l8��#v�E�2CHl�Q��I�d���I�zp�`��DDe	 &&��Tn��u�b@s���\KE2�L��  03�Ja$#��� V�P�C��8&���(4�(QS&��L���U���(I��+���� ����k����v
�<;��T�i�����a���2���(��r�BsR��H�L��HDL̡*_��i`Bd!��͆i�/]1^}i
�U�K��q�u�V�����û��|Խ�6L+MD$���Ｔ}L_՚����R/n�7o+%Y6qVe) e0���([�DDC9BDTPP�([P�P	[`���P���VG��"�%�HI��R��Ǵ���V�!T�T�c֜7�������Z�̌�{5Z�v<UHUI�����V��b��*K� RX�0����b^}�P�*��g��S�Ħ�i�q	e>�oQ��d�Ϥ-�Rl��������
���cJ8���%��ْ�b b4�:M{H� �S�-iM�@cS���YS���3=]<4e�L��&��7��D]Q�2<f-��w�n.�~��G5�,"�mb%S� ����Cx5���k���n��4r�x��O��Z����~��C\~��雟�m�������'PI֛Xg@��=��F"�j��V��w~" O��~M��S4����z�}�,���歯�f͆��ڇ�d��fc5/{TƆ��BϬPeX�2��Q�D��p���� +#h@�!����!?E. �ƂѕD���huRTC��� �"�z��`G�� ��o�����Z�&�Qz�w��y��CUf�<eL���O�xrTd,�X2B����$b�:
�xf�<�3{�D*}K1�ĀAB���0!h��̀a�������D!�����жt����M޻��o�[}����F�,��'����ͻć��ď*A���Rt�-^V��$��%b�p��[HA<a�`� ���tܢ�K��щ�P��-!l*1AF��lbM����l�=Y���
{?�x�=Y��k�
h1o��Ĭυ4�C(�"E���T{OT�ԩf])tj��u{#I���|����) �֬�~��j��|D"R��<�8���8D���M�l"B$��ʼ� ��7S�(�i>�϶լ^�n�ﲹ�l]���{��*���F��* �:�et�볰<+2O�b芚���ĕ(�Q	Py���P��}������ȳ�O��)<x�[�aǇV��~����@���4���n��*�
��5Ͻy�B���4��*���{����z73׍ghq������K������������E1[���
2�P��  ���
��b,�F:� E�Rz�A+0p(��\`��y
(]Yk5����C#��jV��!�׃V�q���#�g*w�ξ(�/pW�j���1�$I @�3n�7�`�@����D�;WDP�@T0�	%[�b)&l+8�b76RT�	��U�h�\�	~'��}����N�25�6��~��	Z�"�	"]��l�
�{��)T��!@��t��i��#Xf��`�
@cy��4@C��-hs�v�n�p�{_�U=4�¼(��8�2�M�[S�XN?�m�(s�5	x.�5>�3��j�I�z�K���O�,=f�{���'��=@5�\�]q�P�#����JNV]R�0��V�V�3BP�t�����^_B&3��R�t ������ߢ��h��t%��2�O����T��^/�k �Tma��0�����?{�J�KM�CϷ��r�若�E�� ������������'���{�	�|�Sx��oy�g���R��޾�gሇ�UM���K:��G�̖"�f�Ve^�~	��!7�l�n[��%�ӂ�-J����ן�)z�+��O7�J�wLZ{Rj���5�X���ʜ �2�H
��N
S�\@�M�Aњ�7Ȥ"(�}ge5�t�@��r�1�A��`�8T��湒V:��}�*�%j�ΐ�E���m�"H���:��`�ύjڽ���D[̀�� �#O�,RD�l1gV�@��5r.�sF))���!R�e�0�-."a`���UjhדX�3���=(*x>V���-LY��u�� ��=�u4� pT&�NвM7
SX��0���vL3(O�<�'j���J�TD  <��:o �%�`�ov ���^rZ�U��Ր�5-mMZ�ЪL�p��Mq��g�n��[Bz��֥��m�h͏��_H}F�Xy�-��׽�O�}��)��a��$	��L77fP��
�����mă�s��2w�v�n��Q&���	6�U�!��o�N�Jj�u5��]�r���5[��ht�ʘj\���AlD���^�Q�2�~�*��~`�L3�j�Q���`���69W`{��$
�����O�G�+����`��e|X�S�
���ޔ|�'$�T�<hIF�kF��PG��r�V�V�̓v.+ֶ�Im���'V���wS�k�ܳ[�u�z�<��/[�]ey�)��ԪI�l���w&�v�@m��d0g(�*��%����6�%P�Q����4`�r�$3����л���ٵ��^&*�W�*ШUi��P�,lM�����Oj��w��(W�kJc�͆ ���Cf�"(U�81B��� �\��{�V0P�Zl��-×a��|Ļ���u��
H��O��T�C��]�rQ�͋�=����v��(��b�.�`���.��9�ƺrD��L��Ϫ	(
� �	�� %�����T "0,��T�2�)��!� V�._�� ���M�	b��GX6�+��:ٻ��5m�*��Z7�6���S�|��β(������h�Z={ċqQ=z�RKK�2��,Dl}�I��,N���9�!0(0r��b��#f�-V"I���`I��7�f���ۍ�<�?`:$�3dN����z��
�:٫��{�����5��x�M�wơ1w"+�[��`�G�����\�3���}4̌��OU�#֌�z�a	J�������9=���G���'�����q��gq�!m@�S�7��T���%����%�XӒ�e��l-=�]����+���f�����j��$��Ic�٬R:�컀&+D�F�¼��,����*�C5Fd@i�DA����2�b�'�f5+�Փ-( R$�FիoP��(2�5��Q��/#c/��2n�G�A���vo����Rf�;2\@� ���l�r�@�Ӣś����O�\ʲ2wj���k=1�B�l@R0b�u��	9<�f(P�le�2Z�p$F(&���d����Lur�Ֆ�R��
�12�����x0(X'�&�-���.���[����J	P�o�Jm�tU�띪�ꋵQz��-g�R�N_Dd���	:�V#���Wg��
��`L�,IrU�TD���*
���n!�-�b��PF 5�����B���O#�-�e	^�@lFT���<'�6N�5׵Z�ֈ��贌����3�L�Z�ZmHͣ�&�+����o�
o��vT((�e!OG�)a�8B�`�7�W�����O�<��֔��|�s�LG��"6q�V�K����YyY�nJ����^��:��*p���T���85�~�4�3�<�ET_������J *5�*˥�v3���k�$9�/!��O����ç�K/�>T
}z�H��'�|�Ki>|���:!�)	��lJڒF�4�Tzh���Bk1�"[�R��tE�uO��V+�����oS�M6,}�[}d}��x��
��!PH=�k%�����(��`�)�X��>6�	!��MHP��D	3� �z�,G� ݮ����,c�f-�|q�5�u*���m�cB��5���+/H� �������Ѽ��x-$R�9�T���9�Br�� 8��ԗ	`A���
)3�
���2z��@�R���RlT-�R0� S��`?r��y�]>�k���ݵߴ=q�e6�Z���<�~��{j��mˡV���Ȧ�+���6*����D���̥� %�L�3�c�j�V��?GS�f`�	 {!*��C@k¤�A��^I2&��0)jߘ�%le�w2�K�C<�<볳ؿ���[;�K<[����V���.��*!��m+��Y0�*aD
D[WHE)���h��!"�3?~�9M�\I�a`!������./���/DH�1����iF�%3�焠-n^�U(��Da��O7_Ջ���׶6'������ڴ��pL��idJ��.o��oK�]�����M��`�Ř��>��9zB� ��o�7_��v����[��/�>����Q誊��/!�Ã��͟+����<�J2�\l�o+�`�D¢Z�E� 5~��$�d�F�-�k�}+v]�D7VX2�W^�J�T����i{�	�槣�!U2�bk��Z'��`�[v��kw�~�%2� n�>�{�8ҌIf$(PM�#�f0pD�4� &�����܎$t��Q^)iՓ�5������Z�t�i�a=�R�P.��	�2$)����<!���JѶ��1FcD@�hID)�T��"P��{�Rޥ*-�K�=�z������(�^�VN��BJ�F�<�u��'5�AD�O���[�q[y{FEP������PB������ws�fԁ��B$���0K56YH� P��8��1�8�ᵕAB�~i��s^���^'���w��DO�ZU��_�.��B^����!��?tf�����0*~=DJ%�>���Ŝ��[�yBN	77Oq�&�֫���k��/�q��BDPR��`���'����'8�(s��4M� ��j�����@M�yW������BS��o���3�(���Bn����\������nșaѪs �_Z��%�ތ\�1�������O��;�����]|v�o5�&|(����������9������<�ђ[R�1b��%�Y\1KY-~�g�7ũ?���@��y��Q�%�ף�(zvh���3!��n�;�@�����7b�線�F���J�Lv�"@z�0{�v@Ĕe��$�P�g5�V"w(3&9b�	%�`W�}��j�����#@JFN�QJ�`��P��r �լ����h�"�(�F�׷�>k��F��Z%�2 �)f��~5\��@�i&���y�R�#�1 F�u����"�!�keA�sQ�T�Ů?FFL� �ϧ�q'˵�H盡��]��8`�ce���4�e��1&K�9��
϶΀e��ʘ��a�:im�|ʼP�T��R7��{U�x ��h� T�ʆ�5T�/D@f�<IP	�o�������c)��%~�i�n�/K��C��nG�V`(j������k�gM�=�S���I�Z:o�v�TK�<"BQ��������equ��d�>}�y*H�#R�8�v�ǓgO��l0������)%��<�\
�	����Gf��%l���7u�,,�%�ô$�َ'9K�@�r����:�җ�3Q��6�h5Z�:;-����)z�LY�u�2]�r=� ��2�������Q��|y���ǃ�+>,����"����]|�o��S����<}ea6��՚��I
�-~���Xr1�doz~d�z���������j-a�3�W��X��L�L��1*#��e���5_]p��aM�5�A{G&�L`����Q2a�#2f�Z
 B�� ;$��5�02�x��F��x����0F�U����W��r�%	���,KZ�v���߮�sk�c	�F�.��j��S�-	�Z7S��pn}�T�JAI�s.AB�H� �(IPf+�4`�ڎA�%F����m��J�5o�HWR��{�'�����e�`�t��S^�g���JʟP��fL'��d��`��ք�Z��e��["�P5LXZ�F��s�X�n{E������9ke+��u�v�1��Q^+�sZ:A��.9�gJ�mW��E�����]��wj���/	5����p���J�Q����R�tx�iNl//��G^�~������ FJO�1��r��a�ʌ�xDJ	Zex�)�sO}���a]���㥯�k�;"��Ȩ��\^c��V��$����z�S�W����I�z�^#3$��6B���?���/������}��O��cߌ>p��������7�v�돤��?U���J:�%�D!ɐ�{2��R��s��r�~��K&o#�j�2 �z-6Ӕ���9x�ڼ�x�h���z�,����|�r-be(b����q,��2n�P��0}��S��j�6���%aFƬ3�L�2c���l�!�pG�C�ц�l ��xF�R���,�z!��OX])t�$����x�,�{_�V��1w�J�
��� �1a@ҌP
B�Z��X )c.Y3rJ��>�gD�F���E)+R*`hQ�ڞ�4�*������S_���5��[h�y��������0+����e"��Q�EiA��iz�7&2Mlg�$��0��T#+t���Ĭ-�ь 5�Ό.!K�5�l�n.�����ڪ�_)�x�ٛAsj ��v��
���F��I�7���W�S_��("]�o���9\Փ�����QE�d�C q@*�<g�R.8'l6#�FpQ�qy}��|�u���x�����}�� �i�8L38D[����	i^�,����3��s���Qp�F��$c���oxnI���J�\�{j5�:+��8n=1L�����\�e ��L	N��
I>�����0=}��}o���x�o��T���%���ax���(��G�|T&�Z��6�	4Z��K?�Lړ��k��S�Qd�� K���Xka���Xv�2?��Kq��/8��V�t��=ʿ%C�6��"F���������ѫޓ�:oAT�X�M��Fւ$3�L]�[�j��z�bε�e�vW���8>@���:C9#�Yp�����S6���εRWt��}�L��n��lb1�w `�)،f�
��֖��c{(KY�KR��X�%�eA��`�C�hQxUkKlԟ�n�?m��
��;Վr���G-�g�hԽ�h�*���! %,^��>FcQ�GҌ[��5-�7�޲��%���q�8�&�ڡ�@�Pڹm
�Ң���[(Gc+Dj��T���E�:/����K�����װ��Y{R�H���3��(��#pzx{�W���2o�C7ԛ���3*�[�@ss@�qq�4g\]]���#���8N3�d#T_{�%�~�d)x��cd���T0�qs{���{�a
��rFN�ĠYd��lRks��t���8Y�;����K���:�������H#���ۺ�I�Z���~���B[�f	�"��A(vn�:m?rI b��t�^��/��>���;�>��ۿ|`
]U������_���{~����h>��2A$�g#����	�j<]!@� �Z��&&�-�D;�5i:��d�V�D�P������e��k���y�H�b:������;�[Љ
;�Ӈ:�KA1��0b[�Q��)����ژT�@�2*�n�aP����lY�(�R$HP䈩�"˄P�B	�C�Ad��$A�%=����!�xe�j�!<d�Bt���&a�1)���u��{+���E��qq���ŦTJ�BEj��"�pE�����焒	4bX:X��Ա�@$BΊTj�
� I	b`��`?�΄cV0�d=�j��P�h�0�e:��I��v% +ͣ�̖��R
��.���?ۗllPh	�U�	`LK)(Z :!ȡ6	1!�4����$"����JMk_]�F&k-j]�
��l����������4�����	����E�֑ �)YIT��ֹ'���ւ����v�m[v�,�Ѣc"]�-L�:�gevF~�>5�n�Y��+;��i�����w�l/����ݣ+l6�4�����f��^������	�b��<���,'�x8����r�m�{5M���#'
�}y���vΔ�q����L���g'���t9 �o�u]����C뫯'��Z~�U�؜�j�$��I~�������������߂����|�o�-�������=���I���t� 5���,Ѥ��-q2B�Y�u�A��ن�W]j��.�`��O(������W5��w�Z���|�$윾�Y��\� ���7}A���[�U-.W։)�M�b���,����f9X'�b���-CY��?:���@��:C���L��E��������� $�Z�o����,ٺ
�nNUa��ߝ%�����D�c�E���m$"d�q��fQ2�T�p HY�&�D"D��`���5z*�\�X7-����o=S<>�K대dzZ�*ζ:XNH�ԖF��=��c��Z9���a��\�Jw�)Ag��^"E! J1_�,fK����rWB����Lw��(�Evk76Hm?��[	(��a����e�`�|v�������a�Ӄ�&�E�5�Q��f��J. �}�j� h�H�S�f8�Q��q����z�-sga�Z�jkKZR��i\ (6�t6`ETPJF�'����#����a�-B���RJ��v��	2�9c�#a�ݠd`;��n�SB��)8��)M�P%�J�!�,,sKe��{�x>I�<Y�;G�����z���c��3���Fw�c/_���>
����:�	l���a.�24-�D"�%A�d��_���y�}+�>�<.}>0�>=~��똏��W��GJ:��Ɇ���#���T�]J��Z��5�^��K�.ٱ���ߟv�[���`
y�1�f�)�=v}rg_��(],����p
�u� m�.�bD`
��jrגd�(�H�ſ�P���EfZj�U�u���Z�EY��U�	a�#�	*���H�,�ea������DKM�Z���0Е!Ж��0�H(�\=j�GV@R��j�s�&��J�zܘ�$"g˼�LP@����Aр���@V�����L���18��ߺ�qCN�����CS>��;���@Kz����q��ǵ�U ���mF�V�3C�2їw_�Gv^�a}�hM;��Ty���"���d"Y�Bɦ���-=y���=�P��� ��"+O�5�i}�W�\=c�)�O�w�V���*I֝�t�m?\��f1�g��i��[_��&@5A���^�j� ˄i>b�#�`�MeZ.���߁����A�f3"��'X�RPJ�dWǨRs�Ob�f��f��}u�V�ק�)�ޟ��q�峽�����Ým��xr�r"_t]]�Ƽ
 *���=.�2�1���O�g���?|�����	�������UzH4g�o�B��$�w�:9M{)Z������dP9��E���U��Xj?������[��7�*rfMU���ݤ����sZ�Z2%���0%�Ɇ���&�B7Nl���i$��5��דs��SR˜O��:#�D��#����<�;ͳ5��d�&�N�������`j�nBAd�z��^/�s�B*�lXw[k�o����[���L�o�m��a� �%�Υ�Bd����T���U��CR׮������x��w��?���Q�]� �����s��vJe�X������֙��������J�+b�!��i��[+�:e��#v-���K^Rm���/�ql�^�:U�
ъ�4/{CZ��v����7BNAulks�AK|v	�-�	�>9�X��*��_���-�R\
3n��|#����)��A�@ ������vLs�������^sr��@���%��n�#�<M�ӌ� ��<�w��u��{KM}ϟ�����-���'��:z�*���V�ja=TÔ5�Xȥ�L�Kӌ m��@Hy�.�����|��o���>�m��'�s5�Z��+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs����|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�f:���E�s�.�L����)������@��w��{n�<��D�^K6�md�c�pcs��yN���I]�$�����i�!�����9�x��=���b��ko@�[��E�S��y�a1�F�bf���W|��	�64졻V�#���޵_���d���є\[���0�h��9N�	���N�!�2�}���2c��?�ߝ��
���{��HI��z$��W}����7S��o=�|ֶ�����]b4�3R. f$ʠ̠\@egJ��%�Ȼ=�T�4�h��]�8T7�1�j�{ȷ#�i���f^���=�d�w=ܲ
	�1Hg�|_��O�Zb#��cE-cm����>AXj��T M�Z�iF��3ي{o�GE�z�E�8c�v�7�n�6��e��I-����#qs��F{J��w`f,�y+ �׽S��=Ӵ���Í�����WV��H7h�!�kO��6վT�#��N�l�N�E��O�2��e9~-�����!�xS�U�׾�19��?W��NH�w�ȥ�"��x{a�p����Zĺn���|r�j������!,}��}cu��o�2�T�6�;�n���1tKY�&�!{��1��]�}zߺ�F��t�*���ER;�H�t����ǯ����z��d�a��x��iW��Hcx��-`�*c�&�b�ns�z$�o�g�{/E$\#>����ЅQ��HIM����+$'�4AZ2O~� ��yM]#�ߌxn���%���L�ځ��ہ�̣��c @�b^�l��1.��cch��}=��&4��ƒD+oB�#��G=t�b��O�Jid�m������>uʫ��C��i�&�T+n%+n圁��){4���g�$��J��kB����ͥ��V�ƃ;�:�J]]w��{�X�?�:�&���=��������O�m�j���*V�����*C�=,�!���*č{��UD��������ݣ��q�=M�\���58.ɚw�iY{���tG����U�-��~���7�O�o~�e���� �il0�C��Ъ��m-r�� {�sB*;P�~�S���� ����x��:П}�{���9 ���r~+��H�X��ԭ4���}�o�@j�#]�^�*$ [KR+�#��W���s�Ƭqtݱ��m�|�6�]�ݲ$�|zYh[=�=��{zQ���f`�{CX��]cX=
�եz�e��i* 5�¾Ag"$����LDA}L����vA��!�Vo��t�2vۤ�o����j���ĭ>�s�����Jk��\,fqO:5+�Y@�����`�083L��&1���e0+r��guU(ߚ=�/��N(d1���WG�1!� �wX��̽���z�ͷ�kߓ�XQ�d�:x����I�H#W޽Y#)���:M̢���t�܈+�$K�d�f�]��D&I^�h9��� M٢>�w-���ugQ��������[�˼`�ŵ��ͫ��}{{���F?n����%��m�4����>��	�s귕��WHպt K���S����TPe��Ċ�#�ہ�Z3!g��tlW}k�Մ,�c��xh^Dp��Hy�Ϙ�)\ER-Z'	@�>Q�ڣ5↳�BU��?��7�������a����^{3D��m#�2ڂ\�������$"�w��;��9�8A�
��r��\ (�N`ڻQ[@y��Ȼ?��?�7�����?�7Ձ �����_�9,K��n�JOr��ip��0���P��NԚ�x!ء�:*K{���G�������c����_���pc����YĲ	k�Yi�L��M�0i�>�O7�77������ɼ,�l{H�7�Q�L�F&��5ܷ�R��0�> �c}����5�%��� 6���m8�/�Nv�j�$~	��A]<a�:s#\WEU=������hJ��-R��y�x>�Ɋ���p�4N���*�f�kǆ��q�'�:G˩E⑏��5�QJ��E��k;������0<�/tv�ֲ�"�PuHޓ��i�l�����'���f�71�:�^��)!!�Y�F�i��^��̮�X.���R�.��*VX^�6�Zl�^X��t�Ϭ�$C}r�n�I-��g�����]��^�W����X�����ӫ\k`�f
p̌R\��>�4�h�v�UR��5ۏjkX*0�Z{V6�͕dG� �_�{���P�u9�I��E���5r3��#�Q���-b7�"]���=j�Q�d��^6��SF*djp�<d�X�4y�������t����w�Agq�����~��K���7~���NzE~�HY���h2�7���rZ=��a�]�o�2�����,k���m�cV9�߬�'76Y�hm.pϫ��Pݶ*�o`�y>���r��e%�y�͐t%� �V�:B�6�I|��9#�y���@N	3^T}x��i; ų�ÓD����5�{�!�l��彘,�^$�)2Ī�uV�M�M� r[<�A�J��`��ŕK������J������@�N	�^��
4��Sww��3�^[/���ӄ=�8��I���Z�:�����������>+�X�����:�^�u[���՝t�+�48�b�/��	>�N���SO�)�&9�5�~h+e0'��m��R�C1��ٌͨ0���z��A��g�y��������@"t��q���z�7�\\��Ū��Vḧ́�ך�_l{�=�$�ު���j\�J���r7������f`8@�V�	)OÐ�V��d3�ن�����u]�P<m)^i,zlp]��v��{Iלޮ�n�l��gA�m+���Kߺt��"������ϻ<��2��	x% R�(�<�ly#�I=�)!BJ�א��s����2�^���A��xS� P���o{���?��~�����|K%��M~W�̓���0��F�Эƞ�j��e{�����@�l��l����]e<�}'H.[�19{xh�gW�z_���
�0�y1��؄�Z�W�ZG����f.���X7��X3#b҂ H�$s�x�i&{���3k��!^?K�ٔi��@���u���:�6a��#^6�x[�sU y�V`n ��y�P������h��=�f���\�b���m��	˲@!�rBNdS����̣*��|�K��]$�W�����f׍y�z�c�S&�������خ_���[���ӱ��f=�����}� aW��e1/�<$��{�잒��!�Ecm�׾�\���@+�2��<	��$���,�v_�쨧��K�6�MX�/����ֵ�][�_;����@�/k�}���~��x�ǟ��vcٌ�_����o�=K e��6�~Y��� MpCI��n͢�Sbp���^Y,(@"F���ڈ��LP�H �)��M�3�،G�{(6?\1�q[�G�H��U�p��9ҿ�h�����8�8��=j�w����!�c��E� W��8O�#�8'(gP��T�<�R�0=��~2��+ǫ{�=���Q�y����~��﨟�9�����Ͽ��?�����"G4,X����C���IA ��۵J�ԇ���R�^/���O�6w��鮘�mB�:�D-�	�.�V>�sQ�Jzh+���R�2]�!�ILloߋglZP?_��IU��b��EO*�����t �4r��mU�g�{}�ȉ�h۞���?��26�5f�!Cү
�MR�Q�Rd�3��n��{���K2V�,��V\^6<)�L��Vۨ�ruh�S �U�d�3 ���խg�!e3D̨i,:��յ���޻�cܧ�g���ՙ��z�F�9��SztC��9z����~���M�A ͞̳�1r�������WkU�|4e@���zw�}-[�;�-���}
��]�2�Ț 9����ģX�0���y�\�|���q�����#i��n?-g��=6�k=��n�z��X��kU���4��"�%'L�	9%;�`�L
挤�T9	@�l�Fk�4r��CY��
z���M�B܈�\�H٣~�������zQ�p��������7�����zU�Yn����n���zU���{�*m�ל���@��(Д�����7�\��mJ{ ����ɟh��}���aqޤ�it"�~����Ư��q�����OO	��1�H��֦�^A����e�B�aH����#T�k�]M���C�7��ƚ�G��.[WF�yzŪ=�ݳ{�_�(Z��Z�V��Y�_���'Q�VJ�D��Z����3�0��t�6v�����"����)ﯕ֜��ٕ�n�9n����X�g�W�ۡ�s�.w+�:Q�M��s���e��+\���-S�n�qy!x��@� R=�n��j/SL)#1#�Aa�2RS�g��L4[;���抔3���L�\@<�6����h��q2���zR�b���M�j�7����Gd���{�CZe�EٚK6.b�֘�(2sF��BW[ߍ�
2�L�T��y���!����sF+tqt�.��y��@/�Z��wz�Q<�]O���zM����Y@���U6��d�{�Q�p��l�x3 s:o�!o����{�Z��li��~�4M`2�k��b�dbO�JV1�'�ͧ�l�*���*cؑ�v9EWEi���O���Q5�e��`|@�����ݯ�*�D7��X�vO��,cF�f�z=Ł�ߏܻ/w.�^�z:]�L}w6c���{p��yO{����0s��e������ `�(~���ެ�it CB�s�(�|]./~��<x����0��ݽ�q�k7�M!��湨����z��u������X���æ�lv�&44���%��t�9��#��4<�ѿO�屛��L�������y�Խi �40��v��`$O(��K��;�m�%v��IM>��=3*(�9�++	�������ٟ{� �:Q�W�JU���QEէn	�������Z�
hJ�1-G\��oy�Ɗ��ZQ[C�L���PB.�zf��y����&X��V@����ē`i���PJ��eƝ�~���W��&�9�f�mk�p�)*�zlN{t	MҪ7��w�Ev������aHٌoej���v;�a�r�l:�P�6��&���N;H���A@*;�i�@��'s�tq	=��.�8����Ji�n��a3�'7�ӣo�`$�\9��#���l���#2�kH�+���p�ѝ��Þ+��I�^���}�Wd��[=���m���b��n����N>��B�x��-��V/n�����G�9m���\�\zAl�
jd����å�>i�H�!��G��,����U~�������H�)Rqs�~�	�ŏk�EG�f��;@��kDJ��C��Ɣ����2퐦�T&�r���i�������S�����7���M�M}�w����s�(>����������K*�	Q����˧���9���e�ՕP��=r`�ʔ,TBCAZ�^�Yվ S?�W�����z�h-�R�ԳC
O���Gچ�\�]�F�����Ⱦ �(�a��B��@�)���j���[�	9�0Q�!gܚv��.pQ�8�=&-��9!��vJ�>'�Z��ۃ��d�ѣ��MW�z���am�{# *r�P�̌&�|D�'���l��{��	g���A����V.�Z��ǓU�i��3�
�Q���a���	mO(��e^���b��dnD*NMq���'2���t+cAc=�t1��}3|��^�E���t�Ve�*���E�x��;��}^wJ}F��NH��9���=\��&{b��кN�y<�i�`KM`�ВВ��!*�߃�'!w��g0JbdΞN�ϚR�y�<��7d��(�ի����U�&��[����Nڣ?�Ag uY0��=?SA��K��郡l*[�N�
�� M7��6�<��#�,H�L�`ڡ���&�,�V�'IR�tEj{��p<][$*O�i�z��CS,�tid�r;��?�z�9���"M�������[Ov�)�S�Z��E�v��6y�.��3aҸX#�}��+Fl_�}��
'���#�����-��:X��D�+�?��2A��\,���`���:�>ޖk��G����S�7�o��C�3�0n������^~��9ܯi��+𣤺K������|�%՞�@nM{ۅ􇗺����V����V�@�W��X���K��m����xo9a��Dmآ�E���ƿ�W;���	9��5�o]�@2#%�BJ�����[�`���T�����3i�e������%v(v%SvO P����=����U��>%�BA���H�_o�̬Tv�DBDJ�oӴS����'䴳��4�ݑ[���Z��¢�V�dJzJl=����`�k(�C��&�s<����&03��Ќ�)�J.���-|�Kh�Q���D6��� �	�+�d��'2�'�����б�������Ƴ�j����ѾǤ;����/xލa߽)����?�+T��n#]6�\lP���*H:���(B"�5���R&P�x�M�4�����m*����S�˧�r@&'�V��o&���5ZU��`���Ƭ AM�A�H9�%e&eb]�E[�*M�*n����������N|�����M�D���'�UIDIUHd�Jċܴ��}��.��0�X�R�)_�̱��� ��?y;��3)Ӕ��_@�p�X�()�	cވ�Z_����dެx�@�!���RaKM�}��M$��IU��u5�!d�(�5�;F��(���F��7������7�S'=`�=#��h��SA�%���r�;�:��ns�3���j�������\��|Ͽ�����?1�2: ����_�ٟ��˸������{�=��$���酪���k��+���q�����f�KI���ja\/"���zC8b�=4z��r{@������G����xiKtE'�zPTm85A�#�d�c����>)I�"��gMH�(^�iyfFJJ9`��\pk���t�|�|@!k� '$0)Zv�>�����������S#JU�-��DG"����> ½�t���!�'�{<pՓ�^K[qF������
9��*�*�T�lҞiwU���v��}-�:�'ngpR�Xt�@p�GiIN��2��e�t\x8N[D��v�D�����E#B*��pk���-­���.����yL��X r��k�ivD�2���MWA���vf����^�E���Y�U@�!��. d*����
��Ҿ��4%�\4��!�"������3v���O@�L��K��'�O�佧��̤��&�ĩ1s#BUEm�.�<SJs���r:��� >NJ�>щ���隠G �rﵓ��"h'-j�,`���W��(���p��C�])�n�����>�|	�U=�&��-mr)��փjۋ�I[+R[��L��$���"�T��HZPX�XG�\���).��)��@�KL��Φ�ժh�J��Ac�>TB����H��nl,��&P����=� �
�V�Aɮ��;�ױH����}���I5��u�g���)#�؝��*S�g���X�H��{��}�E)�K��7��v~��,�Q���w�9���G?���
~���=�f��˷ԁ ������+��q���_hy����m���<1��k�/Q�"%ki�&Hb�0i�N�:���*&X�ܛ��x=��hxI8������V7�U�C&`l �U`Q�PSA&��V�'�W ~�0)R�P�ȔL�L2�0�f1QA��r��i�;�ܙ�`���<!���VA[`�ښ��Y����T���<�Ӄ������5f�� }�2^d�<����h͉+���ݾ*s��n���ҔX.�����2��r��Sʍ�y.Rk���&�eB]
8=U�߯����wcW���������T�E�ITx�j���P�'n)�4/x���Ǚ�JΦ���	9eH3)K&����S�>+n���pkG�mFW"D���+����}��6̨��m�.o�J]ꛣ�^�lm�Ex���~��Z�.���. �Z�����	uf�(�H�V��݄S�q:	��)���gԚ���%��ٕJ�n/|�����S��#_3�Cb<,�����_�į xE��,*ߨN/��[.��[ޕ�)7�,�rc��D¹4"m��kd�e�&Mx7)�De�k�,�jEz�Qr��m�@��r}dL�y*iJ�K�Xu�mn	@Zj˵�,�%�9Km���V淋���R���|�H}mym~B��Vkˡ-ׅuIB�mAʌ�����q��i�����B�N��]ɸ�`\��КE2
d)�vB����hb:]��HPP]Еۈ H��u�Ż+]�����dE�"����Q�;��'�#u�BDS�;oM�{爌Z�q&�a>�@0{�>���>xe�R�#O{�2]q�-�������������R�9�-x�v���Ox���_�{��Oѯ�ҿ���A^�E�� -&�)&<Cb櫶il��R����D��dZ��\���lz�{��f����!���&N��@2AQA3�넂v���z�����+de
��M�1MH�=�N9{�3�JW�c���].pw�w����z*C9!��Ҥ�,Dt��&ί���Μ��S�\N�O	��*��9O'N��ʇ%]ޞ?�3?]�|��r��R3���֟Ih�J���n(������-���Vlr�js�L��'���������9\\�5��Y�q}��YQ�KD�[k���i>��c��[A*Y/��P8=��J��e��yλ]�23@���5��ä�ĉh_wD�/3������?����²]KοNە�9���D�`P���F�1Е�[�pV(�GE�B��:V��� �MՆt:i�_B�	����Δ���K�Zv;�ۇ��R�I��x�s�j��P%���y��SO�r��xI�o�i�Uʻ_W�/���
PK�%���VJie�qj<q�����7e��[,�"��y+��v��	�fc�T2���tЗ#�X��'kgj3P��5�S�L�z���Pv�L��Ί4�EZ�5H���P����"�a������u��Xj�3Z�2�_��m^^���h�۲�g��nk�����T��z(:CeA[ԥ�-���e9��#)���.�*{Bk��:5��m� ���־�D6��SS��' $Ӽ��l�J�#��vng�k)��0A��}��1 h����n<EYi7587"<%��Z,�;��R��xJ;K#��W����^*��J���.>��[�����-w��K���>���4�˸n����?$*���/u~{�si���fH�!��0���n۵b-�=�
�<�����L7��^ �ʱb���߱�l	�W�pya��������+�
����`E6jU��.�֐S�R2�2!sƄl����1+ Ta�
�|�C����%����gO�6����v�2	8w�_Ki����/�gSΟL)����IR�s޵��V=<�T��'>����z[3CiBK�' �g�y�o�z��W�
 �ZѤbYf���=�����^�ƽ|��5?|�Wi̜H[�Z+��L�-;�tGTo�����E�u߄wJ�������rI�3Cs��I�LXTY]S��'��Ki��T�%����z,,`�jR�["�*-��GA��L{�`�-�z/�C�T�R��fPv�RR�uG�}k=�ѓ�Px�&�U�[U�U����Y��ki���R[b�K[�R�)�:/u��~��ݾ�P3�ք_���|Yr������?�z�g����4?q[�p!�ť�|K ��}�SH�ۨ8y����l5����5���?���x~���  �IK���eF���!��m/����y��Nz���г�������;�����<�xWP��@��Y󤏧X�+d�RL�XeW��Rk*��tD=^��%��i����������R���f7�Y�t���A�0N��st���6C��P<r�3�X�\� `��X���/�6ʀ���ƞ���P&Fd��N6��],���H��i�������N����������Oķ� ���G��w��~	iaҧ����.˿�d����&�TZ;B<N*�y7��f�M���G�X��+?Yŧƞ]�.�^A�!�⣴�͏Tتe��ײ�ի������z}�Wu����
h"̲`>��Dؗɫ��r�dNإ	S*&/��g�j�(�w8L�qQ.q�p�������S�Ň��ʴ�r�ʧ	��=�_�����WN��i*{-��|���~���r�0��	���	w��^�w�RI8=8�x\p}\���}������Z�ڽ{�ݿ�w�S��,���=,�	��D��,hMH�uB�ɋM�D�o\1e��.�rb�2A�k�+Q����c�i��~�wW�ֻ���-�N��d�x޷$i�95��Ě�sK��wAV��&a�=0�o�{�M�7\!�*)TD�6�(�q�nr�n�r�ׯ<���8����^�_k�
�gk��.tw�6P��2��O��/t~�{��S�[O���3�[���ew@��HE��}�F��7z������~�+XN�X���f`>bz�I��5˼�\�$e��I�i�z�b�E}7P���4�ҔT�����j|k�C�j}�&�,G���ꅔq<U\_/&*����4pݴ��6�c�F}*�����T� �#&��Z�u��Zunqs[|C
ٍK�Q�H�����5�m��
ǽ��vS!T�^�m�ZJ�۾�T.>���.��?�����C�,���#o�R�'�[�@���/�P2�_��SU����j�ai�;[��&kaZ���R����pk5�9Ϗ�$x.�+m?��O���#޾����6�ի�{�+|���k�W���Ҁ�r�um�>�S�������*6PD�]���p�i��~qUP+ �q��;�{�$��}Wn_�zpk��������y7}\���~��_�}��اtwH�����l��t���^���Ջ#ꬸ���)�N`͠�P�x��5�EЈQ�RFk%��u�_b�9����6L��z���X��^~���p��C���ⷿ�{s�U��g>j��`��p�O?�=}j��km~?D_$�}����\?�;�F�|��x�,f8���"g�����Ԅ�i�i^��+�
���r��;>&�%&y\=�]�pm{��u-�+�P�yʜ���M�Ȥ/{�ڏ�o�~��P8%3+��J�B����bG)#s��8�\v���)���xˋ|���?5���Η>�1(	��5�O?��?�aY�����I����iE�I[��XߢV�0�}h�o�ӽ���X#U" �/���i�-��ke�"�
WU������#��W��'�bC)���QR���(�$L����!>�b`�&ȑӄ[��ؕ���jŔn#c�D	�/���~�ٯ=y��������n�����ҧ_���$4��sϾѷ4��B?�a���{
����an3Z[px�����{���%Ǉ/��J��K��Z�k���bAkC&��^�M	�
�B8͋�N'@��i3/W�Zsx�����F%\�I���+���'�9#%B���d����)���pLލB��Z�l#Y}��	 2��4ٰ�4������k9��J�WA����>���8��-��7�������@�/|�ؽ�i\��h�G�y�����^�N��wf�ߩ�h�����Ui{�Z �Td��^��G��7mܫ��#��f���a�
}������J׆������,*�#� jC|��I��WhRQ�u�K���%d6�f���i���U����\���w��;O�}�c��̻>��/}�ݓ�s����p���7�6A ��_�E �VA�3�y��镯���t�.>Ȍ�6ײ���{ҖI*�r�2� ���s�>m�P���ٔ7��@��xS����]�>�
U�b5�UKIu�����e�i�GǞ�2��qA�x��y+RE`���{ΩW��(/�r?O��r��/Q��H��r��;���/E����=�;��O���`y������SO�vz[m�gAx*ߣ��Է�ջ"� �C2IUXUX��h��d5�㒮��R���Ůq4%+a����{�}�EM`B\���� �����MLPb7MP.>�E-4�4�\�����������������O��,������e���[Z��?��O �^�����>�j~��[o� <xG=]�u��
�>��{���і;m^��T8^�Z5u����54��mmV5�&�'o
�v�k�z#�����3!�U���(q#2��ܵ!o(��p�˔�g��I�.�,̩��2_'N��k����?���?���^�� ��}��F���t~��[��?�ҳ��P��׸x�S}����[h�Ro�N"����P}Z���[*8a�������խ����c_q��
���7�.?IB�,�m��*����>�0��וf�����m���5-˂��Jɨb�1S.Z�W%O��������px�s���/�{�ٷ�-�<�����o�� �g�ԧ���x�|��� rxn�,�����6�<S8�J�U��o"z��o�N�Ts���(��yO
�jz6O���"������
�6C����ܭ-nk�$))aۤ>�i�2"��2%%NB����J�f%>�
����K�ӗ�����qY꧙���F�^|I_��R�L�Uo{���ѷﷄfw�/|�v�j5��@� /����#K]�&�h�Y[M�IRQ6�g"�邈n�-�iOL;UL
ͤH`Ndc���X��J�d�G�*T�`�FB��5���B}�+��De�8-3��#�*�2�~�'�V�J�����<����������O������/�u�4��|��ѷ"�JT�}�8�M����p��~�N��p:ͻZka���:�D�ۙ���������nI�Q�h�k�y^��T91133)"�b��f��@�Y�Z�\r΀���W��X))1	@ں�-�1QQc�
�
�3���9�gN���U��N���,���>+���S�S^��N������¯��'�
�����w?�Y�؏��}�� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��1�Ӓ������   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X    IEND�B`�PK
     !M[d��   �   /   images/a262aa33-74c4-460b-b0ad-c746896f6744.png�PNG

   IHDR   d   d   p�T   gAMA  ���a   	pHYs     ��   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X  �IDATx��{y���u׹���Z�j��ez�����L�b'������2�eH$BaJ�@�dC��`�@��![G6NlϒqO{2��=��RU]{��ۿ�����1�'��n�u�{�[�=�s~�w��ʥ��1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�l�c@�a�z��Ti�R��)�|�H)����]ǧ0�Vg�¸K�F�Z���=:0��y��8L^a�&����4�"ϨH32ʐv4������>Y��6����=�n� ��w�H��)�~�����t�g��!�<T~V�Yz`�����j����ר�����Z�:@N�NF�ޢ���,S�ޠ��NY<�Zk��J��� m
& ̡T�nW���]����{}*f��>s���m�ݽ㯐[����u��)h~�����>�����R����h_�М�NݴC͠���ޘ�g>�?���g�~��P�R8葉ڤ+�T�O�8�,�`�UZ�	!�n�6�a���y6O"ǭVk��D o�D9~G��[�m���^�u�'^"�[^���O�N����+ DF�u
��v�����/M2�P���&���8\��
\��w�z��V�K3�K3���h㇟|������~ݟ����W���f�ȉCD�M"�!Y֕�.���n�Sf�	ch��G�&�q�H5���*o/��%�ݼIj��KI�Z����.J[�(�\ׇGk2�j�4���X:
A�tԿ�M?�Yg����K_����pkC通K�23�*0o�g3�$����0�v�g~�/+�W7��|��ּ�,un_����� I;���\��u��_},�~�n@"��-ob+b�v��X�I��f�L]�Һ^��U�8�E'?vV�x�C�k�;���M�}$�DLi�S����mQ�Ņ�:��(_Ug�����F�����	��ġ`VcrDqf*��q
4SU�NLm&U^�������G��i�8�3�.�۩.tؙ9|fp�[�D����W)�lSg}�����ѡ��0���%�]���pa�[���>PD���~󧢵�� �v���ԡ�����?�j�UZ��ε��@��_
��e���,�=McB�'�pt�&���.���
{^�K�zst���t��I��#���\N������r���4a�8&:��i�M����fS޻�0�*N�� ��%
V^��'B�%���w�1�@��Yuh$L�wQ&�0�3��	B8f��e�wA���Hi��%�?�p-,$|M^�0$ln���ÃN��'���S���;u���}���~g�| ��eP�>Gӧ>�����)3���I�+Q$d���򼴍�*ձ�aѣ�x�M�"D�ܤ,=E��Cdẝ��HKb�=~���kur��0!�-�)���!��D��)�px0D!�`����!��YҞ+sU9��x�T�J�,�OR@do6v�"�J��:������gB�K���E�����Ԡ?±��� ����s�Kh���+��7^mn����&]
wV�:{���i��u�Z�|�I��'��&��=�{��֠}m�r�<�r � ��c%ED��*�	���8k�0�Z��5�׃S�w����i@�g�ׅ�âz��w[�D'��I�Ar<��a�L*�އ\M����G�+�+��߰s[�����
��T�l1�z��=��.� �v+r�v��[�D�KO��c�	�K�N����[_|���S\�m#$ł��y��s��~)�oR�"�qm�ߵU�/�ԃpw��
"��U��2��Nڦ�<���w]B�^�X�U�F�ozZ�3d��(w�m����&�ҳɂ�d^J��)$��D� ]��X0�*\KIy,`Z�S�oا\G�څ��k�ԫ����G(4ED�+�i8���\r;Y_�Fa�bn���V�`���܉'�n��z �}G����#7��{�B���/ga�`:��v!{�%Z�A�q�P�w���~CYT�UM@u�C�D&�����m�O���KY`��Cs5�e@Q�f�\Z�m��-�%*$4�H`ٟ�i2WD�L]VCq�)�~�dQE�:�)IX˵喝
��O=E>U�)��:[[��Bβ�saȜF3�`H)E1��>>CN�?оs������=��;k�.�$�ҩ��x�~���p��_Α7�p�&q�@NTNu����	yф���ά�K���	]�WQ�6���p^S7����N�z��7e�WY��G�95�F��+�ÁBሚ�t�D�,UX�/��p $o�T(M{5�ր�2�gBrNa��r����
�7_׃s̟z���S��\!3X#߳�7��0��p�3��<��D4��Y���b4~�:��˝�7^�H,P��J�ܰ�K핛tv�y��'�w���y�����a2UNQ��8���/#z��!X�4Ee�w�.���9��� �ޙш���.U�5rI?��H�>��!���~�
S%6Y!
F��[ͪJ�亢�"PNтĚ�Ҿ��\�*Ȫ"�윬c�*#��%j��}���y�����﵌r+���Q����5��#w�<� o`Nٰ]M�꿞=��3������i#$�z,�Sm��}ݕ��}�{���ޑ(P���̄ZP^U<P��7�E�)s��p� �Jg�"L��s���8=�8�&Q&	�A@����d��U��Z%p@ e�w�C�� jT���xbn�[惟^��.�ӶxmhI�R�8��X[;��Dn�E~�^��WR# j.�5�RX�_�r�+��]�ʜ-��"���^�t늬դ^��G� x�s�⿸���ԉ?��Q���:�o��� j���g㝫���8��/�(���E�a���r��j�Tܻa/k8S�PY$����I:9s��;��1�M��0RE��<�Rھ��DR�y�2���D�*��$�ETdF�(�8*4�uD)1{6G�����@]-��=F���r��q����0��؜(y�s����@onm/;1�y�&�'����YH��.�KT]xP���SY2�A9qE���	r��������������έ����{>�����@S��/�c��eu��ʘ���	9%�Qڪ��x�"�4a�$ۡN�o��t���"��Z�m�O�ȉ�/SmΞ���%���b[�Ap�����29?gi�IH+�� p"��� xH_�\U�#�8 �=���� �Ʈ��Π�P|9�G�ex����)ݥT�$��5����)L��H��=�c-9Q��3�C���"��BS��4�=w9Z~j;�~����i�ě�}Ű"a��$�ڝ{<��X�1x;"g U.�*Y-���$�0��=��FG*��wi�f���zK�l^���~M��!t`����E�ޗ��5@���R�3�7(T�rl��<��T��;D5�PD��ѹ���d����\�p�!ё�I�#&��Hn=�Afa������[�M�����ox(�}��jߑ5*8�ҷ��D]�kduƵX���E��e��g���s5��w: +�KaS��q��0Y*rc�dZR��+J�*�G�Zc���"4A30��7���ޯ�Q�/�޸D���xs��D�p���.a����6�9%�3ա��XYn�"L[�˭"� �� 1��MR��(a�F��Pcs�6���w�UD#�ƴ�k�:&g�ɻ��P����]^[U��գ�W�s�%���@X���f�S�?��:	���.�B�r8�魐��57�ڛ'�G�͢�k�$�\.�Ӳ3�������|�R�|�|�܁�ڴ���P-���ץ�+Qhlo�)�^��˹!;�S��1C'�aT����Uz+�t�$½�;j�9�d(t��x����m�0H�Հ�"�Yi��BT������5���8R��/6�̽L�FKn�M_r;4��<�\�؊K�E~�%ut���ص;�2��e�@4�����*kY4S���X/���9������
�Y
p=���8�8,Xp��ͽʶ,�{F�>Q�H�Q�Ĩ�SCsnF���g���T���胁őX���}d�$PJR�_Ξ)�
���֠�hGh[���j����'M1��'�>�Hd�D5��8R��,
k"�Y!���C��\Ŕ�AqY�(7��=�b�H�Kr6���e�Nو+_2Kc�����]9ڪ�£���a�Y)@+[3N���?�u@Y�I��2�a^I
��a�|&R��e/Ki�Y����������<}8���$i��{{*2m��"��ZjF�R9\ c�YZ���V�#�j)y�*j�Pj�T))6�����Q�Ƥq��(؟���Z�K�כ�ό��bЃ�l%"w6�s9j�k^\	�m��J� ą�|�(�MҜ[_$9��.e�h5e��ؾ�eJ�F�M0>ߵ�����C���W��4n�&8A�{�^�U,|^x[]��~{�/ۓ��S���r�*��VM:�Ibh*,J2�{`PY��-s�&BU�S��!b%f6zx�"(���u��_NM��ϯ�]	p���[ِ�������C(A��ʚ�&V�%n��Ҳ��m��XZ)�77�lH>�~X���w>�ⴇ�P8Y��e�z��>�!,�S�}%�[��˕�P$+!g�0��Qd�F��-¬��X5�@�iPE�vٟa�T�r7����hޅme���-�a�����Ɣ��;GМ��`��?��{��~�ɿ��'�������C�r.r��Hf@�޾�ѹ���J�ƲЛ�J8����1��� B.N0���=6ۈ3ei��0����E+<÷�V�sI���ϋ{=)�[Q�����#�Ap$�r��q�a(�`�FQО�Y��jî1��X�~�ʍ����C��V!��e���z�3�r�[)W�`�'��?�%��_x���gg�~�Gk�7l>�UH��E�ǡ.J!�dv��:�Ք&�6N���&�1�Ri3צ��=#*�!>�
�mI��P�{�0$j����쵲�ABf�Y֒#����j�����K+GDA�iy_dv�Q��M��T�b���xm.��P�vű|����g�e�X:�JP�W�})B����qQ���H��=���t{��?;�U2�1�	���`���'�~?l.���!Q�w+gD��w��<F��8� ��#$�I�G^�Aa)�un��-O!
c�	����ԋ
�	i(6;��R��	�����|#M�RJd�sRa��
VO^'ANL��Y�k���PY��6��Z��<mMf7�4�t&{,E)�*v�t$F[��1!,�Y�y�s������}2;7YW�����c�q�u�x��T_,.y�}?}�y��,�Ӱc���Z��团�`����)&��|,Q�%�3�Z�T���OD�R����M�όy����|DJ�s�<���O(]��Yx�L�|��X�ǀ�ANY�ؘ 2��H0/n]��z�̍�s�B$+D���"Ys3�T�
Z9?�`NY�h$�(ͲQj�cIQe�_�)��T�~.�t�̳�z�U:�����!�����(��+/�����_s���n�E}��P�{o�����\P���r���J*@S)GG����Ae!ȋ�G\^���P4l�ݞO��+�;�,�}!<��F�R�L���=T`��v������[C�����8/QV�I��@�[�%���-s"� d����uH2��<�P1��:h��gI>�b��I�ѯ�Ch5�������7���st�]��\�v�~7-_x�K��c����YtH��O�-��:�F�"iK�\Ŀ�׏���4�ϐ�x��
�d���Y���Oi+���V���!���h�w�e
 Ң)�;�YِR;@nom��@O���#&���V��UBq���ͯE�.E��4�΂+�5YO�{�F��`d�mp_>��A�Q/���t���h�(��;�_�Ï�|���|����k����W�n�u�1��H꿡������H1��;�^�[��dQ!G��Ȇ2�@qN��A!)�k�ҶVE�V��u2��f�u�k$xn��(0p��]6�F�DSFF!^���+
��l��?W�yn��\Ԡ)v(�6�r�u$��k�
PEO!���$c��'�,]
�Q=�st�t�\���ׇ^�������yo����G����!�v@fg��k/����?���������S�ҡbЅ��e�~i+e%BVG��b�f�n��Cb,�N�w���Ƚ �T�k\�K��'���V��h���]�B�� ^�>]�����lM+�wJ�2u������5)Ly�2�MR�UI5�}��L��k1����k�	oN9Vy�߇�#Y1a;T�&�.����í�~��c������c��i���?0��e|�)�u�T���[itď��FC��'�Oūx��i�\�s����3Μ�-���'���*��jו�6$���-��4��"k����z��J�Z��sը�Pvo]B5��\Q�{߳5�[%g��ٽ)8�eC��0�,~F�_�J��@t�4U�*(�R��#��>�M-�hQ�3�܀�t�m�e�l�a=^s��������~�wx�̇�w�������K��|�vV.��}�?���?b��;����"�e��=�f/.��kT_���En��u:��!j֏H����V��|W;^�K���MD���*��4���AUy���Ss)�f������|��#;���.�u ɎHw���.!��#К��BZG�����8�%��N5O�zGSY�u'�}����O\B� ��Ȯ�H�N���a�'.j�.Ҝ�g)�#p+Ti-Qe��E����a{c��n.�������ճF��w6�S'�������:���H�}R�sn)���>���z�&�3�Uϣ�?M3�����Go�V�3����W_s+��&��N/�G�+���Q���Yz���k۝f�f�����@{��㙄�"����Ju��9�r�i�v������������X��� �:��LT��N{�/)<L����l߭;�f�y�5����ߗ{�<r����.��y/��^"�@�ZI=�F?s �<8^0��U�s���t�s;���H�}oJ��y�V_y�q�����d�����~�v>��n�%G GS+]A1��4��x*�������D�ۊW�=W��k�>��/]�򯷛G���	��P�_'�*�.kqgv{��RoQ7�d�*qR
}EQ��0�і���|�>9Bൕ�e2�-�i��,�bؕ=>'K�w6h8�KG��� `<PRvP<�)���y���?�ɠw��G%�:��=SSt�0Eu�婙�H�Z��S�z��M�yם��?[�N����s�<E5�X�����w3���}ȁG�CwΝ�J����is��*4������V��6}���ȼ���T+�����ڌ)	w�9�_����W~��W.�C��%ZlP-h������}/^�L?N/|�b`|P��֚l�nܜ��U�y�ؗ��ڇ2�[��}�[����<t9`@K���w:�W_���BՇ�{典H�o�4�f��2-��_���[�p�C��
��9.'u!\1���tz�5|�|��>t���W�9��D<����Auߙ'�~�s�"�?�7i��D�����G~��_{)�]D�D��.
ɵΦ��j[Mz��ץg�͆t����q����r�N<�m�W.~���CTi�݋�%�W�ƉluKu�P����FS��5����� ~i�~��wt�?�}�w�����O��O���wf��c�W�c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2f�D�{��w��    IEND�B`�PK
     !M[�c��f  �f  /   images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png�PNG

   IHDR  �  �   ��ߊ  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  a�IDATx���|SU���M�M��ޣ {��Dq�����~�V*�~���(���(�"{�Q6-�-�M�{�'I�M������K��{onn���cU{�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!@��-[a츱�aC�5?�q8�^ݺ"���0�
�"���l�a���>C��p���Oo��vn����"��mE�9F�1\���?ۛ�����(:���c�X���_wlP(�ʔ{���=��|+��#}�Y��mo�w��k��]�o�������?�O�0�?���'�Q���W?s��3��"Sڶo�dՊ�}�I���i�f����gf^�t8Z������^d�g`���>�n�q�0K���k|=Ϗ���5�1��}���I0�p]�y��U��'3r��~'_{���G���ߢ��h������1o��v�#�����޵{�I��z�}Պ�ged��x0'""��!;;�߁�������t8�ADDDՎ��4���N����E�l4"""��L�����QQ���ԿTP�UK���	���sn������BDDDՓ}����{�������H/�=��|!'""�c�4a��sh׮ݔ�#F���u�}�?_+.q��p8PPP��o�O���m+�p���DDDG�}ǎ툯0;+k����C���PA܉��\��+z��I#<r䑓�\y���O5�Q�?�^D��R]�]R<�5k����q֦=11Q�s�*Yǖ�Ull,���0�C�Y6'"�`V|֠g�HKKS�o����T���Ύr���������GXd$���(T�:����=3+Y*��D�~2+3K��H�h#"���sx���_����`:͈�����O��;r��"""
f����6.��p�)�ggg��oDDD�����R�7Mgx�'�����"""
n�Cii����p:M{�'��]��QP3��SSѼE�8���,�3�:gOݟ�F��:�������y�
�DDD���";+;ơzI2�kff&���(��j����H�4�L��at""�`&��:���K@/3�^�a�Љ����nC����E��J膻��0���(���*w�^���(@VV���(���*����:��D^^>���(����p�Yo`� ��;w@/;�����FDDD�Mr�0��mPP�ϵЉ����iB��'ԭiՆ.������Q�V�%""�Qt/w���^J�&�΀NDD����m6È𶁴�{+�Qp�/^�T���t""��g߾m�*���6�Q𲧤�H������]��1�'���i��*w""��g����m*`��r���/��Ä�m�����NDD���3��G@g�;Q�S%�Æ����˝��(��3�����G����ΐNDD�Lس23��i�I��S��)U�ge���'{�3{NN�
����%�;Ճ������zdDD�i��K�DDDA�T=&&Ff��Н*�;Y�NDD�L{xD�t�S�:M�~Q��l6;|T�;�&L�Љ����=L��*w�Su"""
^v�a�ax�&�܉�����0�QN	�U�DDDA�T�\J�׉e���U�DDD��.K�|tV�3�|�i�̽t�U�DDDA��%���F��8tV��rK��U�DDDǀ�����t�K���˝��(���K�z���X���(��E�{	��7���t�,��ʝ��(�ٝO	�:��:űʝ��(hI����4�r��YB'""
fv��a�iz	�n?7�)���(�ٝ�sm��NDD��r���SQ�n��^�n��GDD�쐕�L��T07Љ����)U�J8|�r�Nq�DDDA�n+/�K�g@����<����@=?""�F��0;�*��乸ҵ033ii��k�.$'�@jj*>�����9	�QQ��S�ѨQC4k��6���\���1%>�|��%rpq��+�*3��?V�Y�?���Eb��-طo/<���<W�C=��,|��\`�!6&u��C�V�ЫWO0 }��A�&�f�1�Qȑ��i[�I@���p�{�W�܌���X�z5���;�:��V�ޯJ��(��Q�w�{�>)ͧ�Ė���/s0i�$t8�#�=�\|���ܹ��v��D$<�����pU���Ʉi7`��r��s�C��\�U�^�x1�����n�n٬��E�ۆ�)����`�E���Oq��W���GR���yv"��\�g.~��w|��g���;п_?�i`7нN��¹�}�\�-[�b����Gcǎ�p�W�����=轢������i�O��P\p���������O���u����拓�'�S��o�T!����>���2>�͘����3������_��p���T�Y���tf������ذq#��nԉ�cP'��'������ix뭷�|�2]�Y�^�z���'��2���V�{!�Pz^�0���*RS�µ��Gݷg��g'a��Mw���������{���#R�۟���#G���x䑇Ѡ~}u"
Zy���7o&��f͚���8��yHo���;�1��&��ޔ�y~&M�\�f��`�
���hܸZ�h�:�E˖z8Z�*UGGG#7'�z8ۆ�n�:lݲU�TU�[�Z�QV�a����HOKǨQ#� 1�A������K�,��߁�����Qi�tn��lC�C�����g�><����!??�oF׵kԸ1����3���&M��v�ڈ�{o���b�ʕ�a�:�~�:w���Gf ?/~�$��'�@LT�:�Ca�^��,���eʐ�0���or�gf��_�G*��`���9Q'>�>n��V=��v�Z�ϖ�|/C:�5i�H?�~n��L�<S>�\��S�5��s���[h׮n��z�~Y�(�2+&K�"��n�f9U��W\�Á�U	x���s���Űa�p�9�v\-�_+Ƴ�L�׭Kg�;��|2��֮�ù�J������ѱc�ؿ?K�DD!Nt�s����!�{Μ_���~�2�M�!����#г[7�_+O���/�	u�b��aX�l)�36�6��ѥK�� "�P�c�i7���*w]-̀^�n�ꫯb�d�z��L����p�Wb���hռy�Kƞ��u�@����~�H޶�����{�	�_xK�DD!ɕ�۝�i���q����0��)���_Q����p�����FTI0/N�}�Yg�����ǟ@���(�/3p�@*�y�m�4` ��cP'"
9�����rg��#���,F�9Y�.;ѵ[�G�M�VG%p��,2����/�L񲕁?���?���%]""
I�L�곛�k�Ԛ]B����i_c�jo��L������ރ^=z�R�'�N݃~�os�o�X��3��0s�L�{�DFDT��y�"X�X���x�����X]��:Ne��.��� ״������͞�}���[8�2{�u@|�ٸ��K�ɲ'8�w�{���O��������m=�c���xbP�p�ٟrss�����f��u&"B=�ߞ��y�v����y���Cn^���OV}���a+���N�[�8r��!�1�(ǲ��V�Nq�|����EFxȹʵ)p�>[u�rm��ץ���u}]�����OC��:����9�?���"��\}��ˌ���^��Пc�{�hU��)}>޶�R�5RT�y�s�C~J�@~�V�,�[9C�����57"��_@��U�?ϙ��+V�ۭ%cͯ��zԍ�?�7�/&:�^v	�M��C�0���-lطo�-_���Y"v���X�vV�Y��6`��]f��S�P�,�B�Z�ШQ#�n��:u�q�uD�����JZF233��]ۺ		:�*�>��)�f���X�x֩��s�N�I�##"�{hѲ:v�^�{����k�}^ŏ�r�*,Z�k�5۵k���t@����36o��{�@��]о];Ԋ�����u�8��W�3K��t�	�H��r��!���Q�X������u���lչ5m��}ջW/���u�9��a��5X�p�>Ύ;�q$C�����M�4E��ѭ[7$%��k U��{2��3-=[�l�K!�9n۶�))�����C��(�OL�3A��E�ΝѦMk�V���~�:��.�����MIJ�)���+T���6mB�>y��zK�D��f͛��,�u���㐘X��ZT��gVvv���}<p����_�X�����)�T��21g�(��t���k�8t�(���S_om�&���O<�R�>}�]}�������֊����m����ޭ{w�P��螛�J|���f̘����[�nEzz�����u^��t ���x�s�98��S�P%���w���x���٧��U8r%���5l�/��2ڵiS���C�o������
+T�g��>އ�";4h����õ�^�A�����8;U��n�����/�l�2���w/�k����(u�p�)����N>�$�R�ؑ^�/���<iR��r]d��_��*Hz����ᇙ��/�x�b��>>_�͎z�����5�\�s�g[O��J��`��F�ܰdrd�$���q�#T�T�9���u�	�$xUU��\�M���5�'���X�d����Hp�uT�.�6P�]O�ё"��*�W6�{�U�~1#G�ҁ�0��j�L�#�<Rbd�<������ս>Uw�MNNF���zoR����Z�.�1�sp��#�}{���� ���'��o��H׌2*��ґ��,X6�����?��v��#����.�С�)��^��C�`�l�R������;�ޱ�A.ǭ���*�4h�=z�K1�tP���>��U�ɫ3U[����{����z�g����t��.��c�JXd:ܛo�Y�ʮ'� ��%�ϕ�X��$�9[�
y���N��r��z�8�ޭ2�|��~��^v)U�gR�ve�]�b���ٳ����:���q�*w{�6|���0�Ǚ�Zɇ�J�͎��T%���_��u���<�+�ȿ����_�sGvv�_�+�lʾ��5�����y��ǟxݺv-���I�����B��Z�'_�.w�ځi_}�9?��ŗ\��{I����'g�k�|���z9ϕ+W�i���-�����nՏg�T���p�������KGb�*����?�{���K���Uk���̾R�����'[[��>'�dIAa����G��o֙)��L��M�����Z[j�֬^�u��T&��ge�ԯ���(g�pKU0߽[� �=�%~�q�I�������5�گ�GZ����[=�m؀�^{��9N;{$�6%������/�E]�r�Z����5�m��֩��,ǘz� ^U��7����}(���\�;=���}lٲ�����]J������7'��^��=�ܯ��5sm�?5o���ά���:v���)푆V*4u��p����N����|���f�?c�u�!�_L�[�n����|��"�>� /���]ŏ��VJx�n�\��cǢo�^��r&�9�UeXe�sU�-//��<{s][ɠIFsŊ�駟�裏�_����2��-�S�-��⟩��]x��gT@��&��̊ٵ�̮Z��?���H,���>��I����6��x���r�#����D�Х�2���>���:wB��m�Ӗ���[*J>�9*Q{z���믿�^�)��2�J(2���ч�R�J�H<�!C�v'T�%���'�x����d�k����~����@?���B����3�{5j��4dee��2?E�q80��oUf-�Ox�<�$�*�9
o��ffT�|ſ���Gzo�3�up��8���J�/�_R���>������O���$}�+S%57�F���Ƕ-��f�x��r��0��iذ~=�}�\tᅺ�_�SXO���/�£�<Zl�)��m[6]��������۶n�NjA@�����:lM.��t�t�2[�зO�׉�:�\jf���C����໻����m���WJ�Y��d��bX�w��_�h!��^�����_���*ڋ�	Z�1�w����a�B^���t|߁�'U
�4q�Q��-,���1a�J�=U�9�����NJ��= �r]���1��W0��	�ζʼ�������yx�����K/�Nco��^;i(��?��@���u�ȑ#�h�#!����F����9�[f��zH��������|���ū��s��z�
���zg㪫�
�gYڌ�3K�b�c���+�������Ǚ?⥗�cܸ�������eR:����ǝ�Tk��g��Ѝ�bz͹xť��`Ϟ�^����B�.]t5o(]!OR4��Y:t6o� ��ê ^�~��8ӻw4k�u���UT�h��]z���˖��]	��=gö����Ï�k{�E��T�ק�~��%���#"Ѵi3�B]Su���7';�R��Ҕ�n���VS�JЎ||�ɧ8���|�
_/�]	hLl��h��m�"11QG����uo�;v�;�Yg|�T�H��E_�.�W����=u�4LU%9W{y���D�=M�4Vץ�>o�$��RSS�a�l޴I��[_W�2L�:_r�
��0�L0w]���u�4G����u��n2�Jz��]�V]�dx_�X����(��N8�_�������ȑ��v� ���N��B��I��K�.�3�����Qڵ7oެ۶�'|��C�.Fq6=���=�;�^�I�$��t�2L�<����\ރ|O۴i�{�K�HG�C��r�򹦧�y9w��LӁ��}s���c��A>�G���}��/��\=�7mܨ�[�d��%�ף�t�S�֭[6+��)s���2>�����ak2�H!�ک��H 5��_�|9�?5��`�Db���T%�W^y��#פtu���ԗW��M�:����k�Nx�;�oÓO<�F�h�8Ce�Ru tu�+
�R��ۯ/���J�v�ih�����̈;)q�P�9����oM�R�1�f�Ϟ{n֫���]7�
�u0��3p�:N�޽Ѥq#=��s9���6�k\�����}{���#Ìf��:��^��"�>R�s�v.
�a*A�ޣ7�P���[�j�;W���W�dΤcۤI�����e�	�34t�x̘�طgRS���v":�N9�\}�U�qӦMu	�s]dH�֭��ݷ�����W`���"C�O���}zW����3�ǘ����yp'��o�駝����,���!�1�S��߅�����Y�,2K�s�{]VN����y"����}��ΕΠի� g�u&.��b=�q�ƺ7���zA~>RTfm��%�����H�Qِ�o�}�]�pB=����m곸��{p�-7���]���;u������gj��Q#1��u?�Lɐİ��?��kf@�R�+���D6Х�P������*p_Ub'�|*~�a�q�@Ĩ���'9��x��W�������6g�l��X��mX�z%�W	�۪�Ѩa�J't�P�\��T%���;q뭷��JPQ�L�p))�҅<������>V��t�Q%�����[���x��Gq�E��P��8R"�ݳ�w�'��?��*SeyUR��N�m\�а�8T`�*�G��"�*�ȃ�Եi�Jp�+c�\��-[��u-q�
�R��
�e��B�u��l�kޢ�=4LW97�_��K�jת���ҹ���N�ñ��?��IUb���{�͚4���^֬߀ѣ�ww����'�n��s�mh�2c��:��&������Izʿ8�E/�(ٰr�r�S�O|�Mԫ�P�{]�냅�Q������O�Ї���멈s�m�y2��|�q��aʔ)5r�:�����$C�j�9��nE�Bf��Gq��Յ���2����4��>A�I	��zg�'�q��ϬH�Zž�b���u���1}��qc�}˻C<��&g<�[��c�=�i_M��8B�)�|�ɧx���T�V�6j�Q�G��7�Ꜽ���R%����믿�vxz���T��^��K�DwZ�VaoǑ`0d�`]���۱g�.��lܸIWG׫�$.֊�K|ݺ��8����I����[Ǥ$<���X�n}���H&�ƽ8�{��1ͅ-���?U�1c���nƖ�-�c`��d=#�t���a�ĉX��[�թJ��1b�H]����ɞ�V_]O�II��V�	V��3f`�*9ߦ2��Q��J��u�_��T�3�9?o��!�Ho��]Z��~oSKK��|��:��^��X锸��Zzj|j^�9bz.w��멚�)N:rI��+�['P2�HL%&�6�i�ܵ��.2K5�u7p� =L+�]�#z�����J��t5���H{�|�ǨK/��\gW{�C���]����ݯl'��I�ᤷ�*wk�.=��`^ѡ���:^t�:�D�g=6X�z�J�+��;�w�q��ů"ץW������1F�t}��H�[O<�.8�����{��N��T`�>��C�aݺu8EmW���]���-��V�e��O>����+0��g���L{����t�{�+6��hˬ��z(��g֥〥)�|��a�葅����h*�I��K/�K�,յVs�H��c��	�N���Ց]���g��m�vM_d�p/SfVWs~��ŋ�[0�j��숃���V�ǞxLw[�'�([)�l~��ttx�� u��8��tӍ�ڸ��A�L�������mE��ύ7݄s�����9IIpР���O�x���1t�=iK'��֝�RʖL�ۓ�Fj�>x���J\~�e>k,���*�O�4��C("7JG+����S�#S�Ju�Ν�U���|�M�A�n+̋�Ƌ/�Pw}a����$C}��1�����Nt�p�Zb���W^#�j�G�)S�m�U��y�f�?p $k,��Ͱ�۳�&��KG���l[�V��P�i)��~��7�Y��~i�'�T.��SN�|;�����}�}�a���k�������s7�p�n���qM=%�u�]W���:w�&M���`��G'Z�l��.��2:$�~b}��f���A]�&"#�����)�Oj�V�Z�:�y�xm�>C�u�Ǒ���w�5)P����蒤�NS�*	����2��:wŭ�ݪ�D��.���o���f��.�+K��e:��^�\���0��$��a�k׮���B�{��]��Cꚻ:�ѱbJ��M&a.GMkC�_:Qe����B�+�ۄ�y���$\q���L��OI�.��=��?�:�X�b��5hr�9�<����uĀJ�엨J;�u@_�u�SO;�U��� �p��z���L��U-��V�[a���+���ؼE/S|��s��ǣg��*�JB����m�uQ��^�s��Uj+�2�aa�ͼC��z\�ަuk�{޹z� ��ҿ�.�M���[�5h�Hw@�L�kO@�*yw��	�M�n����̬��б�>k��]/�jb�db��[J�6�`�=D���3�:�[�
h��Kz��w�y�c�UU����0�!�^}UB)=g+P"UF�a��^����r�#��.N����72C��- �>=z�@�J���u��$��ye�лO�J��/���KH��uY�C:�z��(���3o�<����^v��F���,u��x�	i�8p &�5�G��ۇ*�"�Kf�c����(�;YAN'���*s��"1tL�v���u9�����M�>f��ܵL�*�W�L�b���:2ɔ���B�F�4i}�7\�c,XY�K�}9���B:]�t��{��_�׶BSO��1 �Ԇ���qb�>/A+�g��IV�mV�5�ef�U������U+Cw2S׿V-�m��zQ_v�ك��Vx}�k�nh߾j�Hr7M<����J&ϑ9�s�n��^r�ש�������"B���VMcNgH��Ւ����yU��n��sTt�ϭ$G*������٧�`)Î��z�Y���j��ڷw���n٪�l.=����� �+KWT��{�ԓ�4k��e�����H:�1u"ݮ]�J��}]t3���A�?�l��%ǩlgTڶ�ː@���;�`0���I����K[7o�|�y�w53+���m�Fe
7O�d�$3lU�.�Ռot4�_˫r����$ш�Yb1��4W�Ȕ���ɬ�i�u}TsV��]R�����<�b�0��;v�eJ��(qq�t'�ʒ�k�')=���y?�u*�픡��&ޛD\%t9Ve�U��쨌M�7##����=\��[Uj�_��d`�e|v�ڭgᓀ~dLDFE�q��Nz%�*ڼ-��b��/�$t���g���3�I�!���*s�I[]%�Ƃ��͝��Y��4C��I�oU�	��!+�Ig$�6:�t����W+N=j��IЊ�=�Z��k\�V2TU-Zer�t��*S)&	�nݢ�}�H&j��=���_�HaS��L�*�Y��?x�S�W�8��A�@L:TD������YCg&~U���JJ2��M�����۷O�U�w��`���4�eɼ޲�CU/BӴi]��(�8��;��[��.�?G��X�(U:�N�H���Q��H�������܇�}޷G��YO�����Ǐ�믿T�o��ѽ��z�����d�1�F��(8I	�^4o�L��]KJ����MWz]=��i�suj);�7�����/�yJ�99e�2�:Oα2w�T�JG��&�;F5J�$�v42 R"=��M��R�&��x#�k2��q6e�&5��؏�d����j�k�#�\m�5�m�Q�ƈ�]���:�i{�w��`&��[�M�*>
U��1���Idsr+7,�nS�+�����]M��W���e<���X�����z�Uѩ��jH	���n����dLm�zu�o���.;�Ɂ������O���V��G��*@Ib���C���l5s��J.�J�*��<�f"W]HG���e��@u�*��d�;Y����r{��jh@o�X퓒�F�3^�kv$Y6P��7o�3e5o��u�`>?��>�P`��+\��U���Q�*��SNUC�1G9��qk%�Nӽ�0���pk���a��򎥚�gϞ�V�;���˗/׳N�`��ʒ�F^}�5|��7�бz��޽{��%�KOfo3_IU��`)�hf��0HR��g=9�!c��5>�'
��L���C�v�\�3G�f3u���@T1�Yn���5��^*�K`?�a=fu��eض-�:f��#%g�/%EO��c�6����l��ZĐ�3z��K/����)�N�p"	��(�H�`)�W5�s����OT͝Oǎs��
M�?��$&�?f��:U0��8ӟznC�u:N�n[`��(�mHNކ�9�]�]��7�B<�*=Ʒmݬ���ڷo�zi����A�p~PzȘ*�gdT}�_��Z+�و���Ы��`^+�{'O�0J�\h�8��TT�Mu�H�ʽRU}'�zY����?���_�e��]	؇���%����t򓕮�ԫ[O�Ѷ��(��Ν;u�۪v�59���v��1̍f63�٤������Y����mT�:1������]޵Ls������U���v���_�d�R8�rF[�nÌ߫�J�̭>RS�v*���� Q�������*K:ffe!.6�J����]�N�L*Svq9������m�2��Uږ����۷��~�]���R����ft���;�-^��k���Æ�;vbʔ/зO�c6C��gb����|�z���#q֠Az-i�O�^�zhּ6m�^�e�Mz�}\_s-������6��u2;�$x�����BNN�I�d�����K.�Z�%yd^�#��n�Ն^3'��%k�r�U)}���^��u��]vN9i�Q�b��yr2>��s���d6�����mZ���O�܇gq����1��_,�"��u�֣e��
[�n�ƍ��mXY�֭u��(ڨ�^�nv�*��|#d	S�z������H���.���R� 'AIa�������������t�m6\~�e��/�q�:��ٰ=y^z�%t萄���G�)�L@1y��X��?�7��s���0{;�������`�1�Х��Qe
N+LtE�i�쟱{��>���٫�^~��ߊ �y���T@�a񬁕+WaŊ�8픓z\��������s�~��*cQ6@�&MФqc�h���:�����N~3u�	[yU�5��]�}�Νqɥ�`��qz&'+�&M������ȣ�e�i�l���{((��L&�hּ��'A��9���[q۱}�f�*���]wމvm����ٻ3�NG>���ckšO�����}'R �=$�����s����>uON�2����.\�_���Ԕ�أ�d/:��]�>�p�'�se6s����巽BL��:/l�
�W]}��6�[��e����+HHH��s"�ë얔m�*�?�̳ػ�[�z"��.��{�*w�R��ۯ�;��f����0u�T64`S�����|K/���ŤI��úw>ё����3�w��S8�����^ݗ�^���k ��r�ÙY���U0���;��2�UI=�S]�h�����z�I�YN�l2����~�m�a�S��p���؟��}N_��o����W�|�^�/��,^���dNt��7�|�.e�:ݎ^��?�|UZ����&m�'N���N9�J�/9�e+V���^Cf�� ({+JO�s�=͛5�B
$��ڧo�4�GX�1�=9/�8mޜ����W|e�Q���o�nW;g�uV��i��ЭÏ4�y�d����Ə:sJ"\݀7� ��*O��+/��6]���O�^<p?ڵi��	D ����3Ĩ��x��`����E�.]�>�Yg���y�υU_��[6���c�L%rmZ�:���j߇^��*�[�V�hѪ.��|]�
���O��UW_�y��!+Ӻs܌�CR�x��'sd�Lxz��^�cǎՙ~o��N���5ADd�^��j1���<�Kܒ%�ωe@p�v�����ª���n�{�X6d��a�oa��ŸM��SZ������6�I]6mقw�yWW��L���NJ�W_}���
�۞eY
��oT���*�;�����J4�0t�0�ya:�kW�DN��c�.<��p|�ŗ��l�$,,�^{-�w��`NU��s��_���V�z~~�|��G������n|���ҫ�ɧ��?{�j�v��|��hP�~���ccbi�?��}���3rM����t�SB7ٖQ��XRU7��0l�CؽSz�Z}A}����O=���'�����y��'�u�V��c^r9��,lܸ�~����5V�Ҭ����X�W<s }����}���~��3>��S��e%��_���}��GqҀ�^�&��Zi..Z�J*���7��/�p��	'���E�������{J��}��WGw��.:s�����q�
�����"G%_��Q����g��Y::{�ٺ�����w����<k�̾t�����z�T��n_���N�e�U�Zn	ݕ蒇L6q�嗫l�	��jއ��Ds~�	���;Z�j�~���G�����84i�1��:�K)\������{�`ٲ�X�d�.�oS9��Y�|��LO��1ϣm����}݄x�Y�իWc��%�J䤏��ٳ�f�\}�5�����!)Ig ��N:mڼ	ӿ��>�[6m.�WYN�l��?��^�`NUi����{���#��]z���eMM����q���~-[�@���}f��`��ǧ�->��l\���8ѵ{<��Cz\zM����j�ɢ֭�z���];q�}`��i�ԩ���9����ߥ�q�1��+�ak�r���6`�ZD����_�uz���F`�~�+odC��v�����٧vĨĠN|��)�H@�ǲT@Vw�����}�߳|�I'�ŗơO�^���ӫWO�5��s�^��[-Į�;0�����T/5+��e<�L#����g��)Y�p!�'o��᫆����`��0���@T��b-*(�y�ر};�y�/C@��z���xRe�'O���w��4j�	ut'���=m�r����زe�*I�.��{�F���SO���WMIg�}Ʃz+U��s�^�ru2���4���as��2q�i������G��T@/�#�蚢*\����$��z��c\r�˗-��Jg�[��d!�Çӽl��J���0���{�y1�Yt��9 7�9C�F���裏b��M�ԥ��k�v��~�=�UxD�c����<��Ư��M�5�SÇ��T����hеR*0H&2?� ���C�v�m�#遽i�z���˯��uהφ������3#��y�&x��q�X���d������u2
���X|�\������{�a���HP����z�Q^���ß�Rsx��e�^�6mZc��Q�q��ɖ��\+o�:W�L�ÿ��[q��w�I�FKdH��a�����ß��E���^)z����I���ʕ[�ҵ�J܆�63���&%ntlɽ�X}wF??J��ߞ�6�I/k�Mi�W��*�+�[^F���mݦ-�����
�\�����G��X����f
�))ػo��Ŧj�
��k����={b�ĉ��������H�|=�ze��W��SO;��s7�W���$��;g�^Fv�8���-2����U�9�s��:�	���K����ݺu�Čp�3���^��:�=��Ӻ���W^����aZ� X�E�ʻ���=22��q�}�����DU�]N_�#�=���{?v�H��A����HNN>f+\)���ˣ�����?��ުґCf�[�j5������G���!O�[OO[y�5W��s��OH�۽kL��:��x������,l.�H�M���O���O9�]w�^�F&�����^!N����5Z��W�������@�S�Z4���q��^��z�Ksp�	�>����*�e���G~y]lt4n��z=c�dοV���7��~?3��C���
�Q1�ر��Tw���6jРR���Ɏ�{��^�Z���bu<��qD��Is�|��F��}\(oi���9nӦ��=Opv�A�Н�����Ti����õ�K�L���m.���lݲUw�������HH�G�vmq�	'b��A�ӻ7��M�[�*Ty_҃]ޓ�������3�`�?ر}������К�fG�
�mU�\f�2dN:i �={+}��^�[�e�v:�zᜰ��Wmʾ���t�ֽ�LWr��I�V�!5r���֭[�kWu���Ǒ��S�Jur��=�d�%�v��!`��ʔ��{�,�w9���� ̋.׿Es�믎Ӷm�A�Hy�:��2r�sz����9?��ʕ+�����ɽe\
Oa���Eb�D����w.NS%r����Vi�٣�
n9% ��e��/=���tb릮yZڡ��/Sjk���W�\i^�fK��|���i�Oزy3���c��B��Zj3dTP||�����K����]],�J���մNG�s��gC�t�8�3t�;v"y{�^&TƖ������Y���HH�ڵ�PO���5k�\y�W]�fw���[�9��&w���ur�v�Y�F�N�e��Y%#=]�Ws�$*�j��^f��ر:w�W��#d����׫�	Z2���$�뮻���V"""W��+�I���>����QQQ~�ŕ��qϊ]�#>@���S�/�r�p��}e�#������-7�d��|b��+}lԵ�N����6m�ڵk�z��}�����lnn���bս.�=˒��ڵC'��v�{�Z�Z�
��s;��S��w�-kO�\�����S�|��/-�%� _��C�:�����Sqݮ

�����~%'�:u�ѨQC4i�T��1�2�S�
Ԭr�"�W݌�*ˣg����ِ\���5���@$��A)J%J2�Qj�����_��%�o��>�]� C��2w�zߒ ��� ��Ë����}�u�Dӓp�:�ʪ���qU{�o�VD�=��������"�LU}��qq�Q��)�/�I���&=ⳳ���ס�}��$�(:yHf˰�O�H/����r�;P�7��aUu<O�Tc��Q�9��k������΀^)f�K)C�\����b?�w,��#��L�im/��;�hݥ��8��|��8ގ)�ňp�z�����<��58��0K���0�~L��6�@;�\{u�yy�PM����Ni��f7����YB'""
f�S\�[y:�Q�ѝ8�)������^����3�-ӯ6�|v�#""
b���������(�ٝN��ֈ���7=S\�[�,HN�Љ������W~	]�9:����T:v���3M�r'"":�����,�Tn�7+�O"""
�K�ݯ8-%tFt""��d��m�::QPR1����DDDAKW��UBg�8""��e��˝Et""��U�:#:QP���U��8t""�`&U�~lU�?"""
F��ΈNDD�̊��3�)݆ι܉���;��~e/w""�����,�NDD�L��YB'""
jXm�m�DDD��"���������r�z�DDD՞S�r�5""����U*�}�k�r'""
ZR���VN�f,'""
fz�5?7eX'""
V�ߋ�0�'��,�U{�˧2�5?�r�܉�����m�r'""
b��U��DDDA��Nq�����(��~W�Q�b�;Q�Ǚ∈�B g�#""
~�C�˧2�+��^��DDDA���2DDD�ʏ�\�L��NDD���ΨNDD�����*w""���*w""�`�ʝ��(p�8""����kb=S+'�܉��B ;�U\m������K�p.w""�����\�DDD���X�U�DDDA��Q��LqDDD!����,DDD�*�˝m�DDDA�ɉe�������CgX'""
R�
T�Q�͉e���B��m�&�܉������6t"""
F�U��Gk��DDD����܉����
t�#""�`���WЉ����Dh�m��(񃈈���aT$��UBw8�HKK�!�p���� �`PS
Q���c�=�l����j���둓��ז�n��0l�C��Wæ�5�������]8
�������p����*�&6���e��-�8\yS~U��^�t1����h2�g�.��6��sDDDt�I��f4��&��� ""��JJ�:�烈���+UB7��͖n:�� ""��Hfsأ��ege�U;6�-3:::�^�n��������{�g��0=""�I&������K���;w$�Өqӻ<�t^^^/�4cTD��u�ƪ�3*8���c:1ϑ��g�#|���g��OF��x���$�����jժ�y�����W�<l��k�ŧ�O����;v����LP�F��]mn�G���E��l6�&m�v��0�æ�`ap�4�����rd��ϫXf��Ta���
�+����ſ�F�_JoWl����l�	�Q�k1׉x����󇢿B�8*�g�J����b{/���}����(:f��Qxn(���.u��{�`[�~���0T�.b�ҥ�{v�
/���G���NC�&M�T�^n7TWr�֬Y����[f�������=��ILl�o�Nɟ�f��MX�<[Q��}y�~����1�\4%�Y�wϮ�����,�{������vW��3K���yxv�c?%�l�Kb�R��\��W���)|q9��,q%��[����ĮK��}���n�a���{��_�]�r)�'�z_/)���N�l�b+��(�-6-�Y�b����J�-��ڨ�9��G�}{ΧԖ����t��pJ�e���%���-:�b�G�J�JM����.rџ�ݠ��:IϹ��\�������0̘�hg|BvIIs�����Saw���ʇ���G4�΅�Ϡ ?W?j"�gY"P������Ӑ@�p��ÐB�l�S�t8W pr�����T$u:�Õ��p?����w���&���\]$�b��$�o�^ܙ���kѾ����m6�����u�]o�ٽ�ً\t�Ÿ��[Bnn�;z��͸�λt"Q���N���on���'�<�������OOL�<O�EyUw�g��&�%�f�L������õ�Y�I�?\���u����hY<u���	S�,�;u):/��s�]6
ӛb�r�����
_��G���R�����̰�^����kc��4�ͦs�6Wy��-5�0�\�����6�]^cs[�e�._�CA��o��0RB�zHٿo��>�S?�� O�l٪UH��7�

���Vtx�is8t��4��J4�m�j��m�w��/�(5�_�O!_ega2�J%J��#��X�]<�g�إ{�i�'6�^�٧�Lexb�Y��Z�;�'���|��������Jl��2y�.�-�܌Ȉ��Zu#WD ��x���\���j�ژ��~̯s~Y߿}���E���[_a��p�2�mW|�ҥ�R��(�P�F�s+��(��/��(]�*��2�M��x�k�9��?ós�t�<�t�B�{��#�?=�Og^�{Tx6�k��F��'�����ܙ��r����w��=��M\�C���x�y0e[��|�}������vU��2��pU"R��Ɂ�
��c8�Զ��r���گ�S������r�Jt�ܹ�ug����e�,���o��� ����W;����"�#

�eF���e���سgZ6o�/S�T婌���o�c��-]:�mҬ�ks�u���'`��u���+AD,Щ���T<�$$$����J��ʬWr[�l���kt@�`.�;���*CS���f�^��?�>��t��6��{�Q0a@�2ڷh�ǞxR�����v��V&����a�?�`��A�>������_<��sػG��R���Jn߱ø���vh�] "
F�d�q�&�ݧw�_|�^�ڵ����������:��m;����x�駱j�
������f͚���/s�~y��6�w�� "
6�d)-��p|n���V���]*�J[�j5�nۊݺ�:ҝ���1f��y�l�i80ԫW��O>��/��Lꐄ�cǂ�(1���N�#:&f�
�y*�G��¦;�-Y��������λ����(�	N����h׾ݘO?�$%'�0���:Y�6�6m�ʔ���#���5*�M^n6����\s"��Q����{���K���@��0�=�Q��o��}�'�?�fM��;�"�`ŀN�.��b\{��6�#""|Wf��Ȫ/���K����^�jӎ.�bي�1b$��މ��\�����g��w�;��>�Y'>�G<"�`ƀN^����۴9�����U��Uv[�n����t@�$������ѣ�d�b�	�JtTTr��-�L�655/;DD�:y����`r�ڴi�Ff�*;ͫ��b�e8���Q���㭉1��o`5���W��k�.���� �n��O?"�`ǀN^}�~.����j���s�yyQ��q8�p�"���"*22��g��oLx��ٰ*�׊��ѭG��Np�����޻o���:`@'��M�ݺ�@TT�&e~^nS�v�U+Wb_J
Z4k�`�i75r����`��y���ϛ�����C��޻Љ��`@'��z�\vŕ��Ď�QQ۳27-���m۶bÆ�A�u��~w��b�vs�ݞݰA��+W,[8��G�Գ;n��jU��S߾}p�ק�<{�Z〭�%�:tK�.����`$����˒�����|�)�ߓ���mxi� "�N�ɧ����
���e�Ͷ��뻗�t`ѢE��ɑ�AՎ.'+��'�h7���]ٮ}����-c��� "���ɧ_�͚�D�:�W���g��^�j;iG߻oZ�h�`�״����p���n7���hܴ�����)_}��K�aԨ "�n�ɧ��.B�=l˚ի����Xt��۱~���	��SRS1z��^Ǜ6�,����\�պ�k0�|���K "��Щ\	uиq�ݪ�%=-�M�-����y��y�5�fϓv�I����v��:uz��/�ʱ���)�����b@�ru��I��9�U�a�Q�c�t`������Flt�1oG�v�7&L���[��#���7o�r�/?��y���ؽsN?�tUW�T.w�8�{�^�򚣠� �j�U+Wa�޽hӪ��x�#Gc��vsy6���s�͜�����O��3O���:c@�r͚5]��@|B����������e���ؾ�֭?f��<�`�E���_{�����/���w'OQuǀN�:��q�7�t:��/]�+++�n٭����v��:��(���y�EtL̎�mڌ�����0 ��Qv;"����_�z����/��?x�`�mLӡ�S���BlL�QoG�����7����`n���7i������3#����`ND!���Ҹi�rӍ��:���l��]y�e���ػwڴnu��MB�Ju\�j߻w,�����P��'�<��AC�1۶m��oL Q�`@'�<��Ø��iG_�J�9y+�Ihݹs'�o�p��������`���n��]�v�g�������q��_3�QHa@'�HǸ�I���Y����J,�v�e˖��AgU�9I0�/(��＋iS�I�?����#�7i����[2���ѳ[Q#��ÀN~��q=��t"۵�߅�2�3,�V3��ѳ��sƣ�4�g���k��΄U����s/�`J��]�v�Z<x߽ "
5���m����n94��S��`5��X�z��KA�U3�g��u6�y�w��˪vUX��]��Ν;��釙Y���� "
E����Cҹ�ٳW��av�� ?�2��x�M7VY@��JO�ر�������n�ڢeˑsf��)�a��_����Q(b@'�=8t(>��+ԩS{UDDxFA~^�	f��Ұt�2�y��*9��~�?|���0M'���e6���Mz��W�r�x���0⹧AD���o���Z�i���M��ѻ�23�Xm�׽*�G����ܹxy����̀uU���s���Mxz�3�5�[��ND!���ֿ�?^Ƥ����/������m�5�Wc_J
Z6o��K0߲u+F��m[7���m�ڷ����{�r���_���?Q(c@�
9����1))�s�n+m6���Hޖ�M�6,�K0����K/��彩�-�����4m�t��?��9���дi\q� "
u�T!��ɨ];			K#""rsrr"�n�jG_�l�vj@��0M|��g���>���U��a��~�ĩ���K/3���1�Y��Q���N2��3q�"22r}dT�����&V������%K�������J������k>^�"2��[���ۻ��*�<��?�����n4$kBGMk׭�bv�r�s'k7��f�v�Y�j^Rlk�Uh3#l[��dE!0�&"��*'8��e7��s�[�<|?3g8����w��9���L����ܶ�3� ���~�>*J���k������%��8m�F�Y�Dz򃴘מ���5k��\���G�|}[Ǎ�� ���T�|~�3y��' ���~�6�f��ҥm�3�t��_`�Kjj���ٳ
����Z:;e}F��������zWxDĎ�~����
� ?_�n� �pB��oK�zJ[`ƞp�m%��e����A�%-�-RRR"���;�jQ��y_v��]v�����	:���cGW@@���1��v:��Ç%.>ABCCK||}�m6k�����V)*:!]6�x�}:��W���Xa��MY+��f�����	�����Z�N��M*{��:�m������gŠ7T;v��J{{���_�|%M�&�w����74HRR��*+�^Q���ᆌ=|��W^����አc@�B�d��Sr?ʭ���0�Ӹ��*����	z_h1���ƍ�$���<��
�?w�?����/�k� W29�$��ϲ.%��*�~���p3J�su^ZZ*�Ϝ��s�ݷW�l�"6�U<͛�Un���o�ަ��RXX(��� �pE�1 ?��DG��M�'����X-���q6[�?^$֧�b4��禥�Dq�$'�H���t�����=>�Ճ���; �.\���x�ጠc@���f�~��������k�X:�=]Mk����-�q];��,)�k�d�	����N'QQQ{�WO�?c��v����+ �;��������L1u�
�k/{�$?w��������&[�n�?�#�}��Z!�!E3�e���hjn�m��  A� ����c�>bޙ�uZ���{ڨ���(��e2c�t���ҝ��'37HW�7ڢ�r�K�Z~:yrʮ���t�3R[^..  A� DDE�,0��_�Sl��~�����(/���EEb�Q����{W���%yM����Iϭv7��Fo׍��;�צ~x�;��Ȋ�� �_6w�,���Hxxx�ȑ#-�W�~�o�����XZ��亠����F6��Jj�:���/�Ӽ���ZdT�;�ߙ�>����%9�� �w:L�"uz\����-��dn�����R[S��o����)ٻ����i��%A����3��^{�g5���*� �C�1`�G����>Ѿ^��Ω����t��_� {��S�Iz}O���]��.�X����s����s�bc7�d��ߕ�P�1���y� ��:eF|��
h	)3��6���8m]��۷K��Y2g�,�8wN��$u_�WK/��i���_�Т7W�|�.�,~H  �"���ks��y��t����ߔNj��%=-]���$c}�=rD<=��]�GFF��=gv�ƍ�N����
 �cP^߲E��#gΜ)�;엺�����򤪲J*����Ԗ�u?o8j��֙�fnX���g�!�>yR  �t��%�n�Nʻ�|\z��t~�)�'��MR�e���i�L�]���훶lq���ɯ�<)  �:�d2ɒ����������ں��tz�~���w'L�X}Ͻ��ݺu���ݻD�d;A��tZ��J�:m��/>q����ā��%�GZܽ s�����j��u�̝@t�'��˧G���;�x�iʦ���X�V����`0J\|\ުU�v,8䊈���� �aC��?��{\Ǝ���?���b}�.�K��`4��W�Ǜ��j����pF�1$��^��:f츎�G������q���>��K:�n[xT��i�ؤ���[� �Cf�Ν��ޮm�r�������T����C�i�+��<�����-�  ����2˖,��/���s�J�ط���w���-���*<!!��]wߕ|������� }G�1���ِ������l�X��m�I=��������3>m�^9��ŕ���*/���  ���cH͙3Gv��-oeeɁ��"_�$�ݑ�]�Qn���z�;f�y��g�9��ӈ9 Aǐ[�x��d2���D����t:&8�UN���|�����`4�1��Eǋ���ʤ��V  C��8UZ*:�QBCB�'LL375�X::��lA:�����'wtp��u��wZ,�z�j1M�$ ��!���86ih��^��������dn�:V: `�:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
�O��Ր���    IEND�B`�PK
     !M[��EM  M  /   images/d3694a2e-5bba-40c3-8069-8db85c4c9209.png�PNG

   IHDR   d   d   p�T  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  cIDATx��]	xLW~��d�(%�J"��}�%(�Z���B��_[y~R�R[u�E[[����J����ҿZ��j��B)��'s��;��Ĉ����>���=��s�s��-�37:�PTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��AW÷&��z\I���7�)I*�Ev�Z�:d;iJ�3mtRɲ�������V�$IY6��"a[�d��$}/����~�l���99��t.��$u0Z��d�M��(��5D��a�}0�*�
��?���h��dY~�`ȫq+��L��yY���@���[���������ƍ����0��`�Aк�C��"�|<B&�������r����t�PQ:�;w'N�{˧����a)y���3�t>���ʂ
E@fB\yyP� �f�3b�1�(p�3!�<ÃY=��䫄(�d���?0��&1A3vH�JIi�	�YCd��c,�p?��0���g�Ж���lqtws���%b�G��ɒ�2d'jaxR�v�Zl߈s��S�����_C���2Js;�i���8�f�ɒM>�Q.]�����С�x�g/�5J<����зO̚=�g����f6.:6lX�t]������B��5�D��;ѽ[7���s�p�0g�,�n�=_x��(���E��~/���u{���F�m�6�2�h��!����v����;����dX�i5�7�}�����ٿ�2~޳?��#n������1p�@xV�$��u˖�Ѳe��H�zi��|��u��,�Ν'�����ԩ3�/�5PP��7o���,�_���C�޽ѵK���ǚ5k�t�:>�,^|q 4�XȺ����7!&&�+{�_�~��d��ǎ	SԥkW�o؀������A��n��B�p2�7n����Na��>$3��ARLN�G��&����~�� �����QQ��wq�������Тe+xU�ºu_ lQ������͐�լ�K�.����ԙK�.��9����(�QN4|���X�p&M|�����5�OLLDu��x�"�.Y�9o��&�l7ww7�b�rD�c�)��?��޽E��jO����[���a�0�?B��ۿr6n����o�Y�}��E�E�:uh@lAZZ*�i`5]�ر�u�9Ǻ��<s�4�V���ի۽��1�Q�n�:AƢ����D�?O�F�g:b����a� i4puuÑ�#������W��u� ̜�iL8^<H�Ȏ��ʕ+Bui������®�v�u�zS����u>l�ФΝ�P�U�@.��+��������^M�5c�L�L��S��nW",�Y��e��'""#�|���'B�B�FMТœ8���	�R��ӓC��w��t�b�_G�R׿ƛG߭~=L�6U��?���קў��ݻ[��Z���\�rLd0�q�	��o@Ey.D<kI��
2^U��~�zB�!C^65V�E�6m�W���$!-^�j� ��溃��������͂�٤������m׮j׮����{��l"��e����G�fg�AQ�%{ΫbM�6��F�흚6m"�.\@�ƍD���]P��	��g�ΕG���e?h�V��\��ӊ�����ٳq"m���`1i.�[8c:fd��Y����<P��6���׻�2�sq�{dDG2kd'j	h�͛��)2;U�jW��%�=z|j���)�b~b����!JcӁ�L��+$3�i��ߪ[�Fc�8����2�F����~~���dG��?��%\�9���ɡ���3lw[wGDD���Ç�6�V�Z8AQ?��6U_"���YԢq�0��$��_M�i������W[P��@�nns+�F*Z��@'����!����ǤI��`�<a�CI�>��p������<*T�[�Cɩ�1K�,>�>}�/�h�M�vhD�*��89�-�aq�֭�M0m�t�jQt������5k?C��M�ۻ�Mk5���Z�e����ZSVY'�����L���������'����F����g(4�Ŷ��P�^G�>|<(��p������_�R�VUDK</`9rr��WhI�6��E^��9��~��΁�ʧ(��K�c��K�^���}Ѭis<���b�s���J�efp �e
���,���5��<�5o۶oD��h���%.�sab��F��%a�ȑ4I܍��u�Ȗ-�!00�==̤?�9@���������A��"���K�T����J��2
�������r�̋h���C�Шn+���\�t	�i~`�'t�dA�����Ӄ|�'���GEDCQ��z�5{zP�gA`�@��?�h����\�h*��5���]�r^^^pbb(��1��[ޒbo�ػ^8�s4�叽|�4�@����4}�#0(h�my
?A�#����Mg�<��7��?�il���_ �2Eto�����"����j�37-N^��4g��)�8����&��'�*JBCLQ�JH�C���=d��,���}X5D�2`�����0��g窆(&Q#,���!�.o���e�TF��[���9ʲIQ�[�<l�M�V��|/="D�xOR���vG�_G�3˚��7��aj�gE��s�6��ˋk�Q'I����܊�GBEiB���j���QCG�h4Z�D�$ݢY�-R��By%�V+i�T���I|3����4����ĉؙ}���2r����)���Om�fk\]�zH�|�R�iO�l�Mۗ�I6_dْϜf4G��Fk-匷�ݥe�k�\𛍶���V���_�3���X:�-�b(ڴ#ݾ���KĤ����h$�v!VI~}��+s�^����xg��p�h4"�E@�Ӈ$^N������1���	�����ǁ=j��������o��qbZW�?��i�1��wI�t�G��v��e��^3�x޹���k+�t�w��`-;q<3��rJ�r�##���Κr$55G��޶;�a�±c_�ٿΜ�V�{J9�Ԕd��=�(B���}�\�.1�7����׭w�^v�.\�[��"{x<����̣������{�"o���]�|ҵ�"#��[v��n�ٻoޚ>�Mۢ�̛;[�A���(Ks�#�����@�V�s��I������׸��������gn�fV��8\��@�*e	%F��#�n�����8v� �2�Ǎƙ3�2+yV{<6���ܜ����#d9�¡��ȏ ""�z�ז-_�M���^nzjJ�QNk��i�܇��#��~_�Z(_��?���&��2�G9��ɡ�=�gge|�yx�fY$�Q�/R~�'������ll���<����� ~�N�z�����t
s�PVQ��<^�q�s��mOrrJ@�=�t-���K		粲24x6�;�;�%JHJJ
*�|D��-KKMN!p5�olI�x��ݺ�Ge�F��kǏ�H�"A�ռ!i\�xzz�/_�<�R�u�7�u�����U�F��K0��N�rx����̬L�(B���^b���x:y9��}���E������k��%u����QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB����Blg���    IEND�B`�PK 
     !M[������  ��                   cirkitFile.jsonPK 
     !M[                        �  jsons/PK 
     !M[�qE�>  �>               6�  jsons/user_defined.jsonPK 
     !M[                         images/PK 
     !M[ZR�y�Z �Z /             ; images/f51f6ed9-d8f0-454d-af8a-e11415a94f15.pngPK 
     !M[�����"  �"  /             �w images/53dea2ad-2eb7-451c-84a6-1b4fef66a2aa.pngPK 
     !M[��F�} �} /             �� images/b63deb06-c33f-4ae3-8f73-25229955b1c1.pngPK 
     !M[���  �  /             � images/a5640015-ff5c-4848-bb8b-6d4b42e5489b.pngPK 
     !M[�wp�&
  &
  /             #+ images/1cdb40d8-22d5-4761-8204-85ee5f97d036.pngPK 
     !M[!��Ů  �  /             �5 images/9ee875d8-7c7b-435c-a3d9-92ac29f03ab9.pngPK 
     !M[����� �� /             �8 images/99708c53-ae63-4787-a3c4-6dca09af2b7b.pngPK 
     !M[��P�#  �#  /             � images/62b25533-4940-4036-93a8-d94b028d26e9.pngPK 
     !M[	��} } /             ' images/bbfae99c-8036-4c5e-89fd-a87441410720.pngPK 
     !M[d��   �   /             c� images/a262aa33-74c4-460b-b0ad-c746896f6744.pngPK 
     !M[�c��f  �f  /             ;� images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.pngPK 
     !M[��EM  M  /             i,  images/d3694a2e-5bba-40c3-8069-8db85c4c9209.pngPK      G  @    