PK
     �)K[3��C� C�    cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_0":[],"pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_1":["pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_1"],"pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_0":[],"pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_1":["pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_1"],"pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_0":[],"pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_1":["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_1"],"pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_0":[],"pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_1":["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1"],"pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0":["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0"],"pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0":["pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0"],"pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1":["pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_1"],"pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0":["pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0"],"pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_1":["pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_1"],"pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0":["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0","pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0"],"pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_1":["pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_1"],"pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0":["pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0","pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_0"],"pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_1":["pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_1"],"pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_0":["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_2"],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_1":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_2":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_3":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_4":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_5":["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_16"],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_6":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_7":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_8":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_9":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_10":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_11":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_12":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_13":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_14":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_15":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_16":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_17":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_18":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_19":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_20":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_21":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_22":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_23":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_24":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_25":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_26":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_27":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_28":["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_15"],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_29":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_30":["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_12"],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_31":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_32":["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_9"],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_33":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_34":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_35":["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_0"],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_36":["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_6"],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_37":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_38":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_39":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_40":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_41":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_42":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_43":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_44":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_45":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_46":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_47":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_48":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_49":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_50":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_51":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_52":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_53":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_54":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_55":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_56":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_57":[],"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_58":[],"pin-type-component_101dbdbd-a855-4798-9242-a7c17a09d383_0":[],"pin-type-component_101dbdbd-a855-4798-9242-a7c17a09d383_1":[],"pin-type-component_101dbdbd-a855-4798-9242-a7c17a09d383_2":[],"pin-type-component_101dbdbd-a855-4798-9242-a7c17a09d383_3":[],"pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_0":["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0"],"pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_1":["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_0"],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_0":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_0":["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_35","pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_1"],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_1":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_1":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_2":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_2":["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_0"],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_3":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_3":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_4":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_4":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_5":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_5":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_6":["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_36"],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_6":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_7":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_7":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_8":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_8":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_9":["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_32"],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_9":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_10":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_10":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_11":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_11":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_12":["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_30"],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_12":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_13":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_13":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_14":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_14":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_15":["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_28"],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_15":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_16":[],"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_16":["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_5"]},"pin_to_color":{"pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_0":"#000000","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_1":"#000000","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_0":"#000000","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_1":"#000000","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_0":"#000000","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_1":"#020202","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_0":"#000000","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_1":"#000000","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0":"#000000","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0":"#000000","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1":"#000000","pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0":"#000000","pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_1":"#000000","pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0":"#000000","pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_1":"#000000","pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0":"#000000","pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_1":"#020202","pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_0":"#ad0000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_1":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_2":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_3":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_4":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_5":"#1a1a1a","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_6":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_7":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_8":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_9":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_10":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_11":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_12":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_13":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_14":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_15":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_16":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_17":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_18":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_19":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_20":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_21":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_22":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_23":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_24":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_25":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_26":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_27":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_28":"#1a1a1a","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_29":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_30":"#1a1a1a","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_31":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_32":"#1a1a1a","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_33":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_34":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_35":"#1a1a1a","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_36":"#1a1a1a","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_37":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_38":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_39":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_40":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_41":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_42":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_43":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_44":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_45":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_46":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_47":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_48":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_49":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_50":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_51":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_52":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_53":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_54":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_55":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_56":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_57":"#000000","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_58":"#000000","pin-type-component_101dbdbd-a855-4798-9242-a7c17a09d383_0":"#000000","pin-type-component_101dbdbd-a855-4798-9242-a7c17a09d383_1":"#000000","pin-type-component_101dbdbd-a855-4798-9242-a7c17a09d383_2":"#000000","pin-type-component_101dbdbd-a855-4798-9242-a7c17a09d383_3":"#000000","pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_0":"#000000","pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_1":"#1a1a1a","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_0":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_0":"#1a1a1a","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_1":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_1":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_2":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_2":"#ad0000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_3":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_3":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_4":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_4":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_5":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_5":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_6":"#1a1a1a","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_6":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_7":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_7":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_8":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_8":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_9":"#1a1a1a","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_9":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_10":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_10":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_11":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_11":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_12":"#1a1a1a","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_12":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_13":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_13":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_14":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_14":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_15":"#1a1a1a","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_15":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_16":"#000000","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_16":"#1a1a1a"},"pin_to_state":{"pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_0":"neutral","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_1":"neutral","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_0":"neutral","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_1":"neutral","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_0":"neutral","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_1":"neutral","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_0":"neutral","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_1":"neutral","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0":"neutral","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0":"neutral","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1":"neutral","pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0":"neutral","pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_1":"neutral","pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0":"neutral","pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_1":"neutral","pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0":"neutral","pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_1":"neutral","pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_0":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_1":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_2":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_3":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_4":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_5":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_6":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_7":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_8":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_9":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_10":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_11":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_12":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_13":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_14":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_15":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_16":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_17":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_18":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_19":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_20":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_21":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_22":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_23":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_24":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_25":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_26":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_27":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_28":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_29":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_30":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_31":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_32":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_33":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_34":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_35":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_36":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_37":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_38":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_39":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_40":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_41":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_42":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_43":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_44":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_45":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_46":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_47":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_48":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_49":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_50":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_51":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_52":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_53":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_54":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_55":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_56":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_57":"neutral","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_58":"neutral","pin-type-component_101dbdbd-a855-4798-9242-a7c17a09d383_0":"neutral","pin-type-component_101dbdbd-a855-4798-9242-a7c17a09d383_1":"neutral","pin-type-component_101dbdbd-a855-4798-9242-a7c17a09d383_2":"neutral","pin-type-component_101dbdbd-a855-4798-9242-a7c17a09d383_3":"neutral","pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_0":"neutral","pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_1":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_0":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_0":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_1":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_1":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_2":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_2":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_3":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_3":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_4":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_4":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_5":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_5":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_6":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_6":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_7":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_7":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_8":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_8":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_9":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_9":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_10":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_10":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_11":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_11":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_12":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_12":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_13":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_13":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_14":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_14":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_15":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_15":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_16":"neutral","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_16":"neutral"},"next_color_idx":2,"wires_placed_in_order":[["pin-type-component_a3ae65d4-c858-4cbe-bb67-1538767c17f8_5","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_7"],["pin-type-component_a3ae65d4-c858-4cbe-bb67-1538767c17f8_7","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_8"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_29_polarity-pos"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_13","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_28_polarity-neg"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_29","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_29_polarity-pos"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_28_polarity-neg"],["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_1","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"],["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_0","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16"],["pin-type-fake_0","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16"],["pin-type-fake_1","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"],["pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_17","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16"],["pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_12","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"],["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_0","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_1"],["pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_0","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_1"],["pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_0","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_1"],["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_1"],["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_1","pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_1"],["pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_1","pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_1"],["pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_1","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1"],["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0"],["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_1"],["pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_1","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_1"],["pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_1","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_1"],["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_1","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_1"],["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0"],["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0","pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0"],["pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0","pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0"],["pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0"],["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_7","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_0"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_8","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_0"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_9","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_0"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_10","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_0"],["pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0"],["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3"],["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0","pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0"],["pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28"],["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0"],["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_5"],["pin-type-component_b00b0f46-5dcc-4451-a676-221697210905_0","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_4"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_19","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_6"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_16","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_7"],["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_5","pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0"],["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_28","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_0"],["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_30","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_0"],["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_32","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_0"],["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_36","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_0"],["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_0","pin-type-component_101dbdbd-a855-4798-9242-a7c17a09d383_0"],["pin-type-component_101dbdbd-a855-4798-9242-a7c17a09d383_2","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_35"],["pin-type-component_101dbdbd-a855-4798-9242-a7c17a09d383_2","pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_1"],["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0","pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_0"],["pin-type-fake_1","pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_1"],["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_0","pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_1"],["pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_16"],["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_5","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_15"],["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_16","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_5"],["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_0","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_35"],["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_0","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_35"],["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_0","pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_1"],["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_28","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_15"],["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_30","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_14"],["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_32","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_9"],["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_12","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_30"],["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_36","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_6"],["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_6","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_36"],["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_0","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_2"]],"wires_removed_and_placed_in_order":[[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_a3ae65d4-c858-4cbe-bb67-1538767c17f8_5","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_7"]]],[[],[["pin-type-component_a3ae65d4-c858-4cbe-bb67-1538767c17f8_7","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_8"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[["pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_7","pin-type-component_a3ae65d4-c858-4cbe-bb67-1538767c17f8_5"]],[]],[[["pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_8","pin-type-component_a3ae65d4-c858-4cbe-bb67-1538767c17f8_7"]],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_29_polarity-pos"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_13","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_28_polarity-neg"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_29","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_29_polarity-pos"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_28_polarity-neg"]]],[[],[["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_1","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"]]],[[],[["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_0","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16"]]],[[["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_0","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16"]],[]],[[],[["pin-type-fake_0","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16"]]],[[],[]],[[["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_1","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"]],[]],[[],[["pin-type-fake_1","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"]]],[[],[]],[[["pin-type-fake_0","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16"]],[]],[[],[["pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_17","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16"]]],[[],[]],[[["pin-type-fake_1","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"]],[]],[[],[["pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_12","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"]]],[[],[]],[[["pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_12","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"]],[]],[[["pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_17"]],[]],[[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_13","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_28_polarity-neg"]],[]],[[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_28_polarity-neg"]],[]],[[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_29_polarity-pos"]],[]],[[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_29","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_29_polarity-pos"]],[]],[[],[["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_0","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_1"]]],[[],[["pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_0","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_1"]]],[[],[["pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_0","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_1"]]],[[],[["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_1"]]],[[],[["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_1","pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_1"]]],[[],[["pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_1","pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_1"]]],[[],[["pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_1","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1"]]],[[],[["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0"]]],[[["pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_1","pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_0"]],[]],[[["pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_1","pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_1"]],[]],[[["pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_0","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_1"]],[]],[[["pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_1","pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_1"]],[]],[[["pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_0","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_1"]],[]],[[["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1","pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_1"]],[]],[[["pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_1","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0"]],[]],[[["pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1"]],[]],[[],[["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_1"]]],[[],[["pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_1","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_1"]]],[[],[["pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_1","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_1"]]],[[],[["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_1","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_1"]]],[[],[["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0"]]],[[["pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0","pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0"]],[]],[[],[["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0","pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0"]]],[[],[["pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0","pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0"]]],[[],[["pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0"]]],[[],[["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_7","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_0"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_8","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_0"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_9","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_0"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_10","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_0"]]],[[],[["pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0"]]],[[],[["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3"]]],[[],[["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0","pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0"]]],[[],[["pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28"]]],[[],[["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0"]]],[[["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3"]],[]],[[["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1"]],[]],[[],[["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_5"]]],[[],[["pin-type-component_b00b0f46-5dcc-4451-a676-221697210905_0","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_4"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_19","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_6"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_16","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_7"]]],[[["pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_4","pin-type-component_b00b0f46-5dcc-4451-a676-221697210905_0"]],[]],[[["pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_5","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14"]],[]],[[["pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_6","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_19"]],[]],[[["pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_7","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_16"]],[]],[[["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3"]],[]],[[["pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_7"]],[]],[[["pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_8"]],[]],[[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_9","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_0"]],[]],[[["pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_10"]],[]],[[["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14"]],[]],[[["pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28"]],[]],[[],[["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_5","pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0"]]],[[["pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0"]],[]],[[["pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0","pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0"]],[]],[[],[["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_28","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_0"]]],[[],[["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_30","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_0"]]],[[],[["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_32","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_0"]]],[[],[["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_36","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_0"]]],[[],[["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_0","pin-type-component_101dbdbd-a855-4798-9242-a7c17a09d383_0"]]],[[],[["pin-type-component_101dbdbd-a855-4798-9242-a7c17a09d383_2","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_35"]]],[[],[["pin-type-component_101dbdbd-a855-4798-9242-a7c17a09d383_2","pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_1"]]],[[],[["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0","pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_0"]]],[[["pin-type-component_101dbdbd-a855-4798-9242-a7c17a09d383_2","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_35"]],[]],[[["pin-type-component_101dbdbd-a855-4798-9242-a7c17a09d383_0","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_0"]],[]],[[["pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_0","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_36"]],[]],[[["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_32","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_0"]],[]],[[["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_30","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_0"]],[]],[[["pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_0","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_28"]],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[["pin-type-component_101dbdbd-a855-4798-9242-a7c17a09d383_2","pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_1"]],[]],[[],[["pin-type-fake_1","pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_1"]]],[[],[]],[[],[]],[[["pin-type-fake_1","pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_1"]],[]],[[],[["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_0","pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_1"]]],[[],[]],[[],[["pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_16"]]],[[],[]],[[["pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_5"]],[]],[[["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_16","pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0"]],[]],[[],[]],[[],[]],[[],[["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_5","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_15"]]],[[["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_15","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_5"]],[]],[[],[["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_16","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_5"]]],[[],[["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_0","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_35"]]],[[["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_0","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_35"]],[]],[[],[["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_0","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_35"]]],[[["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_0","pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_1"]],[]],[[],[["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_0","pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_1"]]],[[],[["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_28","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_15"]]],[[],[["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_30","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_14"]]],[[],[["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_32","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_9"]]],[[["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_14","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_30"]],[]],[[],[["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_12","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_30"]]],[[],[["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_36","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_6"]]],[[["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_6","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_36"]],[]],[[],[["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_6","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_36"]]],[[],[["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_0","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_2"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_0":"_","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_1":"0000000000000001","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_0":"_","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_1":"0000000000000002","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_0":"_","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_1":"0000000000000003","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_0":"_","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_1":"0000000000000000","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0":"0000000000000004","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0":"0000000000000004","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1":"0000000000000000","pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0":"0000000000000004","pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_1":"0000000000000001","pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0":"0000000000000004","pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_1":"0000000000000002","pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0":"0000000000000004","pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_1":"0000000000000003","pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_0":"0000000000000011","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_1":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_2":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_3":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_4":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_5":"0000000000000005","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_6":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_7":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_8":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_9":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_10":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_11":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_12":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_13":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_14":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_15":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_16":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_17":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_18":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_19":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_20":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_21":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_22":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_23":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_24":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_25":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_26":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_27":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_28":"0000000000000007","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_29":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_30":"0000000000000008","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_31":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_32":"0000000000000009","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_33":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_34":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_35":"0000000000000006","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_36":"0000000000000010","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_37":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_38":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_39":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_40":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_41":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_42":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_43":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_44":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_45":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_46":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_47":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_48":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_49":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_50":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_51":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_52":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_53":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_54":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_55":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_56":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_57":"_","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_58":"_","pin-type-component_101dbdbd-a855-4798-9242-a7c17a09d383_0":"_","pin-type-component_101dbdbd-a855-4798-9242-a7c17a09d383_1":"_","pin-type-component_101dbdbd-a855-4798-9242-a7c17a09d383_2":"_","pin-type-component_101dbdbd-a855-4798-9242-a7c17a09d383_3":"_","pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_0":"0000000000000004","pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_1":"0000000000000006","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_0":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_0":"0000000000000006","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_1":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_1":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_2":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_2":"0000000000000011","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_3":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_3":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_4":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_4":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_5":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_5":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_6":"0000000000000010","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_6":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_7":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_7":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_8":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_8":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_9":"0000000000000009","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_9":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_10":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_10":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_11":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_11":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_12":"0000000000000008","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_12":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_13":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_13":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_14":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_14":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_15":"0000000000000007","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_15":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_16":"_","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_16":"0000000000000005"},"component_id_to_pins":{"f7b311cb-2dd2-4362-af91-c7568e208d66":["0","1"],"c059b081-dcbb-437e-bb8b-813da336182d":["0","1"],"4d0af7ef-6915-4a65-b658-362c305c51f1":["0","1"],"07201ce6-242e-4070-beb1-6b1ecc8e9a32":["0","1"],"2829c8e4-4312-47ed-a029-8eab57667ef2":["0"],"8bc6f0d9-3ee0-4f84-84b0-8d65a769c427":["0","1"],"d430a89f-cf84-421d-97a9-6ef91b5385bc":[],"5078f55d-6889-4bc8-828b-a676a5fdd005":[],"1cf54da9-56c3-4f81-b121-cf75a7c03fd4":[],"3d6d4311-3b96-41a7-9347-33206381a263":[],"9d6a5121-9e9a-495e-ba64-f8cf5049df87":["0","1"],"68792fb0-2eb6-44eb-88c3-d5bd97335509":["0","1"],"5bff362d-8f79-4a23-b1e8-04253d472f65":["0","1"],"a21c1a89-038d-4d33-9463-f2151579a9e0":["0"],"c03fea7f-e196-404b-826d-0177413f616b":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31","32","33","34","35","36","37","38","39","40","41","42","43","44","45","46","47","48","49","50","51","52","53","54","55","56","57","58"],"71023eac-aa29-47f4-a674-909b27edbf73":[],"de9b39d1-1e28-492b-9be8-7de288cd2559":[],"e3e0359e-9bb9-44ac-80e4-66e3c1f30411":[],"49914fee-a25e-42ff-ae99-52a23942b71f":[],"101dbdbd-a855-4798-9242-a7c17a09d383":["0","1","2","3"],"07dde854-559b-49ac-80f5-aa8b57c2b5cb":[],"11263eb5-b485-4dae-b6c9-21c18e7b3a28":[],"72fd138d-67df-44a8-bd00-9e004d450883":["0","1"]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_1"],"0000000000000001":["pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_1","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_1"],"0000000000000002":["pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_1","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_1"],"0000000000000003":["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_1","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_1"],"0000000000000004":["pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0","pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0","pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0","pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0","pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_0"],"0000000000000005":["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_16","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_5"],"0000000000000006":["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_0","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_35","pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_1"],"0000000000000007":["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_28","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_15"],"0000000000000009":["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_32","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_9"],"0000000000000008":["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_12","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_30"],"0000000000000010":["pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_6","pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_36"],"0000000000000011":["pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_0","pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_2"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000001":"Net 1","0000000000000002":"Net 2","0000000000000003":"Net 3","0000000000000004":"Net 4","0000000000000005":"Net 5","0000000000000006":"Net 6","0000000000000007":"Net 7","0000000000000009":"Net 9","0000000000000008":"Net 8","0000000000000010":"Net 10","0000000000000011":"Net 11"},"all_breadboard_info_list":["bf214f1e-c792-43f5-846b-d34128e4e83a_30_2_True_955_100_up","bc941250-d2ab-4f36-99ca-60371a583e71_63_2_True_835_10_up","295e808d-80c9-46a1-9a2f-f0256ea548ee_30_2_True_940.5_145.49999999999955_right","633b310a-2a82-4082-91f6-b1a17256c96b_17_2_False_355_204.99999999999997_up"],"breadboard_info_list":["633b310a-2a82-4082-91f6-b1a17256c96b_17_2_False_355_204.99999999999997_up"],"componentsData":[{"compProperties":{},"position":[268.35808900000023,399.8462299999994],"typeId":"7c3ccbf3-d039-4eec-8ff4-6af5efd4a31a","componentVersion":1,"instanceId":"f7b311cb-2dd2-4362-af91-c7568e208d66","orientation":"down","circleData":[[317.5,394.9999999999991],[219.90399999999954,394.9999999999991]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[268.35808900000046,354.84622999999965],"typeId":"7c3ccbf3-d039-4eec-8ff4-6af5efd4a31a","componentVersion":1,"instanceId":"c059b081-dcbb-437e-bb8b-813da336182d","orientation":"down","circleData":[[317.5,349.9999999999995],[219.90400000000045,349.9999999999995]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[268.3580890000003,309.84622999999993],"typeId":"7c3ccbf3-d039-4eec-8ff4-6af5efd4a31a","componentVersion":1,"instanceId":"4d0af7ef-6915-4a65-b658-362c305c51f1","orientation":"down","circleData":[[317.5,305],[219.9040000000009,305]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[268.35808900000023,444.84622999999965],"typeId":"7c3ccbf3-d039-4eec-8ff4-6af5efd4a31a","componentVersion":1,"instanceId":"07201ce6-242e-4070-beb1-6b1ecc8e9a32","orientation":"down","circleData":[[317.4999999999998,439.99999999999955],[219.90399999999954,439.99999999999955]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[93.13070049999988,488.4428929999996],"typeId":"98d6e125-552a-4063-90e5-58c04872effd","componentVersion":1,"instanceId":"2829c8e4-4312-47ed-a029-8eab57667ef2","orientation":"up","circleData":[[92.49999999999977,469.99999999999955]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"GREEN LED","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"8","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[212.2250186155993,372.84760038547086],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"1cf54da9-56c3-4f81-b121-cf75a7c03fd4","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"330","displayFormat":"input","showOnComp":true,"isVisibleToUser":true,"name":"Resistance","unit":"Ω","required":true,"validRange":[0,70000]},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.25%","value":"0.25%"},{"label":"0.1%","value":"0.1%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false,"isVisibleToUser":true,"name":"Tolerance","required":true},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"string","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false,"isVisibleToUser":true,"name":"Number Of Bands","required":true}},"position":[157.22504875383424,440.6937378115408],"typeId":"72c75556-baa3-04e7-55a5-e13f447c8c5a","componentVersion":1,"instanceId":"8bc6f0d9-3ee0-4f84-84b0-8d65a769c427","orientation":"up","circleData":[[122.49999999999977,439.99999999999955],[197.5,439.99999999999955]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"WHITE LED","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"8","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[212.49349844410642,416.72261565132703],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"3d6d4311-3b96-41a7-9347-33206381a263","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"330","displayFormat":"input","showOnComp":true,"isVisibleToUser":true,"name":"Resistance","unit":"Ω","required":true,"validRange":[0,70000]},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.25%","value":"0.25%"},{"label":"0.1%","value":"0.1%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false,"isVisibleToUser":true,"name":"Tolerance","required":true},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"string","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false,"isVisibleToUser":true,"name":"Number Of Bands","required":true}},"position":[157.22504875383424,395.6937378115408],"typeId":"72c75556-baa3-04e7-55a5-e13f447c8c5a","componentVersion":1,"instanceId":"9d6a5121-9e9a-495e-ba64-f8cf5049df87","orientation":"up","circleData":[[122.49999999999977,394.99999999999955],[197.5,394.99999999999955]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"330","displayFormat":"input","showOnComp":true,"isVisibleToUser":true,"name":"Resistance","unit":"Ω","required":true,"validRange":[0,70000]},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.25%","value":"0.25%"},{"label":"0.1%","value":"0.1%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false,"isVisibleToUser":true,"name":"Tolerance","required":true},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"string","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false,"isVisibleToUser":true,"name":"Number Of Bands","required":true}},"position":[157.22504875383424,350.6937378115408],"typeId":"72c75556-baa3-04e7-55a5-e13f447c8c5a","componentVersion":1,"instanceId":"68792fb0-2eb6-44eb-88c3-d5bd97335509","orientation":"up","circleData":[[122.49999999999977,349.99999999999955],[197.49999999999977,349.99999999999955]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"330","displayFormat":"input","showOnComp":true,"isVisibleToUser":true,"name":"Resistance","unit":"Ω","required":true,"validRange":[0,70000]},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.25%","value":"0.25%"},{"label":"0.1%","value":"0.1%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false,"isVisibleToUser":true,"name":"Tolerance","required":true},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"string","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false,"isVisibleToUser":true,"name":"Number Of Bands","required":true}},"position":[157.22504875383447,305.69373781154076],"typeId":"72c75556-baa3-04e7-55a5-e13f447c8c5a","componentVersion":1,"instanceId":"5bff362d-8f79-4a23-b1e8-04253d472f65","orientation":"up","circleData":[[122.5,304.9999999999995],[197.5,304.9999999999995]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[483.1307005000001,473.4428929999999],"typeId":"98d6e125-552a-4063-90e5-58c04872effd","componentVersion":1,"instanceId":"a21c1a89-038d-4d33-9463-f2151579a9e0","orientation":"up","circleData":[[482.5000000000002,455]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[743.5261630000003,275.2762280000001],"typeId":"a7ff864f-ccec-4557-bfc3-03323186baf4","componentVersion":1,"instanceId":"c03fea7f-e196-404b-826d-0177413f616b","orientation":"left","circleData":[[602.5,485.0000000000001],[587.5021750000001,485.0000000000001],[602.5,470.000018],[587.5021750000001,470.000018],[602.5,455.00003150000003],[587.5021750000001,455.00003150000003],[602.5,440.0000540000001],[587.5021750000001,440.0000540000001],[602.5,425.00006900000005],[587.5021750000001,425.00006900000005],[602.5,410.000093],[587.5021750000001,410.000093],[602.5,395.0001065],[587.5021750000001,395.0001065],[602.5,380.0001275000001],[587.5021750000001,380.0001275000001],[602.5,364.998062],[587.5021750000001,364.998062],[602.5,350.0001815000001],[587.5021750000001,350.0001815000001],[602.5,335.0002009999999],[587.5021750000001,335.0002009999999],[602.5,320.0002070000001],[587.5021750000001,320.0002070000001],[602.5,305.0002265000001],[587.5021750000001,305.0002265000001],[602.5,290.0002310000001],[587.5021750000001,290.0002310000001],[602.5,274.99818050000005],[587.5021750000001,274.99818050000005],[602.5,260.00234000000006],[587.5021750000001,260.00234000000006],[602.5,244.99820449999999],[587.5021750000001,244.99820449999999],[602.5,230.00032400000015],[587.5021750000001,230.00032400000015],[602.5,215.00241500000004],[587.5021750000001,215.00241500000004],[602.5,200.00036450000005],[587.5021750000001,200.00036450000005],[896.4015625000011,430.03928599999995],[896.4015625000011,415.0061854999999],[879.044360500001,427.7600299999999],[879.014945500001,420.51514399999996],[883.4956435000008,350.24113999999986],[883.4956435000008,343.92620149999993],[883.4956435000008,337.6099744999999],[896.4015625000011,270.5561869999999],[881.3795020000007,270.5561869999999],[857.5295110000006,179.9562139999997],[842.5951855000003,179.9981389999997],[857.5295110000006,164.95625000000007],[842.5951855000003,164.99821999999983],[607.8706390000002,140.99075899999968],[601.9109275000001,140.99075899999968],[595.9524160000001,140.99075899999968],[589.9939045000001,141.01495399999965],[859.9435000000003,248.5204999999999],[859.9435000000003,209.38099999999997]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"GPIO26","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"8","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[456.7022493395014,288.4004146975199],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"71023eac-aa29-47f4-a674-909b27edbf73","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"GPIO13","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"8","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[456.5066525413885,332.4462975933936],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"de9b39d1-1e28-492b-9be8-7de288cd2559","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"GPIO6","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"8","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[454.62343403825975,379.73353808062325],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"e3e0359e-9bb9-44ac-80e4-66e3c1f30411","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"GPIO5","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"8","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[453.2046995733484,423.77942097649714],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"49914fee-a25e-42ff-ae99-52a23942b71f","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"PTS645SL50-2 LFS","displayFormat":"input","showOnComp":false,"isVisibleToUser":false},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"C&K Components","displayFormat":"input","showOnComp":false,"isVisibleToUser":false}},"position":[403.99739050000005,229.81236799999996],"typeId":"7cdc340f-5a26-48f5-bb1a-8e6e2bee0aa4","componentVersion":1,"instanceId":"101dbdbd-a855-4798-9242-a7c17a09d383","orientation":"right","circleData":[[422.5,244.99999999999997],[385,244.99999999999997],[422.5,214.99999999999997],[385,214.99999999999997]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"GPIO16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"8","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[477.05839877183263,158.1060918244766],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"07dde854-559b-49ac-80f5-aa8b57c2b5cb","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"3.3v","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"8","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[541.5573437700974,504.91648808548894],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"11263eb5-b485-4dae-b6c9-21c18e7b3a28","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"10000","displayFormat":"input","showOnComp":true,"isVisibleToUser":true,"name":"Resistance","unit":"Ω","required":true,"validRange":[0,70000]},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.25%","value":"0.25%"},{"label":"0.1%","value":"0.1%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false,"isVisibleToUser":true,"name":"Tolerance","required":true},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"string","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false,"isVisibleToUser":true,"name":"Number Of Bands","required":true}},"position":[157.22504875383441,170.69373781154127],"typeId":"72c75556-baa3-04e7-55a5-e13f447c8c5a","componentVersion":1,"instanceId":"72fd138d-67df-44a8-bd00-9e004d450883","orientation":"up","circleData":[[122.5,170],[197.4999999999999,170]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"YELLOW LED","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"8","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[209.0736813496403,329.16743830082186],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"5078f55d-6889-4bc8-828b-a676a5fdd005","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"RED LED","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"8","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[205.9570835169858,284.6440645205774],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"d430a89f-cf84-421d-97a9-6ef91b5385bc","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"2.81950","left":"65.30875","width":"857.41411","height":"544.91345","x":"65.30875","y":"2.81950"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_1\",\"endPinId\":\"pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1\",\"rawStartPinId\":\"pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_1\",\"rawEndPinId\":\"pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"219.9040000000_440.0000000000\\\",\\\"197.5000000000_440.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_1\",\"endPinId\":\"pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_1\",\"rawStartPinId\":\"pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_1\",\"rawEndPinId\":\"pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"197.5000000000_395.0000000000\\\",\\\"219.9040000000_395.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_1\",\"endPinId\":\"pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_1\",\"rawStartPinId\":\"pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_1\",\"rawEndPinId\":\"pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"197.5000000000_350.0000000000\\\",\\\"219.9040000000_350.0000000000\\\"]}\"}","{\"color\":\"#020202\",\"startPinId\":\"pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_1\",\"endPinId\":\"pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_1\",\"rawStartPinId\":\"pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_1\",\"rawEndPinId\":\"pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"219.9040000000_305.0000000000\\\",\\\"197.5000000000_305.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0\",\"endPinId\":\"pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0\",\"rawStartPinId\":\"pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0\",\"rawEndPinId\":\"pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"122.5000000000_305.0000000000\\\",\\\"122.5000000000_305.0000000000\\\",\\\"122.5000000000_350.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0\",\"endPinId\":\"pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0\",\"rawStartPinId\":\"pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0\",\"rawEndPinId\":\"pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"122.5000000000_350.0000000000\\\",\\\"122.5000000000_350.0000000000\\\",\\\"122.5000000000_395.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0\",\"endPinId\":\"pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0\",\"rawStartPinId\":\"pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0\",\"rawEndPinId\":\"pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"122.5000000000_440.0000000000\\\",\\\"122.5000000000_440.0000000000\\\",\\\"122.5000000000_395.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0\",\"endPinId\":\"pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0\",\"rawStartPinId\":\"pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0\",\"rawEndPinId\":\"pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"92.5000000000_470.0000000000\\\",\\\"92.5000000000_440.0000000000\\\",\\\"122.5000000000_440.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0\",\"endPinId\":\"pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_0\",\"rawStartPinId\":\"pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0\",\"rawEndPinId\":\"pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"122.5000000000_305.0000000000\\\",\\\"122.5000000000_170.0000000000\\\"]}\"}","{\"color\":\"#1a1a1a\",\"startPinId\":\"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_16\",\"endPinId\":\"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_5\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_633b310a-2a82-4082-91f6-b1a17256c96b_1_16_4\",\"rawEndPinId\":\"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"482.5000000000_455.0000000000\\\",\\\"557.5000000000_455.0000000000\\\",\\\"557.5000000000_455.0000315000\\\",\\\"587.5021750000_455.0000315000\\\"]}\"}","{\"color\":\"#1a1a1a\",\"startPinId\":\"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_0\",\"endPinId\":\"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_35\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_633b310a-2a82-4082-91f6-b1a17256c96b_1_0_1\",\"rawEndPinId\":\"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_35\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"437.5000000000_215.0000000000\\\",\\\"437.5000000000_170.0000000000\\\",\\\"550.0000000000_170.0000000000\\\",\\\"550.0000000000_230.0003240000\\\",\\\"587.5021750000_230.0003240000\\\"]}\"}","{\"color\":\"#1a1a1a\",\"startPinId\":\"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_0\",\"endPinId\":\"pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_1\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_633b310a-2a82-4082-91f6-b1a17256c96b_1_0_0\",\"rawEndPinId\":\"pin-type-component_72fd138d-67df-44a8-bd00-9e004d450883_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"422.5000000000_215.0000000000\\\",\\\"422.5000000000_170.0000000000\\\",\\\"197.5000000000_170.0000000000\\\"]}\"}","{\"color\":\"#1a1a1a\",\"startPinId\":\"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_15\",\"endPinId\":\"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_28\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_633b310a-2a82-4082-91f6-b1a17256c96b_0_15_4\",\"rawEndPinId\":\"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_28\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"377.5000000000_440.0000000000\\\",\\\"565.0000000000_440.0000000000\\\",\\\"565.0000000000_274.9981805000\\\",\\\"602.5000000000_274.9981805000\\\"]}\"}","{\"color\":\"#1a1a1a\",\"startPinId\":\"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_9\",\"endPinId\":\"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_32\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_633b310a-2a82-4082-91f6-b1a17256c96b_0_9_4\",\"rawEndPinId\":\"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_32\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"377.5000000000_350.0000000000\\\",\\\"535.0000000000_350.0000000000\\\",\\\"535.0000000000_244.9982045000\\\",\\\"602.5000000000_244.9982045000\\\"]}\"}","{\"color\":\"#1a1a1a\",\"startPinId\":\"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_12\",\"endPinId\":\"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_30\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_633b310a-2a82-4082-91f6-b1a17256c96b_0_12_4\",\"rawEndPinId\":\"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_30\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"377.5000000000_395.0000000000\\\",\\\"550.0000000000_395.0000000000\\\",\\\"550.0000000000_260.0023400000\\\",\\\"602.5000000000_260.0023400000\\\"]}\"}","{\"color\":\"#1a1a1a\",\"startPinId\":\"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_0_6\",\"endPinId\":\"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_36\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_633b310a-2a82-4082-91f6-b1a17256c96b_0_6_4\",\"rawEndPinId\":\"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_36\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"377.5000000000_305.0000000000\\\",\\\"512.5000000000_305.0000000000\\\",\\\"512.5000000000_215.0024150000\\\",\\\"602.5000000000_215.0024150000\\\"]}\"}","{\"color\":\"#ad0000\",\"startPinId\":\"pin-type-breadboard_633b310a-2a82-4082-91f6-b1a17256c96b_1_2\",\"endPinId\":\"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_0\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_633b310a-2a82-4082-91f6-b1a17256c96b_1_2_1\",\"rawEndPinId\":\"pin-type-component_c03fea7f-e196-404b-826d-0177413f616b_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"437.5000000000_245.0000000000\\\",\\\"437.5000000000_260.0000000000\\\",\\\"355.0000000000_260.0000000000\\\",\\\"355.0000000000_522.5000000000\\\",\\\"602.5000000000_522.5000000000\\\",\\\"602.5000000000_485.0000000000\\\"]}\"}"],"projectDescription":""}PK
     �)K[               jsons/PK
     �)K[Ȣ       jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"LED","category":["User Defined"],"id":"7c3ccbf3-d039-4eec-8ff4-6af5efd4a31a","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"cac5f02b-fb1b-403b-a5d1-1baa7913483a.png","iconPic":"898fbbe1-f190-4098-9ff7-64122b8b80b8.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"3.48889","pins":[{"uniquePinIdString":"0","positionMil":"5.72076,142.13630","isAnchorPin":true,"label":"Anode"},{"uniquePinIdString":"1","positionMil":"656.36076,142.13630","isAnchorPin":false,"label":"Cathode"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"LED","category":["User Defined"],"id":"7c3ccbf3-d039-4eec-8ff4-6af5efd4a31a","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"cac5f02b-fb1b-403b-a5d1-1baa7913483a.png","iconPic":"898fbbe1-f190-4098-9ff7-64122b8b80b8.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"3.48889","pins":[{"uniquePinIdString":"0","positionMil":"5.72076,142.13630","isAnchorPin":true,"label":"Anode"},{"uniquePinIdString":"1","positionMil":"656.36076,142.13630","isAnchorPin":false,"label":"Cathode"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"LED","category":["User Defined"],"id":"7c3ccbf3-d039-4eec-8ff4-6af5efd4a31a","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"cac5f02b-fb1b-403b-a5d1-1baa7913483a.png","iconPic":"898fbbe1-f190-4098-9ff7-64122b8b80b8.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"3.48889","pins":[{"uniquePinIdString":"0","positionMil":"5.72076,142.13630","isAnchorPin":true,"label":"Anode"},{"uniquePinIdString":"1","positionMil":"656.36076,142.13630","isAnchorPin":false,"label":"Cathode"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"LED","category":["User Defined"],"id":"7c3ccbf3-d039-4eec-8ff4-6af5efd4a31a","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"cac5f02b-fb1b-403b-a5d1-1baa7913483a.png","iconPic":"898fbbe1-f190-4098-9ff7-64122b8b80b8.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"3.48889","pins":[{"uniquePinIdString":"0","positionMil":"5.72076,142.13630","isAnchorPin":true,"label":"Anode"},{"uniquePinIdString":"1","positionMil":"656.36076,142.13630","isAnchorPin":false,"label":"Cathode"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"GND","category":["User Defined"],"id":"98d6e125-552a-4063-90e5-58c04872effd","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1cdb40d8-22d5-4761-8204-85ee5f97d036.png","iconPic":"9ee875d8-7c7b-435c-a3d9-92ac29f03ab9.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"2.37626","numDisplayRows":"3.61380","pins":[{"uniquePinIdString":"0","positionMil":"114.60833,303.64262","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Resistor","category":["Basic"],"id":"72c75556-baa3-04e7-55a5-e13f447c8c5a","subtypeDescription":"","subtypePic":"bbfae99c-8036-4c5e-89fd-a87441410720.png","userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[{"type":"double","name":"Resistance","value":200,"unit":"Ω","showOnComp":true,"required":true,"validRange":[0,70000]},{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}],"iconPic":"a262aa33-74c4-460b-b0ad-c746896f6744.png","componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Resistor","category":["Basic"],"id":"72c75556-baa3-04e7-55a5-e13f447c8c5a","subtypeDescription":"","subtypePic":"bbfae99c-8036-4c5e-89fd-a87441410720.png","userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[{"type":"double","name":"Resistance","value":200,"unit":"Ω","showOnComp":true,"required":true,"validRange":[0,70000]},{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}],"iconPic":"a262aa33-74c4-460b-b0ad-c746896f6744.png","componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Resistor","category":["Basic"],"id":"72c75556-baa3-04e7-55a5-e13f447c8c5a","subtypeDescription":"","subtypePic":"bbfae99c-8036-4c5e-89fd-a87441410720.png","userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[{"type":"double","name":"Resistance","value":200,"unit":"Ω","showOnComp":true,"required":true,"validRange":[0,70000]},{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}],"iconPic":"a262aa33-74c4-460b-b0ad-c746896f6744.png","componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Resistor","category":["Basic"],"id":"72c75556-baa3-04e7-55a5-e13f447c8c5a","subtypeDescription":"","subtypePic":"bbfae99c-8036-4c5e-89fd-a87441410720.png","userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[{"type":"double","name":"Resistance","value":200,"unit":"Ω","showOnComp":true,"required":true,"validRange":[0,70000]},{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}],"iconPic":"a262aa33-74c4-460b-b0ad-c746896f6744.png","componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"GND","category":["User Defined"],"id":"98d6e125-552a-4063-90e5-58c04872effd","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1cdb40d8-22d5-4761-8204-85ee5f97d036.png","iconPic":"9ee875d8-7c7b-435c-a3d9-92ac29f03ab9.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"2.37626","numDisplayRows":"3.61380","pins":[{"uniquePinIdString":"0","positionMil":"114.60833,303.64262","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Raspberry Pi 5","category":["User Defined"],"userDefined":true,"id":"a7ff864f-ccec-4557-bfc3-03323186baf4","subtypeDescription":"","subtypePic":"7be072cc-a725-4446-be13-eff8a797d760.png","iconPic":"d39a4f5b-af2c-4f90-bee3-bb82593c1b3b.png","imageLocation":"local_cache","componentVersion":1,"pinInfo":{"numDisplayCols":"34.99423","numDisplayRows":"22.55956","pins":[{"uniquePinIdString":"0","positionMil":"351.55302,2068.15242","isAnchorPin":true,"label":"3V3"},{"uniquePinIdString":"1","positionMil":"351.55302,2168.13792","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"2","positionMil":"451.55290,2068.15242","isAnchorPin":false,"label":"GPIO2"},{"uniquePinIdString":"3","positionMil":"451.55290,2168.13792","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"4","positionMil":"551.55281,2068.15242","isAnchorPin":false,"label":"GPIO3"},{"uniquePinIdString":"5","positionMil":"551.55281,2168.13792","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"6","positionMil":"651.55266,2068.15242","isAnchorPin":false,"label":"GPIO4"},{"uniquePinIdString":"7","positionMil":"651.55266,2168.13792","isAnchorPin":false,"label":"GPIO14"},{"uniquePinIdString":"8","positionMil":"751.55256,2068.15242","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"9","positionMil":"751.55256,2168.13792","isAnchorPin":false,"label":"GPIO15"},{"uniquePinIdString":"10","positionMil":"851.55240,2068.15242","isAnchorPin":false,"label":"GPIO17"},{"uniquePinIdString":"11","positionMil":"851.55240,2168.13792","isAnchorPin":false,"label":"GPIO18"},{"uniquePinIdString":"12","positionMil":"951.55231,2068.15242","isAnchorPin":false,"label":"GPIO27"},{"uniquePinIdString":"13","positionMil":"951.55231,2168.13792","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"14","positionMil":"1051.55217,2068.15242","isAnchorPin":false,"label":"GPIO22"},{"uniquePinIdString":"15","positionMil":"1051.55217,2168.13792","isAnchorPin":false,"label":"GPIO23"},{"uniquePinIdString":"16","positionMil":"1151.56594,2068.15242","isAnchorPin":false,"label":"3V3"},{"uniquePinIdString":"17","positionMil":"1151.56594,2168.13792","isAnchorPin":false,"label":"GPIO24"},{"uniquePinIdString":"18","positionMil":"1251.55181,2068.15242","isAnchorPin":false,"label":"GPIO10"},{"uniquePinIdString":"19","positionMil":"1251.55181,2168.13792","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"20","positionMil":"1351.55168,2068.15242","isAnchorPin":false,"label":"GPIO9"},{"uniquePinIdString":"21","positionMil":"1351.55168,2168.13792","isAnchorPin":false,"label":"GPIO25"},{"uniquePinIdString":"22","positionMil":"1451.55164,2068.15242","isAnchorPin":false,"label":"GPIO11"},{"uniquePinIdString":"23","positionMil":"1451.55164,2168.13792","isAnchorPin":false,"label":"GPIO8"},{"uniquePinIdString":"24","positionMil":"1551.55151,2068.15242","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"25","positionMil":"1551.55151,2168.13792","isAnchorPin":false,"label":"GPIO7"},{"uniquePinIdString":"26","positionMil":"1651.55148,2068.15242","isAnchorPin":false,"label":"ID_SD"},{"uniquePinIdString":"27","positionMil":"1651.55148,2168.13792","isAnchorPin":false,"label":"ID_SC"},{"uniquePinIdString":"28","positionMil":"1751.56515,2068.15242","isAnchorPin":false,"label":"GPIO5"},{"uniquePinIdString":"29","positionMil":"1751.56515,2168.13792","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"30","positionMil":"1851.53742,2068.15242","isAnchorPin":false,"label":"GPIO6"},{"uniquePinIdString":"31","positionMil":"1851.53742,2168.13792","isAnchorPin":false,"label":"GPIO12"},{"uniquePinIdString":"32","positionMil":"1951.56499,2068.15242","isAnchorPin":false,"label":"GPIO13"},{"uniquePinIdString":"33","positionMil":"1951.56499,2168.13792","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"34","positionMil":"2051.55086,2068.15242","isAnchorPin":false,"label":"GPIO19"},{"uniquePinIdString":"35","positionMil":"2051.55086,2168.13792","isAnchorPin":false,"label":"GPIO16"},{"uniquePinIdString":"36","positionMil":"2151.53692,2068.15242","isAnchorPin":false,"label":"GPIO26"},{"uniquePinIdString":"37","positionMil":"2151.53692,2168.13792","isAnchorPin":false,"label":"GPIO20"},{"uniquePinIdString":"38","positionMil":"2251.55059,2068.15242","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"39","positionMil":"2251.55059,2168.13792","isAnchorPin":false,"label":"GPIO21"},{"uniquePinIdString":"40","positionMil":"717.95778,108.80867","isAnchorPin":false,"label":"PWR-1"},{"uniquePinIdString":"41","positionMil":"818.17845,108.80867","isAnchorPin":false,"label":"PWR-2"},{"uniquePinIdString":"42","positionMil":"733.15282,224.52335","isAnchorPin":false,"label":"BAT+"},{"uniquePinIdString":"43","positionMil":"781.45206,224.71945","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"44","positionMil":"1249.94542,194.84813","isAnchorPin":false,"label":"UART_TX"},{"uniquePinIdString":"45","positionMil":"1292.04501,194.84813","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"46","positionMil":"1334.15319,194.84813","isAnchorPin":false,"label":"UART_RX"},{"uniquePinIdString":"47","positionMil":"1781.17844,108.80867","isAnchorPin":false,"label":"VIO-1"},{"uniquePinIdString":"48","positionMil":"1781.17844,208.95574","isAnchorPin":false,"label":"TR01_TAP"},{"uniquePinIdString":"49","positionMil":"2385.17826,367.95568","isAnchorPin":false,"label":"TR01_TAP"},{"uniquePinIdString":"50","positionMil":"2384.89876,467.51785","isAnchorPin":false,"label":"TR00_TAP"},{"uniquePinIdString":"51","positionMil":"2485.17802,367.95568","isAnchorPin":false,"label":"TR03_TAP"},{"uniquePinIdString":"52","positionMil":"2484.89822,467.51785","isAnchorPin":false,"label":"TR02_TAP"},{"uniquePinIdString":"53","positionMil":"2644.94796,2032.34816","isAnchorPin":false,"label":"Fan-5V"},{"uniquePinIdString":"54","positionMil":"2644.94796,2072.07957","isAnchorPin":false,"label":"Fan-PWM"},{"uniquePinIdString":"55","positionMil":"2644.94796,2111.80298","isAnchorPin":false,"label":"Fan-GND"},{"uniquePinIdString":"56","positionMil":"2644.78666,2151.52639","isAnchorPin":false,"label":"Fan-Tach"},{"uniquePinIdString":"57","positionMil":"1928.08302,351.86242","isAnchorPin":false,"label":"camera1"},{"uniquePinIdString":"58","positionMil":"2189.01302,351.86242","isAnchorPin":false,"label":"camera2"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Pushbutton","category":["User Defined"],"userDefined":true,"id":"7cdc340f-5a26-48f5-bb1a-8e6e2bee0aa4","subtypeDescription":"","subtypePic":"6b6fcb51-98f7-4a52-b90f-3140c0078893.png","pinInfo":{"numDisplayCols":"2.21979","numDisplayRows":"2.98791","pins":[{"uniquePinIdString":"0","positionMil":"212.24038,272.74623","isAnchorPin":true,"label":"Pin 3 (out)"},{"uniquePinIdString":"1","positionMil":"212.24038,22.74623","isAnchorPin":false,"label":"Pin 4 (out)"},{"uniquePinIdString":"2","positionMil":"12.24038,272.74623","isAnchorPin":false,"label":"Pin 1 (in)"},{"uniquePinIdString":"3","positionMil":"12.24038,22.74623","isAnchorPin":false,"label":"Pin 2 (in)"}],"pinType":"wired"},"properties":[{"type":"string","name":"mpn","value":"PTS645SL50-2 LFS","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"C&K Components","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"98e53ca1-f8df-492e-a5f5-3061f52364da.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Resistor","category":["Basic"],"id":"72c75556-baa3-04e7-55a5-e13f447c8c5a","subtypeDescription":"","subtypePic":"bbfae99c-8036-4c5e-89fd-a87441410720.png","userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[{"type":"double","name":"Resistance","value":200,"unit":"Ω","showOnComp":true,"required":true,"validRange":[0,70000]},{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}],"iconPic":"a262aa33-74c4-460b-b0ad-c746896f6744.png","componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""}]}PK
     �)K[               images/PK
     �)K[tM�G.  G.  /   images/cac5f02b-fb1b-403b-a5d1-1baa7913483a.png�PNG

   IHDR  ,   �   �E   	pHYs  �  ��+  -�IDATx��	\U����HΈ8O��`�$fZ����i�<[�3 �<#���i�f�i�x���+,��uD+Sq��TLs��߹{�>��p�3 ���s>{8��9��;k�g=k�k�`.^�X���g11����&@K(�Ν�����~��ݶm�^wuu]���U���ߗ��,��P( V?������c7m�����^+S�����Y^!�%XUk֬ӹs�wnܸ�}����~���U5A�"XB�8y�d��^z)�o��~�Ν�=W�b��ϟ��	���L���r���S\\\b{챲���F���}��m;r�k�`!D��|9|�p��]�.߿�r��iw��5�G�
�e˖5��%�~��XX���r��lxx�|wwwo;;�J�� 
��,�/_�<�WZFFFEM,���#?��C�6mڬLIIi�m���6��Y)$���&BK0��?r����3gN��3�b�+�1`a�����B�`�rX��سg�sM�6����wF<
q�����`ݺu��&B���Q?����W�:���Fw��}"����3<T70��d�C�H��h�`!D�J)+�6�qvv~����ձ�B�
ڟ�i,��p,�-��7o��%X�R[V�.]�=hР%۶m���W�B��޽{�T��,,M,�V)b�~���-Z�XI�TB��*�u�[[���eee��%X�Rȝ;w������T�|�2�� +	q+�\��rl%,�V)dԨQ�8}�jժaaa�Ϝ9�. �A,%^�"rLb���2S]G�'##C\B�b�`�RȊ�G�5x$$$L����9}�tS���jua��x>��<Ye�=t�25+s���&�Ǐ_�s��A�P"��ɓ''�Ȭ�����={�)��z�8�ҫ�-33iHಚ`�y[�l������X���I4e"v	CK0�`<-����!Y\�}}}�߾}�R�XU�X�0�]@ޯ&�޼y�
r�,}�\�4%%��SO=��СCO�ZID�58:88��	%,�o�����o��Ȩ��G|��`M,ama��<j����Χ�]�0ww��$���1����kMz^�"�%�):X�8q�,+W��4�p�>���m�`��E�+Z2���<x�{���ג��B�� �=]��-<�6�`	X�>��W{���9X,Hj����ׯ�"�5.Ǳ�޽���P����+W�T�2eJxbb��$NH�������\��ic��_m�,���*5�i�&�-+�n1�Xծ]�RJJ�krr�-�;y�d<�
	ܵ���`kmÆ�۶m����"��������7n��u	E�X�`�4�;v�>~�������Y�V���<������bbb|/^�X�^�� d��ʺm�k�|�r��#G�:t���4���x����XW%,�s�4OO�h��A)5m�aÆg�M��8}�t~TbiZZZ�{�71>>~&�l���322�43�&��wuu���̬	a��pyfQ�O+"�P���PD�k֬>nܸ'8�)�a!������&A�2~	�ZD�p,�]�p�ԫW����`÷�~�ݷ�z�7�qz|� J,L솪`�\Bi5VB���nnn^ N�y��ڵk�����8q��� ��Ob���)��r��+Vx4k�,�Ν;�X<٪��t N�P�* YdN�P"��իW�8v�X;�Z�@�����A�/6T�z���\áC��w��y������}&�(��<r��`|�*$X��P"�*"lqp�Z{Ġ�.ߤI�A�0888���7n|f	k�=���}}}��~��dIU�8qN�:%����X����r,�2##��&�HD��[��X�������G#��ȩb�����@K��C��Ç�Z�n�����[B����k�>�#vY��5_�͛7%�UB�*"��<==t��e�o�����+��|����r���D���aÆ%>��絋���B���� 7j��
���U�R�(���/�D��,��={v\�lٜ'�|�````H����h� K�.�v�̙�XW���ؼy�,a]���Vԭ[�"Yp�G�m�V��u5��v�Q��x�΂�����U�2��n�#G��'��ܶm�cAAA�ܨS�t ��dk�Gy�}���1b�֑#GZ��zu��$8�7o�ܛ�>�ĉ��jBZ�+n�
א���Sr��`ז'�*R��XgaEN�Xt�A��M~�ot'''�_~iCb�i�v�xyyE�K��c\��;))i܅�傛��X�[�ϟA�w4�s�5l0`�&��A?���+�U9��`Aq�!\�����[znMv���5�&W��{��˃�"ZG��Mbϖ��k�KXdq�5j��[�vm(Y+��Z/�R�iӦ�<��F�$��O��k]\�u�L׷)99y Y��dq��5ű+����YF���&��+�g᡿{
���g������SO=e������|T^%D�� ��n5p��:���رcג�����5~��uz�����`	,X�`jZZZc�2l%���D[ú�	]� \��-=r����د�k�V��+���fKK��n��X`9~�x����VĜ�Oc`�E�(beD�� �s�U[b�����_n�)S�$FEE��[�.xȐ!t��j�bW͛7�Ǻ��k�5����3�F`���~����ʕ�6� �	�����#����?po��K�<�A�Lm"���D���V�ֻw�[,V��������t׫̩S��:��d���y�޶\�@�(cpCO���7#nL�qӞ={j��G%c�|���_�pA��Z�*�q���Z��V�s�tss�� r��h��r���%~eD��n�.]�T�avu.��+͉�\�^W�,�F��Ϗ�1}��Dv-Q��\]]��fW�㚞}��I�vk6f�޽�u��Cu��J�5Ϙ1#3�-��v�f��>�[�����ť�^>�|M^�|d���"Xf�n�9�ҫ.[	�~���u�&\�p��9�X2aUt\���K����=!ZX�R-�t�����/���fkfΜ����7of��Ѿ}�n����F��E��$$$L�p��=YYY�� ���?<�ߩ18,,M�
"X��b�_p��{�ܹFs��]����}/<<��[�+�^�z��`� ����{ձc�o_z饯4�k׮H�����*U���*�+I����颂Iֆ�K�,�E���vT~$q�"�ecԉ���t�R]d���0�n����Хt�f�+�ť�·�7o�wYW��&			�e�N����V�X�z�~�����VߧW�$�z�D�'11qY��O�:�\J"X6�G9鑷�Ѱ����!�y����3q��8�(.���"�|�����k֬��O�P�G�_=���6�� Vd]�ػw��"�?���,`�֭9����)�D~��!$��5j�Hׄ�����H�>��9.C�N����$^s�ϟ�t����u�Թ\��d��^�����.$�����/��·���r(��,Z����}֮]���C��QԄ���Q�	�"ܨȘ�s.Z:.X��/..nZ@@@�9s�V���='�S���qs����k�׳m۶~}���mu�N/5�W``��;vhŔBUX
����-v+f+Cm��N���#�G���N�6m)	NZp)�˔yĺ�̛7/K�{sv�v<�]��cǎG4��#�ec8F���<4�
�oqI]�[�|�,zL�4i�����Gh�I��A���6z��7[s�>�6� A�<'�`Yu�g���~����υm��Q�����m�*���+V��������"驳�k%P�b���w$�1O�a�K�._#�UM��p�\���VnJ�҃u�� �6y��a�@�H�&�_�~Ę1c�}}}C\\\���S�
v[?��acǎm�I���xz>����p��F�°U�b��m2��u
[Y�0/�2�D��W�VY�f�h���G�^�������kq�k�6�f	@{ynzx�s�Ν�+S�����\��v�֭��y�O$�ú�k����
�Bw<���op�1b��G�oӦͯ�({\HTG�<y�DW�>y=<<��������0U�8���c!�`:O��dRS���\q����O��[�n����?<t�P����q[Y\�jǂ�� �۹!���<��w$V{lpm��P���0<Dϱ,�ϑ��bŊ�aaa��L��l�̡������'������k����4��k�����۷/��.C� O�Ѭ �C�1���~sVK4�I�!�a"�P���0���7#D	�Uff�ݛo���v�߰a�����9x�]E��)���A�q�rS$x��K�$''��q���؆�L�c����-�25j�X�m�����rww?@b%�+��2���Sm`AAD�V���իW�µu�־�/��O?u@p�KM�`x����j��R�l��wӦM}����_��R��m�.��{W�Z5�ڵk�p}\7L�D�������,�V9�x����5ӯ_�m�؆I�s�΍HIIy
�+��`<��65n��⥺�*j>[^;w�|���ǫ����N����������s(�>�A�ߵm�� ��6Mr@����ep�v��g=���#��zZ�M��Ȗg�C �qS�6��{���۷���矿��/~���J�=�u9��y���lW�]�]��pk��"X����ի�����_�:J�ݻ�9���@�Ըǰ N�piJ�)PU�R���޽�������v��}TTb\��oC`?)))�I�&gSSS�yf8w�-����w�&� �U��-��i�����:�����+xV
�MpjWe�k��֚����}��������7�<��d����+��&8��B~�ރ���o���"���o��,9bB�D����y��;z�����"W1��/�xU�P��yu"q^�k��#D��I��q��}��=C��ݺu�6(((��G�?\�}A]E��FK�,�IB5�q���薭	B�`َB'(v���'�>�"vHHH�#7�5�mǩ������j���P�G.q�N'b�D�/���ڷo U`�]ؔ��ӧ��{�?ި�#VG�>"X�0��D��O�8�� ۶m�C7�7m0ejOj�,4�`p`��QG<w���C�����~��J��W���O�>�	B>�`=���H˖-Q:�ߑ#Gچ���'''B3���W b�s9v�n%Ǵ8eB�����{�<�6lذ����)~�!*+��k�{I��D�v�}�j��P&i�t�R�իW��~���Z��G��S5��[J��[�S�N�>�b̘1IM�6�h�S�5A03"X%��:L�21((����8���@l�T�bhR�vF��X�y�����V����k�c�?��ȑ#�EDD��9bĈղ�B�C��B�|*=Ɯ<y24&&fnRR�Ȭ��J,V\!�r2'�
�cJ��{Y�H��q����'H�> W1`�ʕ��ҵ���	B��V�6\\\~��$�~�����6l������,wXSj�X]��2B��Y�N�J���S�N5�:u�r��|�/_1iҤ�pZ�o	�A�ѠA�s����P�|�֯_?�\�
�_!�����j!��P��Z�-�C�K��̘1cedd��������xI
�V)����wZL �+x���-[6����\�-+uBunT��N=D��0--����'.��ŋߙ9s�KU�J"X���y���K�.����0�֭[\!��\�T���Y���Q/_�� ݧ�����믯�W��x�5�	
�"X�֨Q�������hѢ)�]������u5�����H�ʤ�������������������x��,
ƈ`	��m�g��MV��;�3�D��:��EIMJ媡�g\��EKu�u~����k͟??<**j6	��)S�@��j�� �%�u�ԹL� ����%��ʕ�j��VbSp�X|X�ت�vY�h�:Y[d�΢�Jr��U�vM�eL	�	6CK�](|�]���g\\�4.'&n��UC�r�)=�v�Q]J����ى,-�+V�������(W)GK�'''Ĕ��MLL|+<<܋D��q	n������Z1Uu)Č��D��9���;���/���!]J%"X��������裏�"�
As�r\݁�`��W�G#y�ĊS �1�.~��Y�\ԩ�&&���G�p�>D��S�F�LZ�?�U���ҥK9��'�Z�O�8݁��-�h(�+���z.X��cƌ�gΜӤI���ʜ�m��Ľ���Ph�\)�[�bŊQ�*��;w��&��Y^p�F&v%���J��ӻ�T�����dɒ�gϞ��ԩS+�5k�J�Ϳ����"�%	4P|��d	�[��������AR�@ �RG%9���.�s�=F2':��'N,jٲ寚P"�̆^9t�k����CCC}N�>ݔ��p�#����6|e�;SS#8��Mf9h����Q\�|�8�ð������)�����ڴi��u�,� 1��D"	�+W�啖�梗��[X���BK몘兞��.��eOb9vժUc��y�慺���4e��Ir+�s�S�:
�EK�z µ�dXxx�Ojj�+����H1xB������=,/,!`k֬F�5���SRR�Z�j�k^�y��Z�h�P�H-/D�����k�شi�~~~!$\.$2e!,<*��A�jٰ��t �q�6زeˠ�[�>|���Ǐ��l��D.�]�A� V���`=D�̃L�5�
z~�nݺA���!�j	����n"ǹ��[j�*[H\��}�ᇃ�6lX�ɓ'�7o�z��!� 1+��4���`]D���Z5C��H��۷o=  �����88ϙ��.rҪ0Ws��4HJJ�ǠA�68p ݦrez���@��,� A�B�[6[hu�l}#""����Os�Ȕ�\�Nr�<�Ǡ ����PYĒ���oܸ��nݾ<q�����5*����]��D���"X�A\�B�Z\����F�m�w�~m¾��.�!. �RO���:I�c]x/��V�Z}�Wv�ܸ۫q#;C��"Xf�����Qo.T�S�`}t��&�/���.Z�����_!��k�޽�s�W.k�=�����&N2e�����j&�ދt�޼^�QB�{�8�:�ӯ��Q�yT�b��B��ɫze��?��C'��͓[y5���ӄ\����i���]�����G�۷�Y�ua��p�D�5�p4��۷�&������X�|���ʖћ2�w[��2��on�s��_�4�H`T�/������rY)�?/���7������?�gϞ�\/^M.�A|���i��ݾ}{uTR���9��C�8����z5,,���`����>��>��Ț��{����! 7���$8/�wv�����b\/L(:"XE�o.�<j[x��t��* �5j�#G�����Y�s��^xN����rK����8'�4ӯU2�-����D((|�j�_�m�HO�֖���C�܎�g��رcO��K�������D��ouT��8��e^��W���g�Y�꯬�4^��.\'�1য়~j=��O?��!V|��htmV��&��*��7��?�K��,���QZr��᰸��٫V�c�Ԟ"�;;�B�pm\�P0��|4��c�oO-6����K��M�׼��u�v�R�{7o���֭[5--X�y��!Tl����Hн�p>vA��_Y�(9u�1Jo���"�~~�^>!!��^�p���k�����e��z,y:�~M�`^D�����?'~m�"`h�N2�l^�\������OL��_����-;kX8�N1��yx�"�?\2�ڼH��C؜����Y����XW����BTT�GÆ礧���QY�r#KD�-9�?�~�r��a�v	q�����o�32�ƿ��W����V�f�陙���٫�a]�;n���gٹ�.�ۏd������ � ��<+�������N�R��
B�U�V�i$N�(�Vd�jl�pA?K�6�{�*�	�j��`>����~pW�ܲ��V����^�0�m��<�L;�1�!�Un֫�O�@�*o�"+��p�n޼����
���
�����-ĩR�J��z���y����cD�&����=n6M(]�v���{��y
c,\�t��2�;�/_����7���ޛ���^�gp��l�^��xX��u����̙3�(Nu�RF�͌���Y�դQ�o|��cVFF�&�ǒ�ZR$Nu<7n�I��CNM)x�81�����X�ة�ٝ��+�J�_�r����,;z�}��U��2?"X�́X]�x�VLL�o�&�P��Q��`�2~-�/��"��,r+�N�6YI�"##æL�����0���V�	���"X�M�q�F�ٳg�6o�|xVVVeN(�+[S\�"���v��n�Z�jg͚C珃�4u�T�u��w��Z�^�&X,�&�={���ŋ}���ުX�"b�e�i�-!�(��F�X�x��SMj׮}n���ú#�B��\]]+J*B�E�<�K`"����CBB�H����`� K���+Q�%��@;ףRgp}2>N�Z�NӹC�����ɓ�q�VV˖-�����1�����`��������i���J$Vv�~�G y�0P���=��Vj�
аa�3���!�F�� �zƍ���n߾]�+.�,���>}�ITT�������u
�$O�2���z0<�X�Z���xU�T��f͚���H��A�F�����+W�O�^�B�AK�|2&&fnӦM�a��q�'ϽS�_r���L�G�X��|��#ӦM[2~���!R��,��U ���J�`	f������ڷo��q� �SS��j�{�kLq�fu�N-��b���|кu딹s�ƌ92Im�ZX��Q�T(8"X�Yؿ���-��С�՚�n��"�n �9��cZ�#x8YT�fΜ�����7c�!���P2��DJJJ뀀��.]���VS��[N9��9v��90olU��݃E���HB����!C4�d#�e;ɸϏ;p�@{??���Ϯ�����"Ǚ��
�X�� V��e�Ν�����˟A�D�J"X�� �����Խ{�Ў;fDGmd�뎎��)�%��A�x2�>�gz�9 �s�����ꫯ~Fb�	�,�$���z������_�$��s'noƖF�L��͹Xd�C�{t{���=z����JJ/"XB���۵kW��E�q"'�]85f�mS'��9��+x��===�{���-�k֠�T�+ֈ`	9�cǎ>]�v��w��.���,ܵZmg�dϜ�ʔ����am�8��߮]��uh���`	�n:	�+AAA���@�N��kRnӮVK�����w�8��y��׷����v���_d�i�`�V)Fm�m۶W���CH4ܸ&�)s�غ�Ɯ��q,5�؍�.7�����ߊ	�m۶=�e�MrC�����Xm߾����O	U;����1e0��<�����!X+�� ��-���F�Z?eʔ�:u:�y�f)),�V)��,aY}���oFGG���k�x��q���2ˍ�[V��%��6��C��ڬY����"VB~�`�p�Vb�����-[�MMMu����tuR2ϣ3u��z���իW�߃cq�
���qo����!T'?��M
�V	b�*11qdxx���6�@8��¶:��Sؽ����%U�j�lw�r��Y�nn�P����+J(
"Xf ����ZTh�NB5����+--����I�çV'(h�1��1�/33��L�:u���gYTg�����`����nQ���F=���$T��L�ޱ���X��Iyď�����X$|wQ+���/�A�����5A0"X%Ւ%K&�Px����7�ߧ�S+|r���Zל'7�%_���r3ƍ�*�q�Ʃ˗/��܈`� HP*��6lt����S�����	� U�\����kԆ�<��EM�0a%�?-66VK!�����	X�r�Jդ�����՛{�ҥz<�g\;*/8/���c��mح[��K�w�����EU�n�t-M,��#Ċܽ*�W��tvv�s��ͪp��JR˼�Ң
� D�}��0�b����T�X���Y���|���������Z�`َ�_�v�ڊ+��h�b�Wǈ[PL���kJ�"X,D���¨����{:88dN�6m����"�+���� X,3`�ܢ��̚����6l8��9�	�,L�3U� z(>��Z�j�AU�[o�_�z����0Ml�V1Cͣ�~���}��	$ZN�~��>�}��3�^�beJMuN��d�������_�Z�k��ޚ ��b�*==�nBB��F�ͽqㆡF�Z���鼄�QG�L��΁u�H�_:r�F����&�,���9M\���θ:�S����y4�z�޽r9YG��_��'�7�u�e���}5j��c�ܹs��y���������!�eؕj�Ց#G�X�f�����O$Ѫ1Q�z~����� ^+į�CBB����Qݺuo�hi�P\��0�AyY?�Ο?�xdd�g�}v��۷˩�SjT^���j|NĴ��x5�9U�F^���^@U<J�L�8Q�����`p�9g�c�G�F����س� 2�U��
�PKè������ի����W��I�>@;w���G	,���=���q�<��K`j�'g���X��	q$�*��j����C̆�̱"X�˷@���!Q��q\��̣~��5�%^pbպu���-3f�j��D�,B�)/T���0&�� VC�(�,g13%��ix�.V���,۪U�����B������رc5Ax���0\���%lC�`qq�5ŀ-2v�b��sK��͛��;hР-Æ�������1N�� �LW�pٽcԺT�S$�:�6�~��͛��ol%��4B�D�ƨ�Vj<�S ,����a���ۡ�� �>}�� ��*+�$"�ec�eĒ�q��Y�N��Cf�k���9ĉ� �P��̭�������
��r��nݺ�!�/⥗^��	|�0-%,k	�w���ƶX��\�=���"��Jm>*�	,�#�,\ ��?l����^^^�ݻw�V���4"�U�:V<���s�=�'66v����!*A�"X6Fu�����{���opǎv��A���2��q�='ժ��ׯ_��!!!�nnn�6m�d�	6�)��!�ea��q���ѷo�������-[ݲe��2���!"g%D��C��_��'�؇����;�U�V'�<*�U	B�`��<a!P.�&L�xΜ9�O<��/k׮�~�XU�I�-ވ`Y�d���X6k֬�...�%&&�\�b
�M(���1�s�\    IEND�B`�PK
     �)K[]�I��  �  /   images/898fbbe1-f190-4098-9ff7-64122b8b80b8.png�PNG

   IHDR   d   4   |l��   	pHYs  �  ��+  �IDATx��\X���AtrV4
���*��B��dD\�1gr*bf�7�٘��h��h���CJ��Ȝ�a��o�	I*�~����z%���}�}]��~�����ݿ���}?���(GRTT$&N�(,X ����ɓ'�gW�T�ȵk��\�~]�w)����D��K/	wwwadd$���ZԬYs~fffۆ���?ċ ���Œ%K ���*�����<8%77ל�*V�X�B�
���@�w1x@���E˖-E�D�f�:�������}aaael�E��nݺ�}��V����a#���8O��X�3���jIOO)))���S,�q�޽{��_}h�!��B�ݺu����䌙�ٹ���7�����999��Ũ�qe̘1b֬Y�XWWW��{�VĽ2����BW�fgdd̏��<x�����s�0���mܸQT�^]t��Q4nܘn�{���a����p�o�����j�*���o���7�x#JnH *W�|3=7++���ݻ�r|ZZ��裏ę3gD�5�ʪ���������Y\a��	 QQQ���T��ڊ~�AQ��Ⱦ}�ġC��rzB��prr
ı��C&#&Թr�8��������b����c�����ܹӈ�F��k�b쐢	 ӧO7n�`�-Z�P�͜9���)�3^��TX�T�������������g�fǎ3ڿ��Ð(6��N�:5��e�����٨�MY�G-Z��	 �[������_���-8��D�������-,,���ť7b�'rQ�~�����
����[�r�0`���3g�B��.2/Q+�b��̵k�V\�C��4x��+Z�&��g#�V ՜q�ĉO�qG`G ���͛+,hРAbѢE����Hѽ{w�t�R�:u�s����m���X�*�����СC�&$$�!� 7�ƸDk�w����Ey�z���،p�n�&M���`�BK��8(��(';;�h�t(fd�z��av.������޽{�k׮��5k�ѣG3��"x7��f.��k׮��jӦMd\deY�5Q�;j �/�|�n�lű��W^�ˣ�������q9��R��X4D�"(T���0�aoo�-�	��Ocf*�����ťK�D||�q�Z���:��x���d��?��!@�u�&f̘!v�������+��`V_����f��x�X�f���]��K���W_-E���?ʯ�2�z(��K;	�$�zDժU��a��:��u�={�<2���/^����2ڴi3۶m�a}�񬖰.S�u�_Z�Edr�,�E�y�T ���z�j@ff�`��ժU[8iҤ�/��2s��)cE�Ν�*0�-��l�2��s��R.���ӧ3a��m۶pI�cPF���^ Q�P���7���@��3 �w�`�Ν�Yv��������SR o�`}4;�e��]����_9������7@(����B��P�t����˗���#[kee�5j�ZL\\�2�GЅQ@u��n�NRR��b��f�ڵeQRȬ���f��NƊ��.d�c�8N@p�Ym/3j9�����ꍠ��_���2O V�!��JFOz��Ԃu܀u�#�ٳg��"z��@���ƍ˂|:dȐH�! fh��F���z���0�`5:0�]piJ�Ҿ}{e,��͛7��:��[��/���D�A].�"i�~�ܹ/����lذa�8 �H.<ɸ���_�t0��ȶ� �.\�=66V̛7OL�:u����J���W_}�\YE�P8�'L�����2AY �X�82.ȹ� \���D��Xs�)S�$��ҹ�|lK)ϔ1@�1TWl߾]����>�|Xddd�l 3�����V�&@x�$Å}������X������رcEy� D���s-}�֭dT�ȰGGG/m�W����.Y��3\�0�pe��av#	���%$$�g����W_	�,a�bP���k�68��B�9��(�$����{�y"o.��2��o$�^ ���+���X���?*cBCC����K�eHA�`����۵k'֯_/>���\X�
��X_�Ċ�k��YL�j	`V7h��0����=���cfO�����%����@e�5����k�pQ��unnn���&!�x�"���6 ��D�n�:�lAϞ=W���ߥ�p ,R[�>Ek@��o`I��zԎ;Ļ�[ ���lpww�0����C����|� ���A9��� \1{��5���䜨��2���N�&�a�nH6��l0��4i�9==�Ӊ�H� ��`l�@�5j4�X�"@~~~9,�h������(����Q��Gi���Jn�*9;;���W�3�X9������T�s����#F����<$�y��0&�. �HM���`1N������Y���L����a�K] Of�E�����4a C�	Em	��Ϭ��u{*���J��Ջ����lժU۳g��w�
���x%���F��L���(�P��L�{����~���u�֥���t���#---$##��_�KUoZ���^u�����\�G�̄�Y�f��y�=�9r�kvv��_]+��>�M�?5[�Ǐ4�kjp�����G X�Q�F)����u`qeȽ{�j>����'�z�������y?�@����%|�F�z<V�EXP����
�Uع*�֢��z���������A ���B�0�433c�9c��q�jii��|�Y��Ɛ3��!lD[�lYE��+��ZY7��ѩS''$�SRR�srr�K1$�
�^���1�g�%%%� ��=16t�d\\�]�i���<��8qrrb�T<�2>m`�������(}�����������ݻw�r-K�(���n��G�������KHH��
��"��){ô~o�ܔN(T*A �e7$K����� "055�Onnn%�+.�<�� �5(xiӦM�u]�Z�<K�[�Ii)7�����������i�jժ�w��^�*�/-����
[�<==#bcc/qɗ���#���, RA,]�9R��e�믿�
ǂ`= ݠPg��:d��G����Zs��@<';���ÕM^o(b��Pq��L�0��'�|�u�6`hA��Q�|d��dPpMp�"�o"""���F��	���^ڀw��\_R��ص[���O?��������	�Y��0���t�gϞU�w��EI�K��f�֏�z�)Kjiee�lZ����ã�8z�hg2Aij0h�N������7zΜ9���S�
�l��cy�,�q~�A@���� �bC�A]:����q��,�6m�����(�0RYC�O#� R:CVI!��@�h����\K�mԯ��]������lZ���.{}iA��}\n�U�b!R٦���7�
 ��m�Vz�U~�E �#����K��".�]���+I!_��X/����\״�4?��2�1�@췵���=|^HH�sX�B��0�I���K�ϯXV�/�X[[�!ǎۈ��~PP���[�V��&�)zm����acc�\�n],g3��|��eGGGe�<88X�Ȣ�Đ�0� ��^�~}�����1;�R���^;�����5 �YH��^ ה��ࠃ�w�%1o  ����믿ք����ꭰ�a��Z��|�o߾$�F8f�l��k��7ʟ�N"g���*    IEND�B`�PK
     �)K[�wp�&
  &
  /   images/1cdb40d8-22d5-4761-8204-85ee5f97d036.png�PNG

   IHDR  �      ��֗   gAMA  ���a   	pHYs  �  ��+   %tEXtdate:create 2023-04-18T17:15:54+00:00SMK�   %tEXtdate:modify 2023-04-18T17:15:54+00:00"�=  	fIDATx���!�Va���1�l�tW�&l&�f�=�Y��`uF NW܁#8�~��2s��<�N}�KߝB$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)�/8�{����a�$_�~^t�a^;'yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yHYN����qr�݋y>���y��r9�WC�ݫa?+����C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C�r���-��.����`�<�!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)�L��<�i���l�6�8�n������f��5IR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR����? bw.g�����9���<pM���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�H~���p���u��$���y:���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E��8�w�q·H~����-$yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)�#=Ng    IEND�B`�PK
     �)K[!��Ů  �  /   images/9ee875d8-7c7b-435c-a3d9-92ac29f03ab9.png�PNG

   IHDR   d   �   ����   gAMA  ���a   	pHYs  �  ��+   %tEXtdate:create 2023-04-18T17:15:54+00:00SMK�   %tEXtdate:modify 2023-04-18T17:15:54+00:00"�=  �IDATx���]N�@@�� !Q���5.ـTg,<;��r��%��z�N:6��0��Ch�1��Ch���ǲ<"�ؕG��U�Ǻ<o�&�3�?"eL��s�?G�G?9�i�1��Ch�1��Ch�1��Ch�1��Ch�1��Ch�1��Ch�1��Ch�1��Ch�1��C�?�-E�w8�%��>.{t��.	ǘ�;�k�2�2������#g�"�*����;�3�KJ��:����o���א.6�*}�v�zju}�.n�&�O�'�aDR���gxA�1��_�ԫr�|�����MK�2���b���:�C/k�u�Z�+���m�����t���.�ʧ��qV�޵�lخ��O;�w�/j�m����ȯ`�!GƮŚ�RC�Y�]Y�|w-��M܎�g{�Y��k5���9rd�}��}���y)����>�4#�/��1��Ch�1��Ch�1��Ch�yQ�K���Oz    IEND�B`�PK
     �)K[�c��f  �f  /   images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png�PNG

   IHDR  �  �   ��ߊ  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  a�IDATx���|SU���M�M��ޣ {��Dq�����~�V*�~���(���(�"{�Q6-�-�M�{�'I�M������K��{onn���cU{�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!@��-[a츱�aC�5?�q8�^ݺ"���0�
�"���l�a���>C��p���Oo��vn����"��mE�9F�1\���?ۛ�����(:���c�X���_wlP(�ʔ{���=��|+��#}�Y��mo�w��k��]�o�������?�O�0�?���'�Q���W?s��3��"Sڶo�dՊ�}�I���i�f����gf^�t8Z������^d�g`���>�n�q�0K���k|=Ϗ���5�1��}���I0�p]�y��U��'3r��~'_{���G���ߢ��h������1o��v�#�����޵{�I��z�}Պ�ged��x0'""��!;;�߁�������t8�ADDDՎ��4���N����E�l4"""��L�����QQ���ԿTP�UK���	���sn������BDDDՓ}����{�������H/�=��|!'""�c�4a��sh׮ݔ�#F���u�}�?_+.q��p8PPP��o�O���m+�p���DDDG�}ǎ툯0;+k����C���PA܉��\��+z��I#<r䑓�\y���O5�Q�?�^D��R]�]R<�5k����q֦=11Q�s�*Yǖ�Ull,���0�C�Y6'"�`V|֠g�HKKS�o����T���Ύr���������GXd$���(T�:����=3+Y*��D�~2+3K��H�h#"���sx���_����`:͈�����O��;r��"""
f����6.��p�)�ggg��oDDD�����R�7Mgx�'�����"""
n�Cii����p:M{�'��]��QP3��SSѼE�8���,�3�:gOݟ�F��:�������y�
�DDD���";+;ơzI2�kff&���(��j����H�4�L��at""�`&��:���K@/3�^�a�Љ����nC����E��J膻��0���(���*w�^���(@VV���(���*����:��D^^>���(����p�Yo`� ��;w@/;�����FDDD�Mr�0��mPP�ϵЉ����iB��'ԭiՆ.������Q�V�%""�Qt/w���^J�&�΀NDD����m6È𶁴�{+�Qp�/^�T���t""��g߾m�*���6�Q𲧤�H������]��1�'���i��*w""��g����m*`��r���/��Ä�m�����NDD���3��G@g�;Q�S%�Æ����˝��(��3�����G����ΐNDD�Lس23��i�I��S��)U�ge���'{�3{NN�
����%�;Ճ������zdDD�i��K�DDDA�T=&&Ff��Н*�;Y�NDD�L{xD�t�S�:M�~Q��l6;|T�;�&L�Љ����=L��*w�Su"""
^v�a�ax�&�܉�����0�QN	�U�DDDA�T�\J�׉e���U�DDD��.K�|tV�3�|�i�̽t�U�DDDA��%���F��8tV��rK��U�DDDǀ�����t�K���˝��(���K�z���X���(��E�{	��7���t�,��ʝ��(�ٝO	�:��:űʝ��(hI����4�r��YB'""
fv��a�iz	�n?7�)���(�ٝ�sm��NDD��r���SQ�n��^�n��GDD�쐕�L��T07Љ����)U�J8|�r�Nq�DDDA�n+/�K�g@����<����@=?""�F��0;�*��乸ҵ033ii��k�.$'�@jj*>�����9	�QQ��S�ѨQC4k��6���\���1%>�|��%rpq��+�*3��?V�Y�?���Eb��-طo/<���<W�C=��,|��\`�!6&u��C�V�ЫWO0 }��A�&�f�1�Qȑ��i[�I@���p�{�W�܌���X�z5���;�:��V�ޯJ��(��Q�w�{�>)ͧ�Ė���/s0i�$t8�#�=�\|���ܹ��v��D$<�����pU���Ʉi7`��r��s�C��\�U�^�x1�����n�n٬��E�ۆ�)����`�E���Oq��W���GR���yv"��\�g.~��w|��g���;п_?�i`7нN��¹�}�\�-[�b����Gcǎ�p�W�����=轢������i�O��P\p���������O���u����拓�'�S��o�T!����>���2>�͘����3������_��p���T�Y���tf������ذq#��nԉ�cP'��'������ix뭷�|�2]�Y�^�z���'��2���V�{!�Pz^�0���*RS�µ��Gݷg��g'a��Mw���������{���#R�۟���#G���x䑇Ѡ~}u"
Zy���7o&��f͚���8��yHo���;�1��&��ޔ�y~&M�\�f��`�
���hܸZ�h�:�E˖z8Z�*UGGG#7'�z8ۆ�n�:lݲU�TU�[�Z�QV�a����HOKǨQ#� 1�A������K�,��߁�����Qi�tn��lC�C�����g�><����!??�oF׵kԸ1����3���&M��v�ڈ�{o���b�ʕ�a�:�~�:w���Gf ?/~�$��'�@LT�:�Ca�^��,���eʐ�0���or�gf��_�G*��`���9Q'>�>n��V=��v�Z�ϖ�|/C:�5i�H?�~n��L�<S>�\��S�5��s���[h׮n��z�~Y�(�2+&K�"��n�f9U��W\�Á�U	x���s���Űa�p�9�v\-�_+Ƴ�L�׭Kg�;��|2��֮�ù�J������ѱc�ؿ?K�DD!Nt�s����!�{Μ_���~�2�M�!����#г[7�_+O���/�	u�b��aX�l)�36�6��ѥK�� "�P�c�i7���*w]-̀^�n�ꫯb�d�z��L����p�Wb���hռy�Kƞ��u�@����~�H޶�����{�	�_xK�DD!ɕ�۝�i���q����0��)���_Q����p�����FTI0/N�}�Yg�����ǟ@���(�/3p�@*�y�m�4` ��cP'"
9�����rg��#���,F�9Y�.;ѵ[�G�M�VG%p��,2����/�L񲕁?���?���%]""
I�L�곛�k�Ԛ]B����i_c�jo��L������ރ^=z�R�'�N݃~�os�o�X��3��0s�L�{�DFDT��y�"X�X���x�����X]��:Ne��.��� ״������͞�}���[8�2{�u@|�ٸ��K�ɲ'8�w�{���O��������m=�c���xbP�p�ٟrss�����f��u&"B=�ߞ��y�v����y���Cn^���OV}���a+���N�[�8r��!�1�(ǲ��V�Nq�|����EFxȹʵ)p�>[u�rm��ץ���u}]�����OC��:����9�?���"��\}��ˌ���^��Пc�{�hU��)}>޶�R�5RT�y�s�C~J�@~�V�,�[9C�����57"��_@��U�?ϙ��+V�ۭ%cͯ��zԍ�?�7�/&:�^v	�M��C�0���-lطo�-_���Y"v���X�vV�Y��6`��]f��S�P�,�B�Z�ШQ#�n��:u�q�uD�����JZF233��]ۺ		:�*�>��)�f���X�x֩��s�N�I�##"�{hѲ:v�^�{����k�}^ŏ�r�*,Z�k�5۵k���t@����36o��{�@��]о];Ԋ�����u�8��W�3K��t�	�H��r��!���Q�X������u���lչ5m��}ջW/���u�9��a��5X�p�>Ύ;�q$C�����M�4E��ѭ[7$%��k U��{2��3-=[�l�K!�9n۶�))�����C��(�OL�3A��E�ΝѦMk�V���~�:��.�����MIJ�)���+T���6mB�>y��zK�D��f͛��,�u���㐘X��ZT��gVvv���}<p����_�X�����)�T��21g�(��t���k�8t�(���S_om�&���O<�R�>}�]}�������֊����m����ޭ{w�P��螛�J|���f̘����[�nEzz�����u^��t ���x�s�98��S�P%���w���x���٧��U8r%���5l�/��2ڵiS���C�o������
+T�g��>އ�";4h����õ�^�A�����8;U��n�����/�l�2���w/�k����(u�p�)����N>�$�R�ؑ^�/���<iR��r]d��_��*Hz����ᇙ��/�x�b��>>_�͎z�����5�\�s�g[O��J��`��F�ܰdrd�$���q�#T�T�9���u�	�$xUU��\�M���5�'���X�d����Hp�uT�.�6P�]O�ё"��*�W6�{�U�~1#G�ҁ�0��j�L�#�<Rbd�<������ս>Uw�MNNF���zoR����Z�.�1�sp��#�}{���� ���'��o��H׌2*��ґ��,X6�����?��v��#����.�С�)��^��C�`�l�R������;�ޱ�A.ǭ���*�4h�=z�K1�tP���>��U�ɫ3U[����{����z�g����t��.��c�JXd:ܛo�Y�ʮ'� ��%�ϕ�X��$�9[�
y���N��r��z�8�ޭ2�|��~��^v)U�gR�ve�]�b���ٳ����:���q�*w{�6|���0�Ǚ�Zɇ�J�͎��T%���_��u���<�+�ȿ����_�sGvv�_�+�lʾ��5�����y��ǟxݺv-���I�����B��Z�'_�.w�ځi_}�9?��ŗ\��{I����'g�k�|���z9ϕ+W�i���-�����nՏg�T���p�������KGb�*����?�{���K���Uk���̾R�����'[[��>'�dIAa����G��o֙)��L��M�����Z[j�֬^�u��T&��ge�ԯ���(g�pKU0߽[� �=�%~�q�I�������5�گ�GZ����[=�m؀�^{��9N;{$�6%������/�E]�r�Z����5�m��֩��,ǘz� ^U��7����}(���\�;=���}lٲ�����]J������7'��^��=�ܯ��5sm�?5o���ά���:v���)푆V*4u��p����N����|���f�?c�u�!�_L�[�n����|��"�>� /���]ŏ��VJx�n�\��cǢo�^��r&�9�UeXe�sU�-//��<{s][ɠIFsŊ�駟�裏�_����2��-�S�-��⟩��]x��gT@��&��̊ٵ�̮Z��?���H,���>��I����6��x���r�#����D�Х�2���>���:wB��m�Ӗ���[*J>�9*Q{z���믿�^�)��2�J(2���ч�R�J�H<�!C�v'T�%���'�x����d�k����~����@?���B����3�{5j��4dee��2?E�q80��oUf-�Ox�<�$�*�9
o��ffT�|ſ���Gzo�3�up��8���J�/�_R���>������O���$}�+S%57�F���Ƕ-��f�x��r��0��iذ~=�}�\tᅺ�_�SXO���/�£�<Zl�)��m[6]��������۶n�NjA@�����:lM.��t�t�2[�зO�׉�:�\jf���C����໻����m���WJ�Y��d��bX�w��_�h!��^�����_���*ڋ�	Z�1�w����a�B^���t|߁�'U
�4q�Q��-,���1a�J�=U�9�����NJ��= �r]���1��W0��	�ζʼ�������yx�����K/�Nco��^;i(��?��@���u�ȑ#�h�#!����F����9�[f��zH��������|���ū��s��z�
���zg㪫�
�gYڌ�3K�b�c���+�������Ǚ?⥗�cܸ�������eR:����ǝ�Tk��g��Ѝ�bz͹xť��`Ϟ�^����B�.]t5o(]!OR4��Y:t6o� ��ê ^�~��8ӻw4k�u���UT�h��]z���˖��]	��=gö����Ï�k{�E��T�ק�~��%���#"Ѵi3�B]Su���7';�R��Ҕ�n���VS�JЎ||�ɧ8���|�
_/�]	hLl��h��m�"11QG����uo�;v�;�Yg|�T�H��E_�.�W����=u�4LU%9W{y���D�=M�4Vץ�>o�$��RSS�a�l޴I��[_W�2L�:_r�
��0�L0w]���u�4G����u��n2�Jz��]�V]�dx_�X����(��N8�_�������ȑ��v� ���N��B��I��K�.�3�����Qڵ7oެ۶�'|��C�.Fq6=���=�;�^�I�$��t�2L�<����\ރ|O۴i�{�K�HG�C��r�򹦧�y9w��LӁ��}s���c��A>�G���}��/��\=�7mܨ�[�d��%�ף�t�S�֭[6+��)s���2>�����ak2�H!�ک��H 5��_�|9�?5��`�Db���T%�W^y��#פtu���ԗW��M�:����k�Nx�;�oÓO<�F�h�8Ce�Ru tu�+
�R��ۯ/���J�v�ih�����̈;)q�P�9����oM�R�1�f�Ϟ{n֫���]7�
�u0��3p�:N�޽Ѥq#=��s9���6�k\�����}{���#Ìf��:��^��"�>R�s�v.
�a*A�ޣ7�P���[�j�;W���W�dΤcۤI�����e�	�34t�x̘�طgRS���v":�N9�\}�U�qӦMu	�s]dH�֭��ݷ�����W`���"C�O���}zW����3�ǘ����yp'��o�駝����,���!�1�S��߅�����Y�,2K�s�{]VN����y"����}��ΕΠի� g�u&.��b=�q�ƺ7���zA~>RTfm��%�����H�Qِ�o�}�]�pB=����m곸��{p�-7���]���;u������gj��Q#1��u?�Lɐİ��?��kf@�R�+���D6Х�P������*p_Ub'�|*~�a�q�@Ĩ���'9��x��W�������6g�l��X��mX�z%�W	�۪�Ѩa�J't�P�\��T%���;q뭷��JPQ�L�p))�҅<������>V��t�Q%�����[���x��Gq�E��P��8R"�ݳ�w�'��?��*SeyUR��N�m\�а�8T`�*�G��"�*�ȃ�Եi�Jp�+c�\��-[��u-q�
�R��
�e��B�u��l�kޢ�=4LW97�_��K�jת���ҹ���N�ñ��?��IUb���{�͚4���^֬߀ѣ�ww����'�n��s�mh�2c��:��&������Izʿ8�E/�(ٰr�r�S�O|�Mԫ�P�{]�냅�Q������O�Ї���멈s�m�y2��|�q��aʔ)5r�:�����$C�j�9��nE�Bf��Gq��Յ���2����4��>A�I	��zg�'�q��ϬH�Zž�b���u���1}��qc�}˻C<��&g<�[��c�=�i_M��8B�)�|�ɧx���T�V�6j�Q�G��7�Ꜽ���R%����믿�vxz���T��^��K�DwZ�VaoǑ`0d�`]���۱g�.��lܸIWG׫�$.֊�K|ݺ��8����I����[Ǥ$<���X�n}���H&�ƽ8�{��1ͅ-���?U�1c���nƖ�-�c`��d=#�t���a�ĉX��[�թJ��1b�H]����ɞ�V_]O�II��V�	V��3f`�*9ߦ2��Q��J��u�_��T�3�9?o��!�Ho��]Z��~oSKK��|��:��^��X锸��Zzj|j^�9bz.w��멚�)N:rI��+�['P2�HL%&�6�i�ܵ��.2K5�u7p� =L+�]�#z�����J��t5���H{�|�ǨK/��\gW{�C���]����ݯl'��I�ᤷ�*wk�.=��`^ѡ���:^t�:�D�g=6X�z�J�+��;�w�q��ů"ץW������1F�t}��H�[O<�.8�����{��N��T`�>��C�aݺu8EmW���]���-��V�e��O>����+0��g���L{����t�{�+6��hˬ��z(��g֥〥)�|��a�葅����h*�I��K/�K�,յVs�H��c��	�N���Ց]���g��m�vM_d�p/SfVWs~��ŋ�[0�j��숃���V�ǞxLw[�'�([)�l~��ttx�� u��8��tӍ�ڸ��A�L�������mE��ύ7݄s�����9IIpР���O�x���1t�=iK'��֝�RʖL�ۓ�Fj�>x���J\~�e>k,���*�O�4��C("7JG+����S�#S�Ju�Ν�U���|�M�A�n+̋�Ƌ/�Pw}a����$C}��1�����Nt�p�Zb���W^#�j�G�)S�m�U��y�f�?p $k,��Ͱ�۳�&��KG���l[�V��P�i)��~��7�Y��~i�'�T.��SN�|;�����}�}�a���k�������s7�p�n���qM=%�u�]W���:w�&M���`��G'Z�l��.��2:$�~b}��f���A]�&"#�����)�Oj�V�Z�:�y�xm�>C�u�Ǒ���w�5)P����蒤�NS�*	����2��:wŭ�ݪ�D��.���o���f��.�+K��e:��^�\���0��$��a�k׮���B�{��]��Cꚻ:�ѱbJ��M&a.GMkC�_:Qe����B�+�ۄ�y���$\q���L��OI�.��=��?�:�X�b��5hr�9�<����uĀJ�엨J;�u@_�u�SO;�U��� �p��z���L��U-��V�[a���+���ؼE/S|��s��ǣg��*�JB����m�uQ��^�s��Uj+�2�aa�ͼC��z\�ަuk�{޹z� ��ҿ�.�M���[�5h�Hw@�L�kO@�*yw��	�M�n����̬��б�>k��]/�jb�db��[J�6�`�=D���3�:�[�
h��Kz��w�y�c�UU����0�!�^}UB)=g+P"UF�a��^����r�#��.N����72C��- �>=z�@�J���u��$��ye�лO�J��/���KH��uY�C:�z��(���3o�<����^v��F���,u��x�	i�8p &�5�G��ۇ*�"�Kf�c����(�;YAN'���*s��"1tL�v���u9�����M�>f��ܵL�*�W�L�b���:2ɔ���B�F�4i}�7\�c,XY�K�}9���B:]�t��{��_�׶BSO��1 �Ԇ���qb�>/A+�g��IV�mV�5�ef�U������U+Cw2S׿V-�m��zQ_v�ك��Vx}�k�nh߾j�Hr7M<����J&ϑ9�s�n��^r�ש�������"B���VMcNgH��Ւ����yU��n��sTt�ϭ$G*������٧�`)Î��z�Y���j��ڷw���n٪�l.=����� �+KWT��{�ԓ�4k��e�����H:�1u"ݮ]�J��}]t3���A�?�l��%ǩlgTڶ�ː@���;�`0���I����K[7o�|�y�w53+���m�Fe
7O�d�$3lU�.�Ռot4�_˫r����$ш�Yb1��4W�Ȕ���ɬ�i�u}TsV��]R�����<�b�0��;v�eJ��(qq�t'�ʒ�k�')=���y?�u*�픡��&ޛD\%t9Ve�U��쨌M�7##����=\��[Uj�_��d`�e|v�ڭgᓀ~dLDFE�q��Nz%�*ڼ-��b��/�$t���g���3�I�!���*s�I[]%�Ƃ��͝��Y��4C��I�oU�	��!+�Ig$�6:�t����W+N=j��IЊ�=�Z��k\�V2TU-Zer�t��*S)&	�nݢ�}�H&j��=���_�HaS��L�*�Y��?x�S�W�8��A�@L:TD������YCg&~U���JJ2��M�����۷O�U�w��`���4�eɼ޲�CU/BӴi]��(�8��;��[��.�?G��X�(U:�N�H���Q��H�������܇�}޷G��YO�����Ǐ�믿T�o��ѽ��z�����d�1�F��(8I	�^4o�L��]KJ����MWz]=��i�suj);�7�����/�yJ�99e�2�:Oα2w�T�JG��&�;F5J�$�v42 R"=��M��R�&��x#�k2��q6e�&5��؏�d����j�k�#�\m�5�m�Q�ƈ�]���:�i{�w��`&��[�M�*>
U��1���Idsr+7,�nS�+�����]M��W���e<���X�����z�Uѩ��jH	���n����dLm�zu�o���.;�Ɂ������O���V��G��*@Ib���C���l5s��J.�J�*��<�f"W]HG���e��@u�*��d�;Y����r{��jh@o�X퓒�F�3^�kv$Y6P��7o�3e5o��u�`>?��>�P`��+\��U���Q�*��SNUC�1G9��qk%�Nӽ�0���pk���a��򎥚�gϞ�V�;���˗/׳N�`��ʒ�F^}�5|��7�бz��޽{��%�KOfo3_IU��`)�hf��0HR��g=9�!c��5>�'
��L���C�v�\�3G�f3u���@T1�Yn���5��^*�K`?�a=fu��eض-�:f��#%g�/%EO��c�6����l��ZĐ�3z��K/����)�N�p"	��(�H�`)�W5�s����OT͝Oǎs��
M�?��$&�?f��:U0��8ӟznC�u:N�n[`��(�mHNކ�9�]�]��7�B<�*=Ʒmݬ���ڷo�zi����A�p~PzȘ*�gdT}�_��Z+�و���Ы��`^+�{'O�0J�\h�8��TT�Mu�H�ʽRU}'�zY����?���_�e��]	؇���%����t򓕮�ԫ[O�Ѷ��(��Ν;u�۪v�59���v��1̍f63�٤������Y����mT�:1������]޵Ls������U���v���_�d�R8�rF[�nÌ߫�J�̭>RS�v*���� Q�������*K:ffe!.6�J����]�N�L*Svq9������m�2��Uږ����۷��~�]���R����ft���;�-^��k���Æ�;vbʔ/зO�c6C��gb����|�z���#q֠Az-i�O�^�zhּ6m�^�e�Mz�}\_s-������6��u2;�$x�����BNN�I�d�����K.�Z�%yd^�#��n�Ն^3'��%k�r�U)}���^��u��]vN9i�Q�b��yr2>��s���d6�����mZ���O�܇gq����1��_,�"��u�֣e��
[�n�ƍ��mXY�֭u��(ڨ�^�nv�*��|#d	S�z������H���.���R� 'AIa�������������t�m6\~�e��/�q�:��ٰ=y^z�%t萄���G�)�L@1y��X��?�7��s���0{;�������`�1�Х��Qe
N+LtE�i�쟱{��>���٫�^~��ߊ �y���T@�a񬁕+WaŊ�8픓z\��������s�~��*cQ6@�&MФqc�h���:�����N~3u�	[yU�5��]�}�Νqɥ�`��qz&'+�&M������ȣ�e�i�l���{((��L&�hּ��'A��9���[q۱}�f�*���]wމvm����ٻ3�NG>���ckšO�����}'R �=$�����s����>uON�2����.\�_���Ԕ�أ�d/:��]�>�p�'�se6s����巽BL��:/l�
�W]}��6�[��e����+HHH��s"�ë얔m�*�?�̳ػ�[�z"��.��{�*w�R��ۯ�;��f����0u�T64`S�����|K/���ŤI��úw>ё����3�w��S8�����^ݗ�^���k ��r�ÙY���U0���;��2�UI=�S]�h�����z�I�YN�l2����~�m�a�S��p���؟��}N_��o����W�|�^�/��,^���dNt��7�|�.e�:ݎ^��?�|UZ����&m�'N���N9�J�/9�e+V���^Cf�� ({+JO�s�=͛5�B
$��ڧo�4�GX�1�=9/�8mޜ����W|e�Q���o�nW;g�uV��i��ЭÏ4�y�d����Ə:sJ"\݀7� ��*O��+/��6]���O�^<p?ڵi��	D ����3Ĩ��x��`����E�.]�>�Yg���y�υU_��[6���c�L%rmZ�:���j߇^��*�[�V�hѪ.��|]�
���O��UW_�y��!+Ӻs܌�CR�x��'sd�Lxz��^�cǎՙ~o��N���5ADd�^��j1���<�Kܒ%�ωe@p�v�����ª���n�{�X6d��a�oa��ŸM��SZ������6�I]6mقw�yWW��L���NJ�W_}���
�۞eY
��oT���*�;�����J4�0t�0�ya:�kW�DN��c�.<��p|�ŗ��l�$,,�^{-�w��`NU��s��_���V�z~~�|��G������n|���ҫ�ɧ��?{�j�v��|��hP�~���ccbi�?��}���3rM����t�SB7ٖQ��XRU7��0l�CؽSz�Z}A}����O=���'�����y��'�u�V��c^r9��,lܸ�~����5V�Ҭ����X�W<s }����}���~��3>��S��e%��_���}��GqҀ�^�&��Zi..Z�J*���7��/�p��	'���E�������{J��}��WGw��.:s�����q�
�����"G%_��Q����g��Y::{�ٺ�����w����<k�̾t�����z�T��n_���N�e�U�Zn	ݕ蒇L6q�嗫l�	��jއ��Ds~�	���;Z�j�~���G�����84i�1��:�K)\������{�`ٲ�X�d�.�oS9��Y�|��LO��1ϣm����}݄x�Y�իWc��%�J䤏��ٳ�f�\}�5�����!)Ig ��N:mڼ	ӿ��>�[6m.�WYN�l��?��^�`NUi����{���#��]z���eMM����q���~-[�@���}f��`��ǧ�->��l\���8ѵ{<��Cz\zM����j�ɢ֭�z���];q�}`��i�ԩ���9����ߥ�q�1��+�ak�r���6`�ZD����_�uz���F`�~�+odC��v�����٧vĨĠN|��)�H@�ǲT@Vw�����}�߳|�I'�ŗơO�^���ӫWO�5��s�^��[-Į�;0�����T/5+��e<�L#����g��)Y�p!�'o��᫆����`��0���@T��b-*(�y�ر};�y�/C@��z���xRe�'O���w��4j�	ut'���=m�r����زe�*I�.��{�F���SO���WMIg�}Ʃz+U��s�^�ru2���4���as��2q�i������G��T@/�#�蚢*\����$��z��c\r�˗-��Jg�[��d!�Çӽl��J���0���{�y1�Yt��9 7�9C�F���裏b��M�ԥ��k�v��~�=�UxD�c����<��Ư��M�5�SÇ��T����hеR*0H&2?� ���C�v�m�#遽i�z���˯��uהφ������3#��y�&x��q�X���d������u2
���X|�\������{�a���HP����z�Q^���ß�Rsx��e�^�6mZc��Q�q��ɖ��\+o�:W�L�ÿ��[q��w�I�FKdH��a�����ß��E���^)z����I���ʕ[�ҵ�J܆�63���&%ntlɽ�X}wF??J��ߞ�6�I/k�Mi�W��*�+�[^F���mݦ-�����
�\�����G��X����f
�))ػo��Ŧj�
��k����={b�ĉ��������H�|=�ze��W��SO;��s7�W���$��;g�^Fv�8���-2����U�9�s��:�	���K����ݺu�Čp�3���^��:�=��Ӻ���W^����aZ� X�E�ʻ���=22��q�}�����DU�]N_�#�=���{?v�H��A����HNN>f+\)���ˣ�����?��ުґCf�[�j5������G���!O�[OO[y�5W��s��OH�۽kL��:��x������,l.�H�M���O���O9�]w�^�F&�����^!N����5Z��W�������@�S�Z4���q��^��z�Ksp�	�>����*�e���G~y]lt4n��z=c�dοV���7��~?3��C���
�Q1�ر��Tw���6jРR���Ɏ�{��^�Z���bu<��qD��Is�|��F��}\(oi���9nӦ��=Opv�A�Н�����Ti����õ�K�L���m.���lݲUw�������HH�G�vmq�	'b��A�ӻ7��M�[�*Ty_҃]ޓ�������3�`�?ر}������К�fG�
�mU�\f�2dN:i �={+}��^�[�e�v:�zᜰ��Wmʾ���t�ֽ�LWr��I�V�!5r���֭[�kWu���Ǒ��S�Jur��=�d�%�v��!`��ʔ��{�,�w9���� ̋.׿Es�믎Ӷm�A�Hy�:��2r�sz����9?��ʕ+�����ɽe\
Oa���Eb�D����w.NS%r����Vi�٣�
n9% ��e��/=���tb릮yZڡ��/Sjk���W�\i^�fK��|���i�Oزy3���c��B��Zj3dTP||�����K����]],�J���մNG�s��gC�t�8�3t�;v"y{�^&TƖ������Y���HH�ڵ�PO���5k�\y�W]�fw���[�9��&w���ur�v�Y�F�N�e��Y%#=]�Ws�$*�j��^f��ر:w�W��#d����׫�	Z2���$�뮻���V"""W��+�I���>����QQQ~�ŕ��qϊ]�#>@���S�/�r�p��}e�#������-7�d��|b��+}lԵ�N����6m�ڵk�z��}�����lnn���bս.�=˒��ڵC'��v�{�Z�Z�
��s;��S��w�-kO�\�����S�|��/-�%� _��C�:�����Sqݮ

�����~%'�:u�ѨQC4i�T��1�2�S�
Ԭr�"�W݌�*ˣg����ِ\���5���@$��A)J%J2�Qj�����_��%�o��>�]� C��2w�zߒ ��� ��Ë����}�u�Dӓp�:�ʪ���qU{�o�VD�=��������"�LU}��qq�Q��)�/�I���&=ⳳ���ס�}��$�(:yHf˰�O�H/����r�;P�7��aUu<O�Tc��Q�9��k������΀^)f�K)C�\����b?�w,��#��L�im/��;�hݥ��8��|��8ގ)�ňp�z�����<��58��0K���0�~L��6�@;�\{u�yy�PM����Ni��f7����YB'""
f�S\�[y:�Q�ѝ8�)������^����3�-ӯ6�|v�#""
b���������(�ٝN��ֈ���7=S\�[�,HN�Љ������W~	]�9:����T:v���3M�r'"":�����,�Tn�7+�O"""
�K�ݯ8-%tFt""��d��m�::QPR1����DDDAKW��UBg�8""��e��˝Et""��U�:#:QP���U��8t""�`&U�~lU�?"""
F��ΈNDD�̊��3�)݆ι܉���;��~e/w""�����,�NDD�L��YB'""
jXm�m�DDD��"���������r�z�DDD՞S�r�5""����U*�}�k�r'""
ZR���VN�f,'""
fz�5?7eX'""
V�ߋ�0�'��,�U{�˧2�5?�r�܉�����m�r'""
b��U��DDDA��Nq�����(��~W�Q�b�;Q�Ǚ∈�B g�#""
~�C�˧2�+��^��DDDA���2DDD�ʏ�\�L��NDD���ΨNDD�����*w""���*w""�`�ʝ��(p�8""����kb=S+'�܉��B ;�U\m������K�p.w""�����\�DDD���X�U�DDDA��Q��LqDDD!����,DDD�*�˝m�DDDA�ɉe�������CgX'""
R�
T�Q�͉e���B��m�&�܉������6t"""
F�U��Gk��DDD����܉����
t�#""�`���WЉ����Dh�m��(񃈈���aT$��UBw8�HKK�!�p���� �`PS
Q���c�=�l����j���둓��ז�n��0l�C��Wæ�5�������]8
�������p����*�&6���e��-�8\yS~U��^�t1����h2�g�.��6��sDDDt�I��f4��&��� ""��JJ�:�烈���+UB7��͖n:�� ""��Hfsأ��ege�U;6�-3:::�^�n��������{�g��0=""�I&������K���;w$�Өqӻ<�t^^^/�4cTD��u�ƪ�3*8���c:1ϑ��g�#|���g��OF��x���$�����jժ�y�����W�<l��k�ŧ�O����;v����LP�F��]mn�G���E��l6�&m�v��0�æ�`ap�4�����rd��ϫXf��Ta���
�+����ſ�F�_JoWl����l�	�Q�k1׉x����󇢿B�8*�g�J����b{/���}����(:f��Qxn(���.u��{�`[�~���0T�.b�ҥ�{v�
/���G���NC�&M�T�^n7TWr�֬Y����[f�������=��ILl�o�Nɟ�f��MX�<[Q��}y�~����1�\4%�Y�wϮ�����,�{������vW��3K���yxv�c?%�l�Kb�R��\��W���)|q9��,q%��[����ĮK��}���n�a���{��_�]�r)�'�z_/)���N�l�b+��(�-6-�Y�b����J�-��ڨ�9��G�}{ΧԖ����t��pJ�e���%���-:�b�G�J�JM����.rџ�ݠ��:IϹ��\�������0̘�hg|BvIIs�����Saw���ʇ���G4�΅�Ϡ ?W?j"�gY"P������Ӑ@�p��ÐB�l�S�t8W pr�����T$u:�Õ��p?����w���&���\]$�b��$�o�^ܙ���kѾ����m6�����u�]o�ٽ�ً\t�Ÿ��[Bnn�;z��͸�λt"Q���N���on���'�<�������OOL�<O�EyUw�g��&�%�f�L������õ�Y�I�?\���u����hY<u���	S�,�;u):/��s�]6
ӛb�r�����
_��G���R�����̰�^����kc��4�ͦs�6Wy��-5�0�\�����6�]^cs[�e�._�CA��o��0RB�zHٿo��>�S?�� O�l٪UH��7�

���Vtx�is8t��4��J4�m�j��m�w��/�(5�_�O!_ega2�J%J��#��X�]<�g�إ{�i�'6�^�٧�Lexb�Y��Z�;�'���|��������Jl��2y�.�-�܌Ȉ��Zu#WD ��x���\���j�ژ��~̯s~Y߿}���E���[_a��p�2�mW|�ҥ�R��(�P�F�s+��(��/��(]�*��2�M��x�k�9��?ós�t�<�t�B�{��#�?=�Og^�{Tx6�k��F��'�����ܙ��r����w��=��M\�C���x�y0e[��|�}������vU��2��pU"R��Ɂ�
��c8�Զ��r���گ�S������r�Jt�ܹ�ug����e�,���o��� ����W;����"�#

�eF���e���سgZ6o�/S�T婌���o�c��-]:�mҬ�ks�u���'`��u���+AD,Щ���T<�$$$����J��ʬWr[�l���kt@�`.�;���*CS���f�^��?�>��t��6��{�Q0a@�2ڷh�ǞxR�����v��V&����a�?�`��A�>������_<��sػG��R���Jn߱ø���vh�] "
F�d�q�&�ݧw�_|�^�ڵ����������:��m;����x�駱j�
������f͚���/s�~y��6�w�� "
6�d)-��p|n���V���]*�J[�j5�nۊݺ�:ҝ���1f��y�l�i80ԫW��O>��/��Lꐄ�cǂ�(1���N�#:&f�
�y*�G��¦;�-Y��������λ����(�	N����h׾ݘO?�$%'�0���:Y�6�6m�ʔ���#���5*�M^n6����\s"��Q����{���K���@��0�=�Q��o��}�'�?�fM��;�"�`ŀN�.��b\{��6�#""|Wf��Ȫ/���K����^�jӎ.�bي�1b$��މ��\�����g��w�;��>�Y'>�G<"�`ƀN^����۴9�����U��Uv[�n����t@�$������ѣ�d�b�	�JtTTr��-�L�655/;DD�:y����`r�ڴi�Ff�*;ͫ��b�e8���Q���㭉1��o`5���W��k�.���� �n��O?"�`ǀN^}�~.����j���s�yyQ��q8�p�"���"*22��g��oLx��ٰ*�׊��ѭG��Np�����޻o���:`@'��M�ݺ�@TT�&e~^nS�v�U+Wb_J
Z4k�`�i75r����`��y���ϛ�����C��޻Љ��`@'��z�\vŕ��Ď�QQ۳27-���m۶bÆ�A�u��~w��b�vs�ݞݰA��+W,[8��G�Գ;n��jU��S߾}p�ק�<{�Z〭�%�:tK�.����`$����˒�����|�)�ߓ���mxi� "�N�ɧ����
���e�Ͷ��뻗�t`ѢE��ɑ�AՎ.'+��'�h7���]ٮ}����-c��� "���ɧ_�͚�D�:�W���g��^�j;iG߻oZ�h�`�״����p���n7���hܴ�����)_}��K�aԨ "�n�ɧ��.B�=l˚ի����Xt��۱~���	��SRS1z��^Ǜ6�,����\�պ�k0�|���K "��Щ\	uиq�ݪ�%=-�M�-����y��y�5�fϓv�I����v��:uz��/�ʱ���)�����b@�ru��I��9�U�a�Q�c�t`������Flt�1oG�v�7&L���[��#���7o�r�/?��y���ؽsN?�tUW�T.w�8�{�^�򚣠� �j�U+Wa�޽hӪ��x�#Gc��vsy6���s�͜�����O��3O���:c@�r͚5]��@|B����������e���ؾ�֭?f��<�`�E���_{�����/���w'OQuǀN�:��q�7�t:��/]�+++�n٭����v��:��(���y�EtL̎�mڌ�����0 ��Qv;"����_�z����/��?x�`�mLӡ�S���BlL�QoG�����7����`n���7i������3#����`ND!���Ҹi�rӍ��:���l��]y�e���ػwڴnu��MB�Ju\�j߻w,�����P��'�<��AC�1۶m��oL Q�`@'�<��Ø��iG_�J�9y+�Ihݹs'�o�p��������`���n��]�v�g�������q��_3�QHa@'�HǸ�I���Y����J,�v�e˖��AgU�9I0�/(��＋iS�I�?����#�7i����[2���ѳ[Q#��ÀN~��q=��t"۵�߅�2�3,�V3��ѳ��sƣ�4�g���k��΄U����s/�`J��]�v�Z<x߽ "
5���m����n94��S��`5��X�z��KA�U3�g��u6�y�w��˪vUX��]��Ν;��釙Y���� "
E����Cҹ�ٳW��av�� ?�2��x�M7VY@��JO�ر�������n�ڢeˑsf��)�a��_����Q(b@'�=8t(>��+ԩS{UDDxFA~^�	f��Ұt�2�y��*9��~�?|���0M'���e6���Mz��W�r�x���0⹧AD���o���Z�i���M��ѻ�23�Xm�׽*�G����ܹxy����̀uU���s���Mxz�3�5�[��ND!���ֿ�?^Ƥ����/������m�5�Wc_J
Z6o��K0߲u+F��m[7���m�ڷ����{�r���_���?Q(c@�
9����1))�s�n+m6���Hޖ�M�6,�K0����K/��彩�-�����4m�t��?��9���дi\q� "
u�T!��ɨ];			K#""rsrr"�n�jG_�l�vj@��0M|��g���>���U��a��~�ĩ���K/3���1�Y��Q���N2��3q�"22r}dT�����&V������%K�������J������k>^�"2��[���ۻ��*�<��?�����n4$kBGMk׭�bv�r�s'k7��f�v�Y�j^Rlk�Uh3#l[��dE!0�&"��*'8��e7��s�[�<|?3g8����w��9���L����ܶ�3� ���~�>*J���k������%��8m�F�Y�Dz򃴘מ���5k��\���G�|}[Ǎ�� ���T�|~�3y��' ���~�6�f��ҥm�3�t��_`�Kjj���ٳ
����Z:;e}F��������zWxDĎ�~����
� ?_�n� �pB��oK�zJ[`ƞp�m%��e����A�%-�-RRR"���;�jQ��y_v��]v�����	:���cGW@@���1��v:��Ç%.>ABCCK||}�m6k�����V)*:!]6�x�}:��W���Xa��MY+��f�����	�����Z�N��M*{��:�m������gŠ7T;v��J{{���_�|%M�&�w����74HRR��*+�^Q���ᆌ=|��W^����አc@�B�d��Sr?ʭ���0�Ӹ��*����	z_h1���ƍ�$���<��
�?w�?����/�k� W29�$��ϲ.%��*�~���p3J�su^ZZ*�Ϝ��s�ݷW�l�"6�U<͛�Un���o�ަ��RXX(��� �pE�1 ?��DG��M�'����X-���q6[�?^$֧�b4��禥�Dq�$'�H���t�����=>�Ճ���; �.\���x�ጠc@���f�~��������k�X:�=]Mk����-�q];��,)�k�d�	����N'QQQ{�WO�?c��v����+ �;��������L1u�
�k/{�$?w��������&[�n�?�#�}��Z!�!E3�e���hjn�m��  A� ����c�>bޙ�uZ���{ڨ���(��e2c�t���ҝ��'37HW�7ڢ�r�K�Z~:yrʮ���t�3R[^..  A� DDE�,0��_�Sl��~�����(/���EEb�Q����{W���%yM����Iϭv7��Fo׍��;�צ~x�;��Ȋ�� �_6w�,���Hxxx�ȑ#-�W�~�o�����XZ��亠����F6��Jj�:���/�Ӽ���ZdT�;�ߙ�>����%9�� �w:L�"uz\����-��dn�����R[S��o����)ٻ����i��%A����3��^{�g5���*� �C�1`�G����>Ѿ^��Ω����t��_� {��S�Iz}O���]��.�X����s����s�bc7�d��ߕ�P�1���y� ��:eF|��
h	)3��6���8m]��۷K��Y2g�,�8wN��$u_�WK/��i���_�Т7W�|�.�,~H  �"���ks��y��t����ߔNj��%=-]���$c}�=rD<=��]�GFF��=gv�ƍ�N����
 �cP^߲E��#gΜ)�;엺�����򤪲J*����Ԗ�u?o8j��֙�fnX���g�!�>yR  �t��%�n�Nʻ�|\z��t~�)�'��MR�e���i�L�]���훶lq���ɯ�<)  �:�d2ɒ����������ں��tz�~���w'L�X}Ͻ��ݺu���ݻD�d;A��tZ��J�:m��/>q����ā��%�GZܽ s�����j��u�̝@t�'��˧G���;�x�iʦ���X�V����`0J\|\ުU�v,8䊈���� �aC��?��{\Ǝ���?���b}�.�K��`4��W�Ǜ��j����pF�1$��^��:f츎�G������q���>��K:�n[xT��i�ؤ���[� �Cf�Ν��ޮm�r�������T����C�i�+��<�����-�  ����2˖,��/���s�J�ط���w���-���*<!!��]wߕ|������� }G�1���ِ������l�X��m�I=��������3>m�^9��ŕ���*/���  ���cH͙3Gv��-oeeɁ��"_�$�ݑ�]�Qn���z�;f�y��g�9��ӈ9 Aǐ[�x��d2���D����t:&8�UN���|�����`4�1��Eǋ���ʤ��V  C��8UZ*:�QBCB�'LL375�X::��lA:�����'wtp��u��wZ,�z�j1M�$ ��!���86ih��^��������dn�:V: `�:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
�O��Ր���    IEND�B`�PK
     �)K[��EM  M  /   images/d3694a2e-5bba-40c3-8069-8db85c4c9209.png�PNG

   IHDR   d   d   p�T  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  cIDATx��]	xLW~��d�(%�J"��}�%(�Z���B��_[y~R�R[u�E[[����J����ҿZ��j��B)��'s��;��Ĉ����>���=��s�s��-�37:�PTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��AW÷&��z\I���7�)I*�Ev�Z�:d;iJ�3mtRɲ�������V�$IY6��"a[�d��$}/����~�l���99��t.��$u0Z��d�M��(��5D��a�}0�*�
��?���h��dY~�`ȫq+��L��yY���@���[���������ƍ����0��`�Aк�C��"�|<B&�������r����t�PQ:�;w'N�{˧����a)y���3�t>���ʂ
E@fB\yyP� �f�3b�1�(p�3!�<ÃY=��䫄(�d���?0��&1A3vH�JIi�	�YCd��c,�p?��0���g�Ж���lqtws���%b�G��ɒ�2d'jaxR�v�Zl߈s��S�����_C���2Js;�i���8�f�ɒM>�Q.]�����С�x�g/�5J<����зO̚=�g����f6.:6lX�t]������B��5�D��;ѽ[7���s�p�0g�,�n�=_x��(���E��~/���u{���F�m�6�2�h��!����v����;����dX�i5�7�}�����ٿ�2~޳?��#n������1p�@xV�$��u˖�Ѳe��H�zi��|��u��,�Ν'�����ԩ3�/�5PP��7o���,�_���C�޽ѵK���ǚ5k�t�:>�,^|q 4�XȺ����7!&&�+{�_�~��d��ǎ	SԥkW�o؀������A��n��B�p2�7n����Na��>$3��ARLN�G��&����~�� �����QQ��wq�������Тe+xU�ºu_ lQ������͐�լ�K�.����ԙK�.��9����(�QN4|���X�p&M|�����5�OLLDu��x�"�.Y�9o��&�l7ww7�b�rD�c�)��?��޽E��jO����[���a�0�?B��ۿr6n����o�Y�}��E�E�:uh@lAZZ*�i`5]�ر�u�9Ǻ��<s�4�V���ի۽��1�Q�n�:AƢ����D�?O�F�g:b����a� i4puuÑ�#������W��u� ̜�iL8^<H�Ȏ��ʕ+Bui������®�v�u�zS����u>l�ФΝ�P�U�@.��+��������^M�5c�L�L��S��nW",�Y��e��'""#�|���'B�B�FMТœ8���	�R��ӓC��w��t�b�_G�R׿ƛG߭~=L�6U��?���קў��ݻ[��Z���\�rLd0�q�	��o@Ey.D<kI��
2^U��~�zB�!C^65V�E�6m�W���$!-^�j� ��溃��������͂�٤������m׮j׮����{��l"��e����G�fg�AQ�%{ΫbM�6��F�흚6m"�.\@�ƍD���]P��	��g�ΕG���e?h�V��\��ӊ�����ٳq"m���`1i.�[8c:fd��Y����<P��6���׻�2�sq�{dDG2kd'j	h�͛��)2;U�jW��%�=z|j���)�b~b����!JcӁ�L��+$3�i��ߪ[�Fc�8����2�F����~~���dG��?��%\�9���ɡ���3lw[wGDD���Ç�6�V�Z8AQ?��6U_"���YԢq�0��$��_M�i������W[P��@�nns+�F*Z��@'����!����ǤI��`�<a�CI�>��p������<*T�[�Cɩ�1K�,>�>}�/�h�M�vhD�*��89�-�aq�֭�M0m�t�jQt������5k?C��M�ۻ�Mk5���Z�e����ZSVY'�����L���������'����F����g(4�Ŷ��P�^G�>|<(��p������_�R�VUDK</`9rr��WhI�6��E^��9��~��΁�ʧ(��K�c��K�^���}Ѭis<���b�s���J�efp �e
���,���5��<�5o۶oD��h���%.�sab��F��%a�ȑ4I܍��u�Ȗ-�!00�==̤?�9@���������A��"���K�T����J��2
�������r�̋h���C�Шn+���\�t	�i~`�'t�dA�����Ӄ|�'���GEDCQ��z�5{zP�gA`�@��?�h����\�h*��5���]�r^^^pbb(��1��[ޒbo�ػ^8�s4�叽|�4�@����4}�#0(h�my
?A�#����Mg�<��7��?�il���_ �2Eto�����"����j�37-N^��4g��)�8����&��'�*JBCLQ�JH�C���=d��,���}X5D�2`�����0��g窆(&Q#,���!�.o���e�TF��[���9ʲIQ�[�<l�M�V��|/="D�xOR���vG�_G�3˚��7��aj�gE��s�6��ˋk�Q'I����܊�GBEiB���j���QCG�h4Z�D�$ݢY�-R��By%�V+i�T���I|3����4����ĉؙ}���2r����)���Om�fk\]�zH�|�R�iO�l�Mۗ�I6_dْϜf4G��Fk-匷�ݥe�k�\𛍶���V���_�3���X:�-�b(ڴ#ݾ���KĤ����h$�v!VI~}��+s�^����xg��p�h4"�E@�Ӈ$^N������1���	�����ǁ=j��������o��qbZW�?��i�1��wI�t�G��v��e��^3�x޹���k+�t�w��`-;q<3��rJ�r�##���Κr$55G��޶;�a�±c_�ٿΜ�V�{J9�Ԕd��=�(B���}�\�.1�7����׭w�^v�.\�[��"{x<����̣������{�"o���]�|ҵ�"#��[v��n�ٻoޚ>�Mۢ�̛;[�A���(Ks�#�����@�V�s��I������׸��������gn�fV��8\��@�*e	%F��#�n�����8v� �2�Ǎƙ3�2+yV{<6���ܜ����#d9�¡��ȏ ""�z�ז-_�M���^nzjJ�QNk��i�܇��#��~_�Z(_��?���&��2�G9��ɡ�=�gge|�yx�fY$�Q�/R~�'������ll���<����� ~�N�z�����t
s�PVQ��<^�q�s��mOrrJ@�=�t-���K		粲24x6�;�;�%JHJJ
*�|D��-KKMN!p5�olI�x��ݺ�Ge�F��kǏ�H�"A�ռ!i\�xzz�/_�<�R�u�7�u�����U�F��K0��N�rx����̬L�(B���^b���x:y9��}���E������k��%u����QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB����Blg���    IEND�B`�PK
     �)K[	��} } /   images/bbfae99c-8036-4c5e-89fd-a87441410720.png�PNG

   IHDR  �  �   ��ߊ   gAMA  ���a    cHRM  z&  ��  �   ��  u0  �`  :�  p��Q<   bKGD      �C�   	pHYs     ��   tIME�#Պ�  � IDATx���{�m[���Ƙs����8��GսU���袍�i�4��A�("�q�6'9�Dq��E�HEVd��HX�d���&�Н��g=��n�}����ךs��?Ɯs����{����f�J������k�5�x��p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8��}�𵂪 ʳwQʄRZ����k��{�Lǁ�%O�h	*T�J�`011@��#�QD
*B)�@ FI�"4"L�Db4��L[�>T	
4AU0����11��*��J���N�L� ��m��l@�(`\m.@aW��7W�G�|������%���<�Ç?���p8��h��@K�J���s�H��K���EFi��_j��R�kh�,A	P@	`   �jQb���!f(PA�U{�B8��W? � �FE}E��z�T�0b��P�t�>��1�yPr�P)[��7���I�����>P�+��T�hT ��ۻL���J��ui� ��5%Nd?#��z�vH
U�w�[��}��rV)R�""�%' ��f�v�U!�bs�!lJ���x�/.��Σ�~�S�����G����7 xD������%b~�]  A�=��~l�,!	"bz���
�*�E �
$S�
t�Nb�Z�L�WaEM����DՀ�Ĭ
�h�AU���!7�(���?��˯���1(��a��%�۽�����]���$���}i8���U�5�ժ��T�[T�GE�C-�J��eC�����	d�VE�RM��F���dQ�liO~M�?'0�w^d^�b�Op�x<��L�$����3x� T"��q���/@%B���w���w��ڄ����k��3o������k�q����:Eӯӳ� e�n|�Z��	U�M"�7h�Yr��((W���� D��@U�����y��䟽��� �6� ���X��D%"H�T�(�R��0+���	|KLO�x��8L����m.��>��m.@aa�]�%����P��/  �Sm/�J��eM�7h.�SD��J�$_+t�RM��
 ن^X�f��@�aJ��QS�t��k��纽o>c8y�l�BqĻx<������{MH��sF����J�v�������U�v�+��K�������]^\��^��������ԟ��|�^�/�-�p����; t�0�>]=����_.���FD�[%���P�)	R
b�K)PUÀq� ̦���2���_�+t�;������2{��W�~N�D�DF���k��q( �fB8�g���90��2�d�����q��o}a�X	�@�>�G�ᗍ�VU����n�./��'�����/%�n���Z�K*%��Pɦ�T d�ά��H��Du�Z�9��yeӕ�����}N�]�v�W-�~��;?��c|���	s)(���QJA�fB�C`036�`6q��F��,��j�@�.�q�}�_o��v�y�~���g��W~Ƌ��Ǉ��q�`ڿ�_�o~��-������<�Β�o�o��V�|����D2��\!���!F\]_#�(Q�W�Y7ƽ˧3]oqǕ�\`S���"ZM"�� J�jTM1+���y����M`��P���ϙ�gƟ��~�Ke�q�1^\!��1��,���;�������/b�]�����U��HI�Z2 ��"	���`^yۨ�j���l&��mH:��@��l�
^P]���u�{	@��9��s��{<��s�7��.���L@��i��%c��؍6���1b�<b�#��E�0�+l����U�_�������b|�_n���7^^���, "���~����g~�G_�2��W����O�����%�v��7�i��|8n��[���R@*��PJC��`�!9���E��^z�U쮯�(��RU����� p� )�z�5���5ki_2����&�5���5�Ye.1WEO�����9
�'����e~������3������1ݾ��}�������o����!����?��9�.��T��9���I�"')�
�慢�B{�g�Z{�^IU��mt�Y�8��ieٮ����$��qԮ�0Q���.~a�9|*���ÌL���9�((#cF�P��BDĆFly����.�<`Ѐ�p��Kx��|}��[����/�~���T�O@)������W�������~�ǿ��y��/a�yʘ��b�]���o�Ͼ��2r�~��p��3,����4�P) ./v�$ bLsƓ�^z��x�ʫ��
� "���ӅA<�t����<���])U��kH��Wy��P��]��� �r��G��C�U�/J?�!�(��#���,o�M���#���#��p}�����u�П���|�G�|���������e��_�|+��*�Z��BHU��(t�ͧg}	yK���*3
�U](y%@hM߯��@���a�y��`��s����N_�8�@IAA���`F �!�b�
��1�6<"P t�J@���p�勏��W�`xTv���8?I<��ƿ�H���4��.��C   �7��+��4�i�p�x�xx<D
�:�ߖ�߭i��A��8o���� � �3��Md�H���#��9g�./����g�N	�^~��������Č@=Q�z�I��;:_���LV6�^�l��H���_׾6	�<vQ q�P��@���Y���q�� �o�D7x�c����@�P���/�*��A_�����폐����_�^�����Ayz�� � �J�h�V���c��S�w�Vν~I5!�)t�j�/%]š� 뤸��P���x=@B"��%Ct��@Q2��j�H1�Z��JI#2fd8!% `@�� 	!d��������F��:��?����R/�t�{C�o���6=~��v��o�~�qw����AU�RP��Bd�p�:s)�ó�?V4��9�ߍi���p��·m)�I��{H:@JB �%�'H�(iF>�Q�H4(�>�@cA�	�M7�i��;()D �%oz����q�9t�:W�dg�o�;��#����u��I�%�X�a���|����(�߮y�#!���@o}���8~vs���[_�N
��~$�}�y��޲,� �Q*��9�%��kXӀ2A҄��4�z�P���oYY����aJ�E�*��j_�*�cYXk�PN��l-(/4;��.�S*7����S�����	��IZ
� H�H�.� K-��"
5�d0�6؅+\�x�W.���xix	�0"`Ѡa��4���g���e��2���x��p����-!����n��K�u����9��3 �����͗���o�*2��O�\~_��o���O�i��N��y"�3Ho�Z 2!�#JN`"��9!��r�0�nn )!��8D��r��E@q���5~�۰���FFV3#R0Yc���Q�.DW��ޛĉ�~��P3	j��6��*s{ͪ���O�u�y�T�����UM�0(�X
�'a:��C�i�ݏ�{|����Ȓp������/	_W��/}�!l>���(�Z��-��D'@Dg�(D$��I�\��%�-h�Ӿ_|�U�v7Zy��1o��B������״}��;��"�ܴMȋ�iT�b B$�j�,�JBT�[J�A�X���B� �غ �H ��`@)B�6(��3o��4��4 �	�kL�c�O��g���8�0��s�Ͱ�~i������w1lw��t-����@��m�$�9���M<|囯5��۫W?6�~�j���K���U��n�O!�-�dYfhI�r��-E��	I,^.9!oq�y
��0n�u����3�4�c��ͣ�-bܘ�#��a�K�J��J�S���$�U�ng9��޳�R_T�9�h�EƂ�@�����OՒ�J�I9D����)㯕0��D�ߺ�<�����~������������O|�ʬ����O�ւ�Z��!�㿡e�(�)G�r�j2[���T�<s��qن�R�T;�Ψ*t���F��9��z�Z&'銢jT�4*���-���9��ւ�Y�]D@PD
�H%�&����Q�VC��H*�b�#Ka�]"�Lϰ��pF��~ʀ(
�y�&��M��7s���Y���t��1�� ~!����g_�t�3�C ¸�Ї��43�3���/�ٳ=��
WWeh���u0����#��̀�rP@b-}�j%A���BH�L@mX����D���Iָ���Z�X�K���jZ����1�}��p�b��`@IJ�A��AT0� Ί�2f�vD���q����Q��0E�t�c���
����v���}����;�y�%��j`���A����o��I_�"��>z=ݾ��*�E�'E��Z�5D8���h�C��	�@��|DIGS� H.ȹ@0�	ДQ�#�t � C���05���uw��"_? �&[T$K||�7�ӄ@������u�{��KoΏ9\����%/D��=����f_tN��;EJ�֛R7J_#�@uF)�e��{�O�����~����~�w~�w�����V���u��o��|���W�|��K�H���"G�L�2�lJ�%ͫn��1F��Ϊ
��w�yL��M����E)��z�ž6^O�:��׾�aU �Z"@�lB��;��,O�@����z!�$(J��ށ ���l���p0R�Ť���3bQ\L��-�����A� ��RB�v������5���������3S��8��"z�oso!�o�?�O?���q(1��%��f�tv"�w��T�Բk�a � J�s�a�q���	L#�iF�G�M3�:Z2r���<�������}��ʟ���G�q���D��2LE��FG�b�c`��B���L��	, )�M��`bb��Y��I ��H�tr��7�>½�
�����_R�U�Fji����P��
U"����V!�K��R]
E� n�b#��:�Ah�t�����p!P �����^������ 8>y��h
n�S� xh+�Q
�60C�~a�.�J�s�JB��g�o��}�f�g��]4b��� )�����/�9^
�Hy@�!��H�q���7��oW�߂r|]U^*%_�f�P�W�Vb�%��@�y�e>"�(ǣy���-e���'@b��%c:� D�4�e����!�@nn��gL9B9X)Z) ��oN��%�T��G�ÛR&��!��Xe�$��nғ�A+��.R�m�e���Ξ-�K��%�i3 c)lT�D@��H��)�''�o.����nz���O��#���a_+|���f-�a�0o����5_)�R�Ũ'�H-+SA˃T]�oQ�a���g�8M�X�jU�X�6ֹ-���s��2�kѩ
Z)�wR��G�؅["D�Ь(�0A� 6A�(g(B��g��#B�dU*`Q����)^C�
�hA��43��A�!��A�^�^"���{�BxF����D�%����ox� �q����ՌF��� r�0��N����N3�W��z���y `_��"����.
D>����d�"ø9��IidC�qP�AJ� �1�C��n�	1��R؍X�S�4A ��(TsE��*7�\5s���C��L꒮oZP�7�7T�/IAbJ]�i*UΩ�Y�(DETUE��Q��q��THJ	�E��,Y@9�EU���PJ�&*��"���T�\��-�˂�-Ƃq,�~�_�9�B�R����٫Z��*���l��r�^�3=��C�<�������`�hH�޽P�E�#��HyՇy��\i�;���9�ΐ־Y�'ת
J� �(%[-�<��#��M	�fS�R ()4%d�ӌ4O��0#猔R�P#�b�R��0����f�� sg8툩9�M�5[���Kύ& ���K�{}��$ԭ����ԍ�ƪ��ηváv�_=]��p�b� �d�I�oU%��w�VDE�n��2��ܼ�i\����zV��*�ӻ�'{�q�M���/i�sH�G(gh��V�V2���>���@��L�QSƴl�N�t^~��۷}JQ{]/1��Q�&�v���^N� ���M^[�f��FR�`l8��#v�E�2CHl�Q��I�d���I�zp�`��DDe	 &&��Tn��u�b@s���\KE2�L��  03�Ja$#��� V�P�C��8&���(4�(QS&��L���U���(I��+���� ����k����v
�<;��T�i�����a���2���(��r�BsR��H�L��HDL̡*_��i`Bd!��͆i�/]1^}i
�U�K��q�u�V�����û��|Խ�6L+MD$���Ｔ}L_՚����R/n�7o+%Y6qVe) e0���([�DDC9BDTPP�([P�P	[`���P���VG��"�%�HI��R��Ǵ���V�!T�T�c֜7�������Z�̌�{5Z�v<UHUI�����V��b��*K� RX�0����b^}�P�*��g��S�Ħ�i�q	e>�oQ��d�Ϥ-�Rl��������
���cJ8���%��ْ�b b4�:M{H� �S�-iM�@cS���YS���3=]<4e�L��&��7��D]Q�2<f-��w�n.�~��G5�,"�mb%S� ����Cx5���k���n��4r�x��O��Z����~��C\~��雟�m�������'PI֛Xg@��=��F"�j��V��w~" O��~M��S4����z�}�,���歯�f͆��ڇ�d��fc5/{TƆ��BϬPeX�2��Q�D��p���� +#h@�!����!?E. �ƂѕD���huRTC��� �"�z��`G�� ��o�����Z�&�Qz�w��y��CUf�<eL���O�xrTd,�X2B����$b�:
�xf�<�3{�D*}K1�ĀAB���0!h��̀a�������D!�����жt����M޻��o�[}����F�,��'����ͻć��ď*A���Rt�-^V��$��%b�p��[HA<a�`� ���tܢ�K��щ�P��-!l*1AF��lbM����l�=Y���
{?�x�=Y��k�
h1o��Ĭυ4�C(�"E���T{OT�ԩf])tj��u{#I���|����) �֬�~��j��|D"R��<�8���8D���M�l"B$��ʼ� ��7S�(�i>�϶լ^�n�ﲹ�l]���{��*���F��* �:�et�볰<+2O�b芚���ĕ(�Q	Py���P��}������ȳ�O��)<x�[�aǇV��~����@���4���n��*�
��5Ͻy�B���4��*���{����z73׍ghq������K������������E1[���
2�P��  ���
��b,�F:� E�Rz�A+0p(��\`��y
(]Yk5����C#��jV��!�׃V�q���#�g*w�ξ(�/pW�j���1�$I @�3n�7�`�@����D�;WDP�@T0�	%[�b)&l+8�b76RT�	��U�h�\�	~'��}����N�25�6��~��	Z�"�	"]��l�
�{��)T��!@��t��i��#Xf��`�
@cy��4@C��-hs�v�n�p�{_�U=4�¼(��8�2�M�[S�XN?�m�(s�5	x.�5>�3��j�I�z�K���O�,=f�{���'��=@5�\�]q�P�#����JNV]R�0��V�V�3BP�t�����^_B&3��R�t ������ߢ��h��t%��2�O����T��^/�k �Tma��0�����?{�J�KM�CϷ��r�若�E�� ������������'���{�	�|�Sx��oy�g���R��޾�gሇ�UM���K:��G�̖"�f�Ve^�~	��!7�l�n[��%�ӂ�-J����ן�)z�+��O7�J�wLZ{Rj���5�X���ʜ �2�H
��N
S�\@�M�Aњ�7Ȥ"(�}ge5�t�@��r�1�A��`�8T��湒V:��}�*�%j�ΐ�E���m�"H���:��`�ύjڽ���D[̀�� �#O�,RD�l1gV�@��5r.�sF))���!R�e�0�-."a`���UjhדX�3���=(*x>V���-LY��u�� ��=�u4� pT&�NвM7
SX��0���vL3(O�<�'j���J�TD  <��:o �%�`�ov ���^rZ�U��Ր�5-mMZ�ЪL�p��Mq��g�n��[Bz��֥��m�h͏��_H}F�Xy�-��׽�O�}��)��a��$	��L77fP��
�����mă�s��2w�v�n��Q&���	6�U�!��o�N�Jj�u5��]�r���5[��ht�ʘj\���AlD���^�Q�2�~�*��~`�L3�j�Q���`���69W`{��$
�����O�G�+����`��e|X�S�
���ޔ|�'$�T�<hIF�kF��PG��r�V�V�̓v.+ֶ�Im���'V���wS�k�ܳ[�u�z�<��/[�]ey�)��ԪI�l���w&�v�@m��d0g(�*��%����6�%P�Q����4`�r�$3����л���ٵ��^&*�W�*ШUi��P�,lM�����Oj��w��(W�kJc�͆ ���Cf�"(U�81B��� �\��{�V0P�Zl��-×a��|Ļ���u��
H��O��T�C��]�rQ�͋�=����v��(��b�.�`���.��9�ƺrD��L��Ϫ	(
� �	�� %�����T "0,��T�2�)��!� V�._�� ���M�	b��GX6�+��:ٻ��5m�*��Z7�6���S�|��β(������h�Z={ċqQ=z�RKK�2��,Dl}�I��,N���9�!0(0r��b��#f�-V"I���`I��7�f���ۍ�<�?`:$�3dN����z��
�:٫��{�����5��x�M�wơ1w"+�[��`�G�����\�3���}4̌��OU�#֌�z�a	J�������9=���G���'�����q��gq�!m@�S�7��T���%����%�XӒ�e��l-=�]����+���f�����j��$��Ic�٬R:�컀&+D�F�¼��,����*�C5Fd@i�DA����2�b�'�f5+�Փ-( R$�FիoP��(2�5��Q��/#c/��2n�G�A���vo����Rf�;2\@� ���l�r�@�Ӣś����O�\ʲ2wj���k=1�B�l@R0b�u��	9<�f(P�le�2Z�p$F(&���d����Lur�Ֆ�R��
�12�����x0(X'�&�-���.���[����J	P�o�Jm�tU�띪�ꋵQz��-g�R�N_Dd���	:�V#���Wg��
��`L�,IrU�TD���*
���n!�-�b��PF 5�����B���O#�-�e	^�@lFT���<'�6N�5׵Z�ֈ��贌����3�L�Z�ZmHͣ�&�+����o�
o��vT((�e!OG�)a�8B�`�7�W�����O�<��֔��|�s�LG��"6q�V�K����YyY�nJ����^��:��*p���T���85�~�4�3�<�ET_������J *5�*˥�v3���k�$9�/!��O����ç�K/�>T
}z�H��'�|�Ki>|���:!�)	��lJڒF�4�Tzh���Bk1�"[�R��tE�uO��V+�����oS�M6,}�[}d}��x��
��!PH=�k%�����(��`�)�X��>6�	!��MHP��D	3� �z�,G� ݮ����,c�f-�|q�5�u*���m�cB��5���+/H� �������Ѽ��x-$R�9�T���9�Br�� 8��ԗ	`A���
)3�
���2z��@�R���RlT-�R0� S��`?r��y�]>�k���ݵߴ=q�e6�Z���<�~��{j��mˡV���Ȧ�+���6*����D���̥� %�L�3�c�j�V��?GS�f`�	 {!*��C@k¤�A��^I2&��0)jߘ�%le�w2�K�C<�<볳ؿ���[;�K<[����V���.��*!��m+��Y0�*aD
D[WHE)���h��!"�3?~�9M�\I�a`!������./���/DH�1����iF�%3�焠-n^�U(��Da��O7_Ջ���׶6'������ڴ��pL��idJ��.o��oK�]�����M��`�Ř��>��9zB� ��o�7_��v����[��/�>����Q誊��/!�Ã��͟+����<�J2�\l�o+�`�D¢Z�E� 5~��$�d�F�-�k�}+v]�D7VX2�W^�J�T����i{�	�槣�!U2�bk��Z'��`�[v��kw�~�%2� n�>�{�8ҌIf$(PM�#�f0pD�4� &�����܎$t��Q^)iՓ�5������Z�t�i�a=�R�P.��	�2$)����<!���JѶ��1FcD@�hID)�T��"P��{�Rޥ*-�K�=�z������(�^�VN��BJ�F�<�u��'5�AD�O���[�q[y{FEP������PB������ws�fԁ��B$���0K56YH� P��8��1�8�ᵕAB�~i��s^���^'���w��DO�ZU��_�.��B^����!��?tf�����0*~=DJ%�>���Ŝ��[�yBN	77Oq�&�֫���k��/�q��BDPR��`���'����'8�(s��4M� ��j�����@M�yW������BS��o���3�(���Bn����\������nșaѪs �_Z��%�ތ\�1�������O��;�����]|v�o5�&|(����������9������<�ђ[R�1b��%�Y\1KY-~�g�7ũ?���@��y��Q�%�ף�(zvh���3!��n�;�@�����7b�線�F���J�Lv�"@z�0{�v@Ĕe��$�P�g5�V"w(3&9b�	%�`W�}��j�����#@JFN�QJ�`��P��r �լ����h�"�(�F�׷�>k��F��Z%�2 �)f��~5\��@�i&���y�R�#�1 F�u����"�!�keA�sQ�T�Ů?FFL� �ϧ�q'˵�H盡��]��8`�ce���4�e��1&K�9��
϶΀e��ʘ��a�:im�|ʼP�T��R7��{U�x ��h� T�ʆ�5T�/D@f�<IP	�o�������c)��%~�i�n�/K��C��nG�V`(j������k�gM�=�S���I�Z:o�v�TK�<"BQ��������equ��d�>}�y*H�#R�8�v�ǓgO��l0������)%��<�\
�	����Gf��%l���7u�,,�%�ô$�َ'9K�@�r����:�җ�3Q��6�h5Z�:;-����)z�LY�u�2]�r=� ��2�������Q��|y���ǃ�+>,����"����]|�o��S����<}ea6��՚��I
�-~���Xr1�doz~d�z���������j-a�3�W��X��L�L��1*#��e���5_]p��aM�5�A{G&�L`����Q2a�#2f�Z
 B�� ;$��5�02�x��F��x����0F�U����W��r�%	���,KZ�v���߮�sk�c	�F�.��j��S�-	�Z7S��pn}�T�JAI�s.AB�H� �(IPf+�4`�ڎA�%F����m��J�5o�HWR��{�'�����e�`�t��S^�g���JʟP��fL'��d��`��ք�Z��e��["�P5LXZ�F��s�X�n{E������9ke+��u�v�1��Q^+�sZ:A��.9�gJ�mW��E�����]��wj���/	5����p���J�Q����R�tx�iNl//��G^�~������ FJO�1��r��a�ʌ�xDJ	Zex�)�sO}���a]���㥯�k�;"��Ȩ��\^c��V��$����z�S�W����I�z�^#3$��6B���?���/������}��O��cߌ>p��������7�v�돤��?U���J:�%�D!ɐ�{2��R��s��r�~��K&o#�j�2 �z-6Ӕ���9x�ڼ�x�h���z�,����|�r-be(b����q,��2n�P��0}��S��j�6���%aFƬ3�L�2c���l�!�pG�C�ц�l ��xF�R���,�z!��OX])t�$����x�,�{_�V��1w�J�
��� �1a@ҌP
B�Z��X )c.Y3rJ��>�gD�F���E)+R*`hQ�ڞ�4�*������S_���5��[h�y��������0+����e"��Q�EiA��iz�7&2Mlg�$��0��T#+t���Ĭ-�ь 5�Ό.!K�5�l�n.�����ڪ�_)�x�ٛAsj ��v��
���F��I�7���W�S_��("]�o���9\Փ�����QE�d�C q@*�<g�R.8'l6#�FpQ�qy}��|�u���x�����}�� �i�8L38D[����	i^�,����3��s���Qp�F��$c���oxnI���J�\�{j5�:+��8n=1L�����\�e ��L	N��
I>�����0=}��}o���x�o��T���%���ax���(��G�|T&�Z��6�	4Z��K?�Lړ��k��S�Qd�� K���Xka���Xv�2?��Kq��/8��V�t��=ʿ%C�6��"F���������ѫޓ�:oAT�X�M��Fւ$3�L]�[�j��z�bε�e�vW���8>@���:C9#�Yp�����S6���εRWt��}�L��n��lb1�w `�)،f�
��֖��c{(KY�KR��X�%�eA��`�C�hQxUkKlԟ�n�?m��
��;Վr���G-�g�hԽ�h�*���! %,^��>FcQ�GҌ[��5-�7�޲��%���q�8�&�ڡ�@�Pڹm
�Ң���[(Gc+Dj��T���E�:/����K�����װ��Y{R�H���3��(��#pzx{�W���2o�C7ԛ���3*�[�@ss@�qq�4g\]]���#���8N3�d#T_{�%�~�d)x��cd���T0�qs{���{�a
��rFN�ĠYd��lRks��t���8Y�;����K���:�������H#���ۺ�I�Z���~���B[�f	�"��A(vn�:m?rI b��t�^��/��>���;�>��ۿ|`
]U������_���{~����h>��2A$�g#����	�j<]!@� �Z��&&�-�D;�5i:��d�V�D�P������e��k���y�H�b:������;�[Љ
;�Ӈ:�KA1��0b[�Q��)����ژT�@�2*�n�aP����lY�(�R$HP䈩�"˄P�B	�C�Ad��$A�%=����!�xe�j�!<d�Bt���&a�1)���u��{+���E��qq���ŦTJ�BEj��"�pE�����焒	4bX:X��Ա�@$BΊTj�
� I	b`��`?�΄cV0�d=�j��P�h�0�e:��I��v% +ͣ�̖��R
��.���?ۗllPh	�U�	`LK)(Z :!ȡ6	1!�4����$"����JMk_]�F&k-j]�
��l����������4�����	����E�֑ �)YIT��ֹ'���ւ����v�m[v�,�Ѣc"]�-L�:�gevF~�>5�n�Y��+;��i�����w�l/����ݣ+l6�4�����f��^������	�b��<���,'�x8����r�m�{5M���#'
�}y���vΔ�q����L���g'���t9 �o�u]����C뫯'��Z~�U�؜�j�$��I~�������������߂����|�o�-�������=���I���t� 5���,Ѥ��-q2B�Y�u�A��ن�W]j��.�`��O(������W5��w�Z���|�$윾�Y��\� ���7}A���[�U-.W։)�M�b���,����f9X'�b���-CY��?:���@��:C���L��E��������� $�Z�o����,ٺ
�nNUa��ߝ%�����D�c�E���m$"d�q��fQ2�T�p HY�&�D"D��`���5z*�\�X7-����o=S<>�K대dzZ�*ζ:XNH�ԖF��=��c��Z9���a��\�Jw�)Ag��^"E! J1_�,fK����rWB����Lw��(�Evk76Hm?��[	(��a����e�`�|v�������a�Ӄ�&�E�5�Q��f��J. �}�j� h�H�S�f8�Q��q����z�-sga�Z�jkKZR��i\ (6�t6`ETPJF�'����#����a�-B���RJ��v��	2�9c�#a�ݠd`;��n�SB��)8��)M�P%�J�!�,,sKe��{�x>I�<Y�;G�����z���c��3���Fw�c/_���>
����:�	l���a.�24-�D"�%A�d��_���y�}+�>�<.}>0�>=~��똏��W��GJ:��Ɇ���#���T�]J��Z��5�^��K�.ٱ���ߟv�[���`
y�1�f�)�=v}rg_��(],����p
�u� m�.�bD`
��jrגd�(�H�ſ�P���EfZj�U�u���Z�EY��U�	a�#�	*���H�,�ea������DKM�Z���0Е!Ж��0�H(�\=j�GV@R��j�s�&��J�zܘ�$"g˼�LP@����Aр���@V�����L���18��ߺ�qCN�����CS>��;���@Kz����q��ǵ�U ���mF�V�3C�2їw_�Gv^�a}�hM;��Ty���"���d"Y�Bɦ���-=y���=�P��� ��"+O�5�i}�W�\=c�)�O�w�V���*I֝�t�m?\��f1�g��i��[_��&@5A���^�j� ˄i>b�#�`�MeZ.���߁����A�f3"��'X�RPJ�dWǨRs�Ob�f��f��}u�V�ק�)�ޟ��q�峽�����Ým��xr�r"_t]]�Ƽ
 *���=.�2�1���O�g���?|�����	�������UzH4g�o�B��$�w�:9M{)Z������dP9��E���U��Xj?������[��7�*rfMU���ݤ����sZ�Z2%���0%�Ɇ���&�B7Nl���i$��5��דs��SR˜O��:#�D��#����<�;ͳ5��d�&�N�������`j�nBAd�z��^/�s�B*�lXw[k�o����[���L�o�m��a� �%�Υ�Bd����T���U��CR׮������x��w��?���Q�]� �����s��vJe�X������֙��������J�+b�!��i��[+�:e��#v-���K^Rm���/�ql�^�:U�
ъ�4/{CZ��v����7BNAulks�AK|v	�-�	�>9�X��*��_���-�R\
3n��|#����)��A�@ ������vLs�������^sr��@���%��n�#�<M�ӌ� ��<�w��u��{KM}ϟ�����-���'��:z�*���V�ja=TÔ5�Xȥ�L�Kӌ m��@Hy�.�����|��o���>�m��'�s5�Z��+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs����|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�f:���E�s�.�L����)������@��w��{n�<��D�^K6�md�c�pcs��yN���I]�$�����i�!�����9�x��=���b��ko@�[��E�S��y�a1�F�bf���W|��	�64졻V�#���޵_���d���є\[���0�h��9N�	���N�!�2�}���2c��?�ߝ��
���{��HI��z$��W}����7S��o=�|ֶ�����]b4�3R. f$ʠ̠\@egJ��%�Ȼ=�T�4�h��]�8T7�1�j�{ȷ#�i���f^���=�d�w=ܲ
	�1Hg�|_��O�Zb#��cE-cm����>AXj��T M�Z�iF��3ي{o�GE�z�E�8c�v�7�n�6��e��I-����#qs��F{J��w`f,�y+ �׽S��=Ӵ���Í�����WV��H7h�!�kO��6վT�#��N�l�N�E��O�2��e9~-�����!�xS�U�׾�19��?W��NH�w�ȥ�"��x{a�p����Zĺn���|r�j������!,}��}cu��o�2�T�6�;�n���1tKY�&�!{��1��]�}zߺ�F��t�*���ER;�H�t����ǯ����z��d�a��x��iW��Hcx��-`�*c�&�b�ns�z$�o�g�{/E$\#>����ЅQ��HIM����+$'�4AZ2O~� ��yM]#�ߌxn���%���L�ځ��ہ�̣��c @�b^�l��1.��cch��}=��&4��ƒD+oB�#��G=t�b��O�Jid�m������>uʫ��C��i�&�T+n%+n圁��){4���g�$��J��kB����ͥ��V�ƃ;�:�J]]w��{�X�?�:�&���=��������O�m�j���*V�����*C�=,�!���*č{��UD��������ݣ��q�=M�\���58.ɚw�iY{���tG����U�-��~���7�O�o~�e���� �il0�C��Ъ��m-r�� {�sB*;P�~�S���� ����x��:П}�{���9 ���r~+��H�X��ԭ4���}�o�@j�#]�^�*$ [KR+�#��W���s�Ƭqtݱ��m�|�6�]�ݲ$�|zYh[=�=��{zQ���f`�{CX��]cX=
�եz�e��i* 5�¾Ag"$����LDA}L����vA��!�Vo��t�2vۤ�o����j���ĭ>�s�����Jk��\,fqO:5+�Y@�����`�083L��&1���e0+r��guU(ߚ=�/��N(d1���WG�1!� �wX��̽���z�ͷ�kߓ�XQ�d�:x����I�H#W޽Y#)���:M̢���t�܈+�$K�d�f�]��D&I^�h9��� M٢>�w-���ugQ��������[�˼`�ŵ��ͫ��}{{���F?n����%��m�4����>��	�s귕��WHպt K���S����TPe��Ċ�#�ہ�Z3!g��tlW}k�Մ,�c��xh^Dp��Hy�Ϙ�)\ER-Z'	@�>Q�ڣ5↳�BU��?��7�������a����^{3D��m#�2ڂ\�������$"�w��;��9�8A�
��r��\ (�N`ڻQ[@y��Ȼ?��?�7�����?�7Ձ �����_�9,K��n�JOr��ip��0���P��NԚ�x!ء�:*K{���G�������c����_���pc����YĲ	k�Yi�L��M�0i�>�O7�77������ɼ,�l{H�7�Q�L�F&��5ܷ�R��0�> �c}����5�%��� 6���m8�/�Nv�j�$~	��A]<a�:s#\WEU=������hJ��-R��y�x>�Ɋ���p�4N���*�f�kǆ��q�'�:G˩E⑏��5�QJ��E��k;������0<�/tv�ֲ�"�PuHޓ��i�l�����'���f�71�:�^��)!!�Y�F�i��^��̮�X.���R�.��*VX^�6�Zl�^X��t�Ϭ�$C}r�n�I-��g�����]��^�W����X�����ӫ\k`�f
p̌R\��>�4�h�v�UR��5ۏjkX*0�Z{V6�͕dG� �_�{���P�u9�I��E���5r3��#�Q���-b7�"]���=j�Q�d��^6��SF*djp�<d�X�4y�������t����w�Agq�����~��K���7~���NzE~�HY���h2�7���rZ=��a�]�o�2�����,k���m�cV9�߬�'76Y�hm.pϫ��Pݶ*�o`�y>���r��e%�y�͐t%� �V�:B�6�I|��9#�y���@N	3^T}x��i; ų�ÓD����5�{�!�l��彘,�^$�)2Ī�uV�M�M� r[<�A�J��`��ŕK������J������@�N	�^��
4��Sww��3�^[/���ӄ=�8��I���Z�:�����������>+�X�����:�^�u[���՝t�+�48�b�/��	>�N���SO�)�&9�5�~h+e0'��m��R�C1��ٌͨ0���z��A��g�y��������@"t��q���z�7�\\��Ū��Vḧ́�ך�_l{�=�$�ު���j\�J���r7������f`8@�V�	)OÐ�V��d3�ن�����u]�P<m)^i,zlp]��v��{Iלޮ�n�l��gA�m+���Kߺt��"������ϻ<��2��	x% R�(�<�ly#�I=�)!BJ�א��s����2�^���A��xS� P���o{���?��~�����|K%��M~W�̓���0��F�Эƞ�j��e{�����@�l��l����]e<�}'H.[�19{xh�gW�z_���
�0�y1��؄�Z�W�ZG����f.���X7��X3#b҂ H�$s�x�i&{���3k��!^?K�ٔi��@���u���:�6a��#^6�x[�sU y�V`n ��y�P������h��=�f���\�b���m��	˲@!�rBNdS����̣*��|�K��]$�W�����f׍y�z�c�S&�������خ_���[���ӱ��f=�����}� aW��e1/�<$��{�잒��!�Ecm�׾�\���@+�2��<	��$���,�v_�쨧��K�6�MX�/����ֵ�][�_;����@�/k�}���~��x�ǟ��vcٌ�_����o�=K e��6�~Y��� MpCI��n͢�Sbp���^Y,(@"F���ڈ��LP�H �)��M�3�،G�{(6?\1�q[�G�H��U�p��9ҿ�h�����8�8��=j�w����!�c��E� W��8O�#�8'(gP��T�<�R�0=��~2��+ǫ{�=���Q�y����~��﨟�9�����Ͽ��?�����"G4,X����C���IA ��۵J�ԇ���R�^/���O�6w��鮘�mB�:�D-�	�.�V>�sQ�Jzh+���R�2]�!�ILloߋglZP?_��IU��b��EO*�����t �4r��mU�g�{}�ȉ�h۞���?��26�5f�!Cү
�MR�Q�Rd�3��n��{���K2V�,��V\^6<)�L��Vۨ�ruh�S �U�d�3 ���խg�!e3D̨i,:��յ���޻�cܧ�g���ՙ��z�F�9��SztC��9z����~���M�A ͞̳�1r�������WkU�|4e@���zw�}-[�;�-���}
��]�2�Ț 9����ģX�0���y�\�|���q�����#i��n?-g��=6�k=��n�z��X��kU���4��"�%'L�	9%;�`�L
挤�T9	@�l�Fk�4r��CY��
z���M�B܈�\�H٣~�������zQ�p��������7�����zU�Yn����n���zU���{�*m�ל���@��(Д�����7�\��mJ{ ����ɟh��}���aqޤ�it"�~����Ư��q�����OO	��1�H��֦�^A����e�B�aH����#T�k�]M���C�7��ƚ�G��.[WF�yzŪ=�ݳ{�_�(Z��Z�V��Y�_���'Q�VJ�D��Z����3�0��t�6v�����"����)ﯕ֜��ٕ�n�9n����X�g�W�ۡ�s�.w+�:Q�M��s���e��+\���-S�n�qy!x��@� R=�n��j/SL)#1#�Aa�2RS�g��L4[;���抔3���L�\@<�6����h��q2���zR�b���M�j�7����Gd���{�CZe�EٚK6.b�֘�(2sF��BW[ߍ�
2�L�T��y���!����sF+tqt�.��y��@/�Z��wz�Q<�]O���zM����Y@���U6��d�{�Q�p��l�x3 s:o�!o����{�Z��li��~�4M`2�k��b�dbO�JV1�'�ͧ�l�*���*cؑ�v9EWEi���O���Q5�e��`|@�����ݯ�*�D7��X�vO��,cF�f�z=Ł�ߏܻ/w.�^�z:]�L}w6c���{p��yO{����0s��e������ `�(~���ެ�it CB�s�(�|]./~��<x����0��ݽ�q�k7�M!��湨����z��u������X���æ�lv�&44���%��t�9��#��4<�ѿO�屛��L�������y�Խi �40��v��`$O(��K��;�m�%v��IM>��=3*(�9�++	�������ٟ{� �:Q�W�JU���QEէn	�������Z�
hJ�1-G\��oy�Ɗ��ZQ[C�L���PB.�zf��y����&X��V@����ē`i���PJ��eƝ�~���W��&�9�f�mk�p�)*�zlN{t	MҪ7��w�Ev������aHٌoej���v;�a�r�l:�P�6��&���N;H���A@*;�i�@��'s�tq	=��.�8����Ji�n��a3�'7�ӣo�`$�\9��#���l���#2�kH�+���p�ѝ��Þ+��I�^���}�Wd��[=���m���b��n����N>��B�x��-��V/n�����G�9m���\�\zAl�
jd����å�>i�H�!��G��,����U~�������H�)Rqs�~�	�ŏk�EG�f��;@��kDJ��C��Ɣ����2퐦�T&�r���i�������S�����7���M�M}�w����s�(>����������K*�	Q����˧���9���e�ՕP��=r`�ʔ,TBCAZ�^�Yվ S?�W�����z�h-�R�ԳC
O���Gچ�\�]�F�����Ⱦ �(�a��B��@�)���j���[�	9�0Q�!gܚv��.pQ�8�=&-��9!��vJ�>'�Z��ۃ��d�ѣ��MW�z���am�{# *r�P�̌&�|D�'���l��{��	g���A����V.�Z��ǓU�i��3�
�Q���a���	mO(��e^���b��dnD*NMq���'2���t+cAc=�t1��}3|��^�E���t�Ve�*���E�x��;��}^wJ}F��NH��9���=\��&{b��кN�y<�i�`KM`�ВВ��!*�߃�'!w��g0JbdΞN�ϚR�y�<��7d��(�ի����U�&��[����Nڣ?�Ag uY0��=?SA��K��郡l*[�N�
�� M7��6�<��#�,H�L�`ڡ���&�,�V�'IR�tEj{��p<][$*O�i�z��CS,�tid�r;��?�z�9���"M�������[Ov�)�S�Z��E�v��6y�.��3aҸX#�}��+Fl_�}��
'���#�����-��:X��D�+�?��2A��\,���`���:�>ޖk��G����S�7�o��C�3�0n������^~��9ܯi��+𣤺K������|�%՞�@nM{ۅ􇗺����V����V�@�W��X���K��m����xo9a��Dmآ�E���ƿ�W;���	9��5�o]�@2#%�BJ�����[�`���T�����3i�e������%v(v%SvO P����=����U��>%�BA���H�_o�̬Tv�DBDJ�oӴS����'䴳��4�ݑ[���Z��¢�V�dJzJl=����`�k(�C��&�s<����&03��Ќ�)�J.���-|�Kh�Q���D6��� �	�+�d��'2�'�����б�������Ƴ�j����ѾǤ;����/xލa߽)����?�+T��n#]6�\lP���*H:���(B"�5���R&P�x�M�4�����m*����S�˧�r@&'�V��o&���5ZU��`���Ƭ AM�A�H9�%e&eb]�E[�*M�*n����������N|�����M�D���'�UIDIUHd�Jċܴ��}��.��0�X�R�)_�̱��� ��?y;��3)Ӕ��_@�p�X�()�	cވ�Z_����dެx�@�!���RaKM�}��M$��IU��u5�!d�(�5�;F��(���F��7������7�S'=`�=#��h��SA�%���r�;�:��ns�3���j�������\��|Ͽ�����?1�2: ����_�ٟ��˸������{�=��$���酪���k��+���q�����f�KI���ja\/"���zC8b�=4z��r{@������G����xiKtE'�zPTm85A�#�d�c����>)I�"��gMH�(^�iyfFJJ9`��\pk���t�|�|@!k� '$0)Zv�>�����������S#JU�-��DG"����> ½�t���!�'�{<pՓ�^K[qF������
9��*�*�T�lҞiwU���v��}-�:�'ngpR�Xt�@p�GiIN��2��e�t\x8N[D��v�D�����E#B*��pk���-­���.����yL��X r��k�ivD�2���MWA���vf����^�E���Y�U@�!��. d*����
��Ҿ��4%�\4��!�"������3v���O@�L��K��'�O�佧��̤��&�ĩ1s#BUEm�.�<SJs���r:��� >NJ�>щ���隠G �rﵓ��"h'-j�,`���W��(���p��C�])�n�����>�|	�U=�&��-mr)��փjۋ�I[+R[��L��$���"�T��HZPX�XG�\���).��)��@�KL��Φ�ժh�J��Ac�>TB����H��nl,��&P����=� �
�V�Aɮ��;�ױH����}���I5��u�g���)#�؝��*S�g���X�H��{��}�E)�K��7��v~��,�Q���w�9���G?���
~���=�f��˷ԁ ������+��q���_hy����m���<1��k�/Q�"%ki�&Hb�0i�N�:���*&X�ܛ��x=��hxI8������V7�U�C&`l �U`Q�PSA&��V�'�W ~�0)R�P�ȔL�L2�0�f1QA��r��i�;�ܙ�`���<!���VA[`�ښ��Y����T���<�Ӄ������5f�� }�2^d�<����h͉+���ݾ*s��n���ҔX.�����2��r��Sʍ�y.Rk���&�eB]
8=U�߯����wcW���������T�E�ITx�j���P�'n)�4/x���Ǚ�JΦ���	9eH3)K&����S�>+n���pkG�mFW"D���+����}��6̨��m�.o�J]ꛣ�^�lm�Ex���~��Z�.���. �Z�����	uf�(�H�V��݄S�q:	��)���gԚ���%��ٕJ�n/|�����S��#_3�Cb<,�����_�į xE��,*ߨN/��[.��[ޕ�)7�,�rc��D¹4"m��kd�e�&Mx7)�De�k�,�jEz�Qr��m�@��r}dL�y*iJ�K�Xu�mn	@Zj˵�,�%�9Km���V淋���R���|�H}mym~B��Vkˡ-ׅuIB�mAʌ�����q��i�����B�N��]ɸ�`\��КE2
d)�vB����hb:]��HPP]Еۈ H��u�Ż+]�����dE�"����Q�;��'�#u�BDS�;oM�{爌Z�q&�a>�@0{�>���>xe�R�#O{�2]q�-�������������R�9�-x�v���Ox���_�{��Oѯ�ҿ���A^�E�� -&�)&<Cb櫶il��R����D��dZ��\���lz�{��f����!���&N��@2AQA3�넂v���z�����+de
��M�1MH�=�N9{�3�JW�c���].pw�w����z*C9!��Ҥ�,Dt��&ί���Μ��S�\N�O	��*��9O'N��ʇ%]ޞ?�3?]�|��r��R3���֟Ih�J���n(������-���Vlr�js�L��'���������9\\�5��Y�q}��YQ�KD�[k���i>��c��[A*Y/��P8=��J��e��yλ]�23@���5��ä�ĉh_wD�/3������?����²]KοNە�9���D�`P���F�1Е�[�pV(�GE�B��:V��� �MՆt:i�_B�	����Δ���K�Zv;�ۇ��R�I��x�s�j��P%���y��SO�r��xI�o�i�Uʻ_W�/���
PK�%���VJie�qj<q�����7e��[,�"��y+��v��	�fc�T2���tЗ#�X��'kgj3P��5�S�L�z���Pv�L��Ί4�EZ�5H���P����"�a������u��Xj�3Z�2�_��m^^���h�۲�g��nk�����T��z(:CeA[ԥ�-���e9��#)���.�*{Bk��:5��m� ���־�D6��SS��' $Ӽ��l�J�#��vng�k)��0A��}��1 h����n<EYi7587"<%��Z,�;��R��xJ;K#��W����^*��J���.>��[�����-w��K���>���4�˸n����?$*���/u~{�si���fH�!��0���n۵b-�=�
�<�����L7��^ �ʱb���߱�l	�W�pya��������+�
����`E6jU��.�֐S�R2�2!sƄl����1+ Ta�
�|�C����%����gO�6����v�2	8w�_Ki����/�gSΟL)����IR�s޵��V=<�T��'>����z[3CiBK�' �g�y�o�z��W�
 �ZѤbYf���=�����^�ƽ|��5?|�Wi̜H[�Z+��L�-;�tGTo�����E�u߄wJ�������rI�3Cs��I�LXTY]S��'��Ki��T�%����z,,`�jR�["�*-��GA��L{�`�-�z/�C�T�R��fPv�RR�uG�}k=�ѓ�Px�&�U�[U�U����Y��ki���R[b�K[�R�)�:/u��~��ݾ�P3�ք_���|Yr������?�z�g����4?q[�p!�ť�|K ��}�SH�ۨ8y����l5����5���?���x~���  �IK���eF���!��m/����y��Nz���г�������;�����<�xWP��@��Y󤏧X�+d�RL�XeW��Rk*��tD=^��%��i����������R���f7�Y�t���A�0N��st���6C��P<r�3�X�\� `��X���/�6ʀ���ƞ���P&Fd��N6��],���H��i�������N����������Oķ� ���G��w��~	iaҧ����.˿�d����&�TZ;B<N*�y7��f�M���G�X��+?Yŧƞ]�.�^A�!�⣴�͏Tتe��ײ�ի������z}�Wu����
h"̲`>��Dؗɫ��r�dNإ	S*&/��g�j�(�w8L�qQ.q�p�������S�Ň��ʴ�r�ʧ	��=�_�����WN��i*{-��|���~���r�0��	���	w��^�w�RI8=8�x\p}\���}������Z�ڽ{�ݿ�w�S��,���=,�	��D��,hMH�uB�ɋM�D�o\1e��.�rb�2A�k�+Q����c�i��~�wW�ֻ���-�N��d�x޷$i�95��Ě�sK��wAV��&a�=0�o�{�M�7\!�*)TD�6�(�q�nr�n�r�ׯ<���8����^�_k�
�gk��.tw�6P��2��O��/t~�{��S�[O���3�[���ew@��HE��}�F��7z������~�+XN�X���f`>bz�I��5˼�\�$e��I�i�z�b�E}7P���4�ҔT�����j|k�C�j}�&�,G���ꅔq<U\_/&*����4pݴ��6�c�F}*�����T� �#&��Z�u��Zunqs[|C
ٍK�Q�H�����5�m��
ǽ��vS!T�^�m�ZJ�۾�T.>���.��?�����C�,���#o�R�'�[�@���/�P2�_��SU����j�ai�;[��&kaZ���R����pk5�9Ϗ�$x.�+m?��O���#޾����6�ի�{�+|���k�W���Ҁ�r�um�>�S�������*6PD�]���p�i��~qUP+ �q��;�{�$��}Wn_�zpk��������y7}\���~��_�}��اtwH�����l��t���^���Ջ#ꬸ���)�N`͠�P�x��5�EЈQ�RFk%��u�_b�9����6L��z���X��^~���p��C���ⷿ�{s�U��g>j��`��p�O?�=}j��km~?D_$�}����\?�;�F�|��x�,f8���"g�����Ԅ�i�i^��+�
���r��;>&�%&y\=�]�pm{��u-�+�P�yʜ���M�Ȥ/{�ڏ�o�~��P8%3+��J�B����bG)#s��8�\v���)���xˋ|���?5���Η>�1(	��5�O?��?�aY�����I����iE�I[��XߢV�0�}h�o�ӽ���X#U" �/���i�-��ke�"�
WU������#��W��'�bC)���QR���(�$L����!>�b`�&ȑӄ[��ؕ���jŔn#c�D	�/���~�ٯ=y��������n�����ҧ_���$4��sϾѷ4��B?�a���{
����an3Z[px�����{���%Ǉ/��J��K��Z�k���bAkC&��^�M	�
�B8͋�N'@��i3/W�Zsx�����F%\�I���+���'�9#%B���d����)���pLލB��Z�l#Y}��	 2��4ٰ�4������k9��J�WA����>���8��-��7�������@�/|�ؽ�i\��h�G�y�����^�N��wf�ߩ�h�����Ui{�Z �Td��^��G��7mܫ��#��f���a�
}������J׆������,*�#� jC|��I��WhRQ�u�K���%d6�f���i���U����\���w��;O�}�c��̻>��/}�ݓ�s����p���7�6A ��_�E �VA�3�y��镯���t�.>Ȍ�6ײ���{ҖI*�r�2� ���s�>m�P���ٔ7��@��xS����]�>�
U�b5�UKIu�����e�i�GǞ�2��qA�x��y+RE`���{ΩW��(/�r?O��r��/Q��H��r��;���/E����=�;��O���`y������SO�vz[m�gAx*ߣ��Է�ջ"� �C2IUXUX��h��d5�㒮��R���Ůq4%+a����{�}�EM`B\���� �����MLPb7MP.>�E-4�4�\�����������������O��,������e���[Z��?��O �^�����>�j~��[o� <xG=]�u��
�>��{���і;m^��T8^�Z5u����54��mmV5�&�'o
�v�k�z#�����3!�U���(q#2��ܵ!o(��p�˔�g��I�.�,̩��2_'N��k����?���?���^�� ��}��F���t~��[��?�ҳ��P��׸x�S}����[h�Ro�N"����P}Z���[*8a�������խ����c_q��
���7�.?IB�,�m��*����>�0��וf�����m���5-˂��Jɨb�1S.Z�W%O��������px�s���/�{�ٷ�-�<�����o�� �g�ԧ���x�|��� rxn�,�����6�<S8�J�U��o"z��o�N�Ts���(��yO
�jz6O���"������
�6C����ܭ-nk�$))aۤ>�i�2"��2%%NB����J�f%>�
����K�ӗ�����qY꧙���F�^|I_��R�L�Uo{���ѷﷄfw�/|�v�j5��@� /����#K]�&�h�Y[M�IRQ6�g"�邈n�-�iOL;UL
ͤH`Ndc���X��J�d�G�*T�`�FB��5���B}�+��De�8-3��#�*�2�~�'�V�J�����<����������O������/�u�4��|��ѷ"�JT�}�8�M����p��~�N��p:ͻZka���:�D�ۙ���������nI�Q�h�k�y^��T91133)"�b��f��@�Y�Z�\r΀���W��X))1	@ں�-�1QQc�
�
�3���9�gN���U��N���,���>+���S�S^��N������¯��'�
�����w?�Y�؏��}�� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��1�Ӓ������   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X    IEND�B`�PK
     �)K[d��   �   /   images/a262aa33-74c4-460b-b0ad-c746896f6744.png�PNG

   IHDR   d   d   p�T   gAMA  ���a   	pHYs     ��   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X  �IDATx��{y���u׹���Z�j��ez�����L�b'������2�eH$BaJ�@�dC��`�@��![G6NlϒqO{2��=��RU]{��ۿ�����1�'��n�u�{�[�=�s~�w��ʥ��1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�l�c@�a�z��Ti�R��)�|�H)����]ǧ0�Vg�¸K�F�Z���=:0��y��8L^a�&����4�"ϨH32ʐv4������>Y��6����=�n� ��w�H��)�~�����t�g��!�<T~V�Yz`�����j����ר�����Z�:@N�NF�ޢ���,S�ޠ��NY<�Zk��J��� m
& ̡T�nW���]����{}*f��>s���m�ݽ㯐[����u��)h~�����>�����R����h_�М�NݴC͠���ޘ�g>�?���g�~��P�R8葉ڤ+�T�O�8�,�`�UZ�	!�n�6�a���y6O"ǭVk��D o�D9~G��[�m���^�u�'^"�[^���O�N����+ DF�u
��v�����/M2�P���&���8\��
\��w�z��V�K3�K3���h㇟|������~ݟ����W���f�ȉCD�M"�!Y֕�.���n�Sf�	ch��G�&�q�H5���*o/��%�ݼIj��KI�Z����.J[�(�\ׇGk2�j�4���X:
A�tԿ�M?�Yg����K_����pkC通K�23�*0o�g3�$����0�v�g~�/+�W7��|��ּ�,un_����� I;���\��u��_},�~�n@"��-ob+b�v��X�I��f�L]�Һ^��U�8�E'?vV�x�C�k�;���M�}$�DLi�S����mQ�Ņ�:��(_Ug�����F�����	��ġ`VcrDqf*��q
4SU�NLm&U^�������G��i�8�3�.�۩.tؙ9|fp�[�D����W)�lSg}�����ѡ��0���%�]���pa�[���>PD���~󧢵�� �v���ԡ�����?�j�UZ��ε��@��_
��e���,�=McB�'�pt�&���.���
{^�K�zst���t��I��#���\N������r���4a�8&:��i�M����fS޻�0�*N�� ��%
V^��'B�%���w�1�@��Yuh$L�wQ&�0�3��	B8f��e�wA���Hi��%�?�p-,$|M^�0$ln���ÃN��'���S���;u���}���~g�| ��eP�>Gӧ>�����)3���I�+Q$d���򼴍�*ձ�aѣ�x�M�"D�ܤ,=E��Cdẝ��HKb�=~���kur��0!�-�)���!��D��)�px0D!�`����!��YҞ+sU9��x�T�J�,�OR@do6v�"�J��:������gB�K���E�����Ԡ?±��� ����s�Kh���+��7^mn����&]
wV�:{���i��u�Z�|�I��'��&��=�{��֠}m�r�<�r � ��c%ED��*�	���8k�0�Z��5�׃S�w����i@�g�ׅ�âz��w[�D'��I�Ar<��a�L*�އ\M����G�+�+��߰s[�����
��T�l1�z��=��.� �v+r�v��[�D�KO��c�	�K�N����[_|���S\�m#$ł��y��s��~)�oR�"�qm�ߵU�/�ԃpw��
"��U��2��Nڦ�<���w]B�^�X�U�F�ozZ�3d��(w�m����&�ҳɂ�d^J��)$��D� ]��X0�*\KIy,`Z�S�oا\G�څ��k�ԫ����G(4ED�+�i8���\r;Y_�Fa�bn���V�`���܉'�n��z �}G����#7��{�B���/ga�`:��v!{�%Z�A�q�P�w���~CYT�UM@u�C�D&�����m�O���KY`��Cs5�e@Q�f�\Z�m��-�%*$4�H`ٟ�i2WD�L]VCq�)�~�dQE�:�)IX˵喝
��O=E>U�)��:[[��Bβ�saȜF3�`H)E1��>>CN�?оs������=��;k�.�$�ҩ��x�~���p��_Α7�p�&q�@NTNu����	yф���ά�K���	]�WQ�6���p^S7����N�z��7e�WY��G�95�F��+�ÁBሚ�t�D�,UX�/��p $o�T(M{5�ր�2�gBrNa��r����
�7_׃s̟z���S��\!3X#߳�7��0��p�3��<��D4��Y���b4~�:��˝�7^�H,P��J�ܰ�K핛tv�y��'�w���y�����a2UNQ��8���/#z��!X�4Ee�w�.���9��� �ޙш���.U�5rI?��H�>��!���~�
S%6Y!
F��[ͪJ�亢�"PNтĚ�Ҿ��\�*Ȫ"�윬c�*#��%j��}���y�����﵌r+���Q����5��#w�<� o`Nٰ]M�꿞=��3������i#$�z,�Sm��}ݕ��}�{���ޑ(P���̄ZP^U<P��7�E�)s��p� �Jg�"L��s���8=�8�&Q&	�A@����d��U��Z%p@ e�w�C�� jT���xbn�[惟^��.�ӶxmhI�R�8��X[;��Dn�E~�^��WR# j.�5�RX�_�r�+��]�ʜ-��"���^�t늬դ^��G� x�s�⿸���ԉ?��Q���:�o��� j���g㝫���8��/�(���E�a���r��j�Tܻa/k8S�PY$����I:9s��;��1�M��0RE��<�Rھ��DR�y�2���D�*��$�ETdF�(�8*4�uD)1{6G�����@]-��=F���r��q����0��؜(y�s����@onm/;1�y�&�'����YH��.�KT]xP���SY2�A9qE���	r��������������έ����{>�����@S��/�c��eu��ʘ���	9%�Qڪ��x�"�4a�$ۡN�o��t���"��Z�m�O�ȉ�/SmΞ���%���b[�Ap�����29?gi�IH+�� p"��� xH_�\U�#�8 �=���� �Ʈ��Π�P|9�G�ex����)ݥT�$��5����)L��H��=�c-9Q��3�C���"��BS��4�=w9Z~j;�~����i�ě�}Ű"a��$�ڝ{<��X�1x;"g U.�*Y-���$�0��=��FG*��wi�f���zK�l^���~M��!t`����E�ޗ��5@���R�3�7(T�rl��<��T��;D5�PD��ѹ���d����\�p�!ё�I�#&��Hn=�Afa������[�M�����ox(�}��jߑ5*8�ҷ��D]�kduƵX���E��e��g���s5��w: +�KaS��q��0Y*rc�dZR��+J�*�G�Zc���"4A30��7���ޯ�Q�/�޸D���xs��D�p���.a����6�9%�3ա��XYn�"L[�˭"� �� 1��MR��(a�F��Pcs�6���w�UD#�ƴ�k�:&g�ɻ��P����]^[U��գ�W�s�%���@X���f�S�?��:	���.�B�r8�魐��57�ڛ'�G�͢�k�$�\.�Ӳ3�������|�R�|�|�܁�ڴ���P-���ץ�+Qhlo�)�^��˹!;�S��1C'�aT����Uz+�t�$½�;j�9�d(t��x����m�0H�Հ�"�Yi��BT������5���8R��/6�̽L�FKn�M_r;4��<�\�؊K�E~�%ut���ص;�2��e�@4�����*kY4S���X/���9������
�Y
p=���8�8,Xp��ͽʶ,�{F�>Q�H�Q�Ĩ�SCsnF���g���T���胁őX���}d�$PJR�_Ξ)�
���֠�hGh[���j����'M1��'�>�Hd�D5��8R��,
k"�Y!���C��\Ŕ�AqY�(7��=�b�H�Kr6���e�Nو+_2Kc�����]9ڪ�£���a�Y)@+[3N���?�u@Y�I��2�a^I
��a�|&R��e/Ki�Y����������<}8���$i��{{*2m��"��ZjF�R9\ c�YZ���V�#�j)y�*j�Pj�T))6�����Q�Ƥq��(؟���Z�K�כ�ό��bЃ�l%"w6�s9j�k^\	�m��J� ą�|�(�MҜ[_$9��.e�h5e��ؾ�eJ�F�M0>ߵ�����C���W��4n�&8A�{�^�U,|^x[]��~{�/ۓ��S���r�*��VM:�Ibh*,J2�{`PY��-s�&BU�S��!b%f6zx�"(���u��_NM��ϯ�]	p���[ِ�������C(A��ʚ�&V�%n��Ҳ��m��XZ)�77�lH>�~X���w>�ⴇ�P8Y��e�z��>�!,�S�}%�[��˕�P$+!g�0��Qd�F��-¬��X5�@�iPE�vٟa�T�r7����hޅme���-�a�����Ɣ��;GМ��`��?��{��~�ɿ��'�������C�r.r��Hf@�޾�ѹ���J�ƲЛ�J8����1��� B.N0���=6ۈ3ei��0����E+<÷�V�sI���ϋ{=)�[Q�����#�Ap$�r��q�a(�`�FQО�Y��jî1��X�~�ʍ����C��V!��e���z�3�r�[)W�`�'��?�%��_x���gg�~�Gk�7l>�UH��E�ǡ.J!�dv��:�Ք&�6N���&�1�Ri3צ��=#*�!>�
�mI��P�{�0$j����쵲�ABf�Y֒#����j�����K+GDA�iy_dv�Q��M��T�b���xm.��P�vű|����g�e�X:�JP�W�})B����qQ���H��=���t{��?;�U2�1�	���`���'�~?l.���!Q�w+gD��w��<F��8� ��#$�I�G^�Aa)�un��-O!
c�	����ԋ
�	i(6;��R��	�����|#M�RJd�sRa��
VO^'ANL��Y�k���PY��6��Z��<mMf7�4�t&{,E)�*v�t$F[��1!,�Y�y�s������}2;7YW�����c�q�u�x��T_,.y�}?}�y��,�Ӱc���Z��团�`����)&��|,Q�%�3�Z�T���OD�R����M�όy����|DJ�s�<���O(]��Yx�L�|��X�ǀ�ANY�ؘ 2��H0/n]��z�̍�s�B$+D���"Ys3�T�
Z9?�`NY�h$�(ͲQj�cIQe�_�)��T�~.�t�̳�z�U:�����!�����(��+/�����_s���n�E}��P�{o�����\P���r���J*@S)GG����Ae!ȋ�G\^���P4l�ݞO��+�;�,�}!<��F�R�L���=T`��v������[C�����8/QV�I��@�[�%���-s"� d����uH2��<�P1��:h��gI>�b��I�ѯ�Ch5�������7���st�]��\�v�~7-_x�K��c����YtH��O�-��:�F�"iK�\Ŀ�׏���4�ϐ�x��
�d���Y���Oi+���V���!���h�w�e
 Ң)�;�YِR;@nom��@O���#&���V��UBq���ͯE�.E��4�΂+�5YO�{�F��`d�mp_>��A�Q/���t���h�(��;�_�Ï�|���|����k����W�n�u�1��H꿡������H1��;�^�[��dQ!G��Ȇ2�@qN��A!)�k�ҶVE�V��u2��f�u�k$xn��(0p��]6�F�DSFF!^���+
��l��?W�yn��\Ԡ)v(�6�r�u$��k�
PEO!���$c��'�,]
�Q=�st�t�\���ׇ^�������yo����G����!�v@fg��k/����?���������S�ҡbЅ��e�~i+e%BVG��b�f�n��Cb,�N�w���Ƚ �T�k\�K��'���V��h���]�B�� ^�>]�����lM+�wJ�2u������5)Ly�2�MR�UI5�}��L��k1����k�	oN9Vy�߇�#Y1a;T�&�.����í�~��c������c��i���?0��e|�)�u�T���[itď��FC��'�Oūx��i�\�s����3Μ�-���'���*��jו�6$���-��4��"k����z��J�Z��sը�Pvo]B5��\Q�{߳5�[%g��ٽ)8�eC��0�,~F�_�J��@t�4U�*(�R��#��>�M-�hQ�3�܀�t�m�e�l�a=^s��������~�wx�̇�w�������K��|�vV.��}�?���?b��;����"�e��=�f/.��kT_���En��u:��!j֏H����V��|W;^�K���MD���*��4���AUy���Ss)�f������|��#;���.�u ɎHw���.!��#К��BZG�����8�%��N5O�zGSY�u'�}����O\B� ��Ȯ�H�N���a�'.j�.Ҝ�g)�#p+Ti-Qe��E����a{c��n.�������ճF��w6�S'�������:���H�}R�sn)���>���z�&�3�Uϣ�?M3�����Go�V�3����W_s+��&��N/�G�+���Q���Yz���k۝f�f�����@{��㙄�"����Ju��9�r�i�v������������X��� �:��LT��N{�/)<L����l߭;�f�y�5����ߗ{�<r����.��y/��^"�@�ZI=�F?s �<8^0��U�s���t�s;���H�}oJ��y�V_y�q�����d�����~�v>��n�%G GS+]A1��4��x*�������D�ۊW�=W��k�>��/]�򯷛G���	��P�_'�*�.kqgv{��RoQ7�d�*qR
}EQ��0�і���|�>9Bൕ�e2�-�i��,�bؕ=>'K�w6h8�KG��� `<PRvP<�)���y���?�ɠw��G%�:��=SSt�0Eu�婙�H�Z��S�z��M�yם��?[�N����s�<E5�X�����w3���}ȁG�CwΝ�J����is��*4������V��6}���ȼ���T+�����ڌ)	w�9�_����W~��W.�C��%ZlP-h������}/^�L?N/|�b`|P��֚l�nܜ��U�y�ؗ��ڇ2�[��}�[����<t9`@K���w:�W_���BՇ�{典H�o�4�f��2-��_���[�p�C��
��9.'u!\1���tz�5|�|��>t���W�9��D<����Auߙ'�~�s�"�?�7i��D�����G~��_{)�]D�D��.
ɵΦ��j[Mz��ץg�͆t����q����r�N<�m�W.~���CTi�݋�%�W�ƉluKu�P����FS��5����� ~i�~��wt�?�}�w�����O��O���wf��c�W�c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2f�D�{��w��    IEND�B`�PK
     �)K[:\�iE E /   images/7be072cc-a725-4446-be13-eff8a797d760.png�PNG

   IHDR  4  J   ���   	pHYs  \F  \F�CA  ��IDATx������?��ofw��q�ޏ�"�E�] �$�1��wM�'�c�IL�y�c�`�A�Ă�w8�z�3����\r��m=��y�n��ۻ/�����~�7>P��[�G�����Q8�v��Z��������������R�pZ�_mpP-o����E���ac;�|�D}`��p��?f���:�s�8^~�����I����O���=��TCݶ�.?P:o���:8X�y�=_�h(�3�_(�(���ҙ�5��O0���������������`��\G�e�*�p^�ϣݷ�|���R3аt^	l,������Dp�"""""""""""""�cj" &����B���e�����
P�I�@�c�"(>)o}6f�<�DDDDDDDDDDDDDD^��9�9��{����CK���J;(%$�a��3�J�q��W:��������������H#���ƹ��݃�y�a�/��	�Ԓ3�p��&�����\N%�/��*,�+(��"lq/�Y�4()%W��t�	�^�����8Q��0�3�箆���k^\J*�hp�ʺt�ص?��@DDDDDDDDDDDDDD)B�
�Qz������U����a�ܙX"~8gAxE(�$Ґ?r�#|ȑ��p����
��w�c�	]hr�h���R�t��iG:ADDDDDDDDD�J��C�H� ��s�>�Xk�\2���'��@lX�8hF�1�&���B���V;��36���(Y����+��g`�_����Қ����.·����Mr�4�կ�v�'��1�0F�^�Y*2�u��Q��r'{�ӆ�h�N�;�.����!'"""""""""ҙJDƊ,�db��8Y�a�G�}�{�.�;ь�N�:�8ഁ������%0�sQ:裡��7��iI�@����Bt�'�������E '�|Ly�,r1Bd|ty��R	�P�	t������N#���xשsgu """""""""� L'�0�P�Y�0Ad���D3 0X��˩(8��Ztb�݈�N�8u�㴂���4'D�����p���,.�������p��-�;�g��8���8��/�p��c�|��Bc�{���Nޱk�ҩ�v�DDDDDDDDDD^P(�-b����3�<@]�b�Q��(r��fqxǩ�j��=�,�}%"""=�iplu�_C��?,Z�	҆>���sϑ+��3+�(��s� ̑;�CDt�bD&�9���KT��T�%�{�)ӈ����������K��1�,1ӌ<��*ַA"�!���f'�UN^�+�p�DDD:�������â�@Z�~����LYy��@b�SS��*
ܝ�� ����a"׊����^�9� ^r*��X """""""""J5����k#�.%�H��D1Γ��8xѮ�3�T�DDD�5[����n��y��� ��@�r$0\�/�X�\_fu��H��(1K�Yg,�;�Xb�� """""""""��6a�1��KV'�B��E�,��[N�ʰ�i iD�;*�t�l �+���y7��ȼ�0���}౉�Ð�k̑8G�d�4��!\����b�;�Kv%�{q���(���������(:��
c�{:y,��ɧ�B��+ćN[{�S"""�����M�c�^��^�y�7���yB�*J�ë�]c����`�)d8������<���T���N���������(l�R��0F�L��7�D~���&���=Xm3�@DD��3o�������� ��^��t�u�����}8[�{�9
�CSfF�����3EN��I{���A�FST'J}���n��p�D.~hNûF~o��n�DDD��q��:�̿��	�o��9��_��|XC�b�K,|��\�}�
x\mǹF1�v�9� ��T��[�q(٠�����7�����.4�2"""��_��s��5/� y�w��w"�S'����9�D�o��W��7��[k+S�DDDDDDDDD�,��)s.3�q��0�K_f�Y�@��ځv�����D<�%s���y�7��,��M<��Ռ�����v\'|H	�E.~��^�m��A��@DDDDDDDD��N���Y�B��KDJ�@�ms"�4����m�F�����2��'�d�5xñ4�����qL3����m���i�b�B!7�0[���&��lDDDDDDDDD)# 7��q�1�SD!�����6��TBg���1��a��MN{D?#]r�D�c��o�:j܅��R�ȗ��X<�B\��U�1ulK�/�c�I�q�B�c(>o�qw�)>F�,�֜�?�;�} �&��zd;ǉ��D��щ�Q$��F�J^�tc�I&�G%�g����%j|�P�L��1	�*Y�kި���c�3��lL|��s����;�Y���W�����y�ʦ�z'$��:Y￼Q��MT�O���T��TLH�$����ޗ,<L3q`bb���"p`rb�������w��wjb�Mot0y��z+&��7%�?#�	�^9��^U��ݗ��m��.�F���MK��9�U�����o�*KʎK��Z���S�^9�S�i����\-�������S���3#���.�}^����F���=3������q��G���D����I*�A�.�q�oN��q��m��6
���%�"ufE��v���CQ�"�~���`���A�̱4��=��W�2�e�G�b��|����W�Ly��ފvGϝ���pp��ͯ>+ӟu��|��q�y�W�x����Xe�?��4�@ŤļRa��=S��l��&�i�z�<�y����>�p�L�>{ds4�f�$T��=qpR�R�Q�	j"��ƉK���7�� |���5	�je�K<To�����4����>+�A��̈́5UTXef��&zf|�;�������R��9�^_'����ԫ�'?*��]�ء̑��n`����;k��#�_w|;DH*�1kq�}���}���qr��� ��8%A볪�Q�>wz�����*�=5A�6'="�i<2�9r}��
�8-1'�x�^��+���%f|Us�CA�5����'_����zuu�1_4ǻ3�R��cؓE�6b����[/�� "�!���;y�,�v6���{۪��lf�XFecl��5b[�7��x�Y���@�Ӱh��1ql��w_ 3�R�?0��3	Pb�c�(��|���6�@nv���g�����D4�ˀiO=W��l7P�&p�~3��Nx�%��bqo��9^_e��*0�&��wƓ_�zm���{�ka������Eܛ�^焔�+(�׈{ح���g�9!�Vv�s�n��e�'Δ�i�Juv������9!cVu���87���QԈ�{Cn��Dܛ����3�ŭw��7�M��p��p�����r���n{-�2���2��ͬ�q��S�2bM��*��z-�2����^Q���Hs_Q�ߑ�Й�-s�j�Z8GQ��xO�_�p�����s�)#޷�P���>7�;\�"��7?|������.2�[���ڊ��*Q�i̅��I�to���X۰�����O��)�to�?q%껚?v�kG���&^��||��caM�V����b�b�u��ϝ�S\0xV�?����uXU���^�����rp�ٸJ.�g�����;p��g�Ӎ����H
5jb(<��_p&>�|#�����tN6`?)o��ᦈ<�М�\����"��N����Xg7@G�lL��\�7$�M`U�4O��&p�n9��z��87����I5��#nMQ���6�-���XO�szPM`Ǌߙ�^�Ļ	��z��j8GIDSԫ�����J�Ό�j8'$�M`��sB���j8Gq���~T��Qo�������P�n�pN��׃a����vį)�α<�>+C�;��ka�9qZ�=F
��z�Ƨ^��sB�lP�_�ϋ_�^�)�p񮷿��}S0U��G|�Os�x��""�����U�2�+o�EY[5l�vgJ(N��)�����?h85ӃZ&���>�������p����?�����n�:�O��{��������ǅ�OƼWn�5������ n��
�q�G�%��4��l(��Y��6홢��MB z'�u�#W����q7��e�:��Ɣm�����WX�z��.����=��z�u&pw�A�׫��j*�]��vP��a$�����؛�^�(�<��a%�M`�U��vg
z&��p��6��tf���HJ<ό��xI9���G1���pNH<��^���3c��	�WS�k��:�!뻟s�Ήm|�F
��{�s���4dc�����c[��8SPo�lr�둅ġ^��sz���4���0�z=8SPo�UoS3��iN�0�����jL�`�� ��^k+����S׌<�`�ᕪ��m�����M��g|�P|r�||z���>����8����iy8�`n��	�����\��k7��=/}�����x`�
<��%�Y�ɝB'�=3�������Kp��[���K1u��䍟��U�����X��Z`��M�蔻^���)�n5'"_�Uo�1�E}��zf�N�ƣ)Z����?��x�	\�����a��Qk�uX�pNH�M�A�d��5�7�3�u	�(�h��	�Ǚ�*�3�Y����X�H=�zf�.��^+�&�᜞bm����m�z�FY�᜞bm����i����ʇ�G9��+��W��F��%�2p��i�Y���Ԩw����YY�E���s�=�)�����.��^M�9!����&�����D��yF1�?n@CDDt�����X�V��^�O��r9�m��q�����8�I�v;Z�9�o�x���=��4�p���?hx��[�������W`PA��V�����ny�;˃��4��a����p��~�{���Xw���#�c��S���c1�����Nx��u6&��ߛ��%"n��Fɫ�v��h�������^��2=r�&�^�k}��	\�YI��	��ѳ�h��-�mX�pNH�g��	���X]f
:�{fl����:�szRM`���#�w���F��-���M�M��}G��-�mS��<Ԯޢ�j���0��Y�0R�j�N��.���-�R�����,�Y�Ի+�z��
#��9���»WGX�&3.�z��4���Ӑ	o���b�(�O|���C�:�$x���_M���x��0CO���Ft�'*��n�V�.��1Y�?������UXB]�B��SrGaU�z�O��t��X�J9�_�O���Y�i��@��9s,�6���E�L� �dy3�0��Wj���#�4�������o��6���`�kz֫D:=��ᜐH����sB"m���)�3�u��iX�pNO��	�c8'����4�U8g����(�鑭�ό�5�����sB"m��	���X]�9!�6Eu��1�I�_f��ԛ�]�5Eu�(c�G���9�˭��.����Ta�OZ)So;Q����H��|=E�L~fN�Y������v��=c�7طotb�zį.�c��^ˏ~���I���l y����o�d'�g�{ݫ�e�p�o�9x�I��!� 9�����S�w"z韽�t�n���X�Fs4�����|����/���.��	<J�:&����p�>���ޑ�����N��s8��p���4���v�HIPo�M`��H!�6�U��5[��e�{&��a��	���癱*�T���:3��'-|�G�P�pNH�g���I5�g.s�l��:s���=3V�pNȀT�w_��jF
q��aԫ{8'D�{��wM*ջT�{���(��:Μӛ�J��A����z���"�Ϝ�0�GM���cs:�\�6x/��-iR�qܥ��:Pa��"8򹘾�`B�gPW�����&?�>?�����g؏��V��msS�;����'aV�D�]�9!?Gͨ0s@�{���uQ=��ݭa5SĦ�=H2`���/��p�4�Λ���h���H|B.�mj������0�{������&��7-�^�<�������	�,a%�鑓�^��3c�%��W8Y�9!}�	<�]Y��$���&p��sB�:8Y�9!}��,ᜐ�>����	�	�,ᜐ����Ϝs��ΌM�pN����#�o��sB�j'c�Gk�&KX%$G�;k���	�m��ד��JYo�Q�M�pNHv-p���D���>S������M9��o�y�	O��Y�Ю�n�����gz�0Caa!|>o΢B�gV�0\�o,;I^ )!���Y���5���1�^,+{ϗ��ת�a{������C�#z�6 3����t��.=�-K"�=���qӘ��������kBt�]x�gq�{A	��W��S3�;�?���\jŧ�� =��4�Ѕg�����������HM`�HI�zU�|��XS�d��a$��ɐ#M��lᜐ#5��-�r�&��l�~'���#M�lᜐ#5��-�r�&p��sB��N�z{i'[8'�Hg�|���=�$<�	�lᜐ#��l��)�K8��9!n����'���W5Eg����k�7��9!Y�N~x�vjכdᜐ�:�<���k�=v9�e������6Jd�Ǿ�� �:P3i|ט�Y�ak����̄eYhnn�1�@^3�=��u�@DG�������p��K��8,1�]���f��^�����#{_BcW�QkL�`�3�^��aw�G�=[CmgSD���TşO�6
9��ܶ������i�/o\J��Zg}_��Xa�Q�[�q �|��Ztb�]�caҋ�{vD���vxx«�{�.Y�Ua�a�w���鑓5�rxX5���M�zo'k8'��頓5�rxS4Y�9!����ᜐÛ���	QM��e�o��}�q�8Y~&p���BTӬgS4�f�9��g�&k8'��h��sB��Sv��u�m ��Ny�>�M�pN�j����P�IV	9�^uY��$o�Mr��Po]�s�M���wx��-�雊l��r�Q����X[�����9���/1M3��\RU������nYs��}�{1�|��Y����q�S���i��/�{/���z��것��Vu��B����3i�_-�Ç����v��@��q��ECNvoߺ���a�.$/q�{5�yq(a��]:�|Z}3��(��/c2̤}ۖ�9f���m�lw�w�u�r˝zR��^oBM�<�A���o�����y�g�${��3�[ ��9!�3��I�		5�����W5	� ��'�3�UM�ڡ�g;'��������M���m?D�#%��t��*�8�.�^�	\9&����>d�b0jM
���[9Q���$;U�i&�����M��	FJ��6Eb�t��H�z�e���]�{����S��L�M��m��GQ6#��}�:��~�����TB:H?�Q�b�]ݨPÐ!C����:\�Rπ.n�)2/V��.~Ç�
'cV�D�x<���,_:������ʕ?ē�W��ۚ�c�?o�������s���7ồ����A��͟��{�>�����_m^�{�>��g�7x��p�3���H\���!�������ZnSS��М�/�E����ou������jI�z+�R��T ��9!jls*���U�j�T%�;D5	3�2T8#����Z���f6���J��:֗j���و�Rg}VM����u�X�59����>���:�sz3��GG�ֆ���pn�oYIwم#	��^��7�(;�@��1DH_�5�b�ӊ��Z�D����@ Џ	�>ttt��k'5��*��NN8���N�V�,�Z��]~�e)�}�ɴ�Ւ+�~3�x���#�����},�W�-\7r.���x�j�Q��;�S?�޾�3���A�@[��卟�"1���y���WE��jF���MF�@z(��=9��\��uވ��������t������ ����m�$|%�.�DD���࿃T�f�炫�h�"��7����Ä��`�,��������a'"�쁷�@�2w�	G4|y���Ϲ����|�{	r$=��a��?��啠�KL�����\%�3�'���9��6G�/�.Q��.�p�1�����M�7���3k��:���Y�7j6���>J}g�;C4�/�4(�3Fh8�^s��ج!G����^�{O��{��=/���:�!�D6,�6��[����a�� pv��~���U�0PrYd��{v=�w�ADDDDDDDDD���cNrgå�1Nd�'�om������l����a�ޗ�x_S8�h�{{Mݖ������l��1&d��1n}>�w��ܟ���U|���`9)��"����~�W�4��h�5W��-��C�d�Ԉ~ǜ�/�E#�@DDDDDDDDD����/雌.7��]�o9� ""��l�˕`��aԹ��Ƈp���m���aHz�{��}���9ٝ}�h3 �P�u#纷;�`T�3(_)������{�]��O�!���U��͟!�XHa��ߑ�������.��Ü�@ɩP�����?	n %�|�s����N��on�A�Óǈ�tpǆ0g�q��gaŜ�p�ߺ!5s��n���>���ۛ��o�^������o������ط���z��7w�9�*������+������~��%�|.�LǸ�!�~乘W<�����=XR��!��r���[�0æ���kS)��;�e�v�V���I�q>�����z�7�4�h�u���D!(��)�p�Q�U�>�㴀��߈�cuv����v:-=̈́��zU��f/K��e��c��H�qy�����oכ��9j�Z�Ϧ\��S��s��+kU�t<�P�_֛�z�������_R�ހ|�M���7����l����z�z����ǃ۫T���|p�1���8��_Y�AD��4M��/���M��J�W���k��������k��5����Z���ø��n�@Q�7\��h�:z}�I9#���>�.*$���n#2����7j6�����iL�`�3ﾣ������+����Ӆ�Ovg��>+�����s�;�Ɵw>��'D&�P�����&~[�G�-w�@��ȅ��cA���f	�:hv�x#8k�tuu #=��X��ؽ����[�Hf��VocSv�zk��i'7��{���]���1}8`��9��:M-�޽�;m�|U�Bz���$�w��;m(�t�>�j}V�+��\yܔa���Ƿ�����O�6y|������;�֠���©�� �b_U��=�����<m�`�v����v��U������p�S�>��;Y֛��b]�;�so��띢�Mr|c��`[G��Ԡ��6y� de��J����]��z'���,�������z��>��-Bn�s�A�zǏ)B~�_�&��8��|=����j��U���4Y��Xt��y��g�ނ�ܧ��q:��ؾ�����%s<�E�6��ؘg�e�kl��#��!�CWW,�r���D|��td���ޫێ�O�����@����v6�3*�l�b�����}\<�\8�d�ʟ���<w�I]b�;���n]��{q��6�2�i�;�ך� ���Ĳ��z���
[�1z�a�ԌB_F��_b��w��=[3�Y���j��9s,�/5�*�eEn4�࿭�Ё�ob���zskԡ�ܯ����'�4Aֻ9�3Ts���NM����1+��u�P�[Q��8jP�ߓgN�i|U�J�+�_�z��:s�߭Q7�Ts�B�+4��0�1k^{cKԡ���Nm�g�8�xm��ǷY���Z�k����UYo��+���W^��ZP��'�Wg�zc�P�:l��!���c[�Us�J�x�^���}�8��jK��)��b}��9�����[�n�w���V��#�Kb�b�W5���Wk��U��u��}�u�!T��+˕�sl�����}��cy��>�%����7�P�jv�=����z$�w����Wֻ�@��@�_r�i%x���Q�Ts�M�7��>m��w[ԡ���SVC�~�[�r|Wo�:Ԡ�ݽW�zC����"P���1���A'�=K�ڕP�2�0%�U5�q�k��3͝٠0-�T��asS��KP�;u[��wgv�Q�����Z����Ϡ��7�����P�5�ɏKAq�@��s|��|k��v���Z.2��y� �:᧷���4N?%�P�
3TV����0eL�4Ч�<o��%⦷fP�j�f_�{�)хTs_5M��=���B��_�Y���O��:�y�?f������0��	Q�8Ts�@e�V㫚�� e4!]�=+ʦw����5yo�ꍶ��6�+��7��J(̠��쓃3��	Q�T�a_y�;��ow�!�&w��{}��c��׫��6�C�}UoP���^jxE��6�Us�`��o�!�P�A�ki5��ߏ��>��g�9C���q��g��޾��A�q�B���i�T�a��Y�K�z�G�5�M`k��r�2���e�3_�4�����8n�)iXh�C�����;+��6���o��1�e v�T�y�#>�&>��
�bh�ߦ��r�9^��>ŕs5��~�g��+B��H����
tj���zU�!������P�!�&�����hB�澩���N����7���v��*=���G$���֭��Bg���n��Z���4�i�k&�z+����C��
�|�FjP�n5S��㫚��O�(���P�[7�3SL�(�ѳ����z#5�l��&�PCh�3��w��קc�BD��p�Ѳ^��>3�PCh�����G��f�M4�f�YV�Utr�9ÐJ=�0G`�]�Jhtm":��t�QX���G����,>oC��h�m�Q��"���؟a�u��PM�Sf�P��>/���\�i34�5���om�;x$�u��6SBT��ԓK�r�VYo�����6�CB3q����0.�74�W�^_�9�ˡ�>�*�p�)ܙ)��}���3�5����[S�^��>�49�o����{}�5�����7��d��m"����\Q���
5�3S�z�x�����=�{8�Ge�z6C�8Vn	o|�h�,nSt�Jr�Ԩw�iݡ���l2ݟ�Cr}�è7���׫�ax#4ӊ�>�V��j����^7L�y�ݯ�[`Y}O����m} ?�#A�) ������@DDD^ ��5���A1����� ��H/�h���`����1Xe���({���GQaV��T�,�d5�(=Ï�E�}�k�ʫ�/8=M����4�
�$G�*�RT�w�Jy����PCAAVX����̰*��W�8����4���7�S�V#;�U���0,�O��Y�¯�
�|γP����_j(��7Y�-p�'������/����W=��$X�U�?�}�e��K�z�@~>��M2l�B�F8��]d�@��8EE1;G��;��8� q{�!ݺ0�"���F1��LPj&2p�1/ٕ """"""""�� ��͈�LIFE��7F����~lq�O����/�G�mbJϙ�E/o�$�@�c\�	a>�.EfghD6ٍ�
tTעsw�վ��孰�K�N�\��	c@�����"0j�H+�b�9�x>�0�`��+v,�5�ѱv�9i��da
�Q�Y��hm�v:�j��M���Dgm��!��n9�����!�9�i�D���FN�0d ٩�������i�EuG��܋M�Do�r��]����-/]h��E���c�X�!Ymq������ۜ����{$��-�{>������k���|�-���%%Fα~=K��"��:�BDDDDDDDDD�<�q�Q�dU�tb�]]�-/�m�>R���X�J�����c��WO�W�夓���w�U�?��#?�6����<�1.1�-� �O�cD�mWɝ�dӌ ^VT���?�a����v�EK� ����xxn񩁢o����6�e'��W�h """"""""��%�`"����߰k:�85�x�i�q�§ދ�A-߹��Z��i%�iמ*��y�9p�H��T�u�X���
�gZsg�t^�h E-���m�i�u��q"ɢ]X,߱¨�Ʈ�O=��t�K����饗_q�(�{�Q<F�������"�>�������������K�aHA�xݮi~ɪ��[��3,Zݖ�t��[����ч�\v�<���qFvRL\i���v�1�pΖ�DZ�l�p�0����	!گ��{�|�34�3"��˓d'ۂ�vE����O�X��s���w/x���xn٥\��\lh&�i�C��b�����������/g1 INvZo7s�ݵ�f�q�����ׯ��80���KF^�|�Js����z�Q��Y�ІȮ�|��Aض��y���H�@�b�\~��sg���@��s|��)���E '���P�9��&{�������y%x�~����~��ߟ8l}Q����_'�h�4�,�;�م�`��	��޽�Q��u�?�ߣ}�3{N����+�����bP4��x��]�������a�4���
S�444����aF�uP���������9q~���>}���7�����}&���ʚ����]v���n^��
�|kے����(~�<��Hh�쓿�<�Fl��DDDDDDDDDԻ����mu������|c��{��=������ƌ��?�sNv�K��4+*�PYY��Ϸ���}izo'""�pN�_���Wڑ|���xM�}2�=2Ǚ���~��oj��ܵ���]�zq�۷p��ߔ�:r�3��O���k���|�������ݗ9:���L���Bg�n�NX�e�z[t������+��uVfZZ[����Ԫ���	�tYaԛ����f謪��|��aԛ���f�뭑��۫���U���]oMM�|�"��o^n�������w|�Y��r�����ŭ5�zs��������
����\445Bgu�m��l�a�� �mԼ���VY�V�j|�����A��vX�s��<�>�}ٽ��6�VXG
�����w��M���H>�x�e��ij����U�-* ����Yd�森�:ki��h{���<�� ����2uMh|�؋vE��;��U~��5�Z��$0��tѭ�1��|�����d���"{=��uv��Dv'�΂8t�5�C��!�d�&�w���/�ADD$_���O�7�A��ǫ��1��#�g� r0��Q3�����Њ�� /[��mV�۰��}�7拹^�M��ǈ,�t��4U�����g�u��#���2��y�����~s��73����n܋�V=�(UV6�Y�oA�㛟��-Ӷ魚����;`֮ߋfMC����&��������fw]]c��+U����ܢgST5��j#x�f`�|�6i:�ղ���-��u���ؤ����ouu=
"�w��M`���������VT�ET�m������ނ���t�W5���#�7C�+�m��������[��MѦ�v��_������[jt����UG8��uL��9�z7n5P[�gӻ��{˪�~����$ǷF��[�ު���(��u|U�a��*��
o}V�/������5� ����������z�]���E�w�<r���	���D#W˩��:ڿ�E4��ò{8�sO9\�݄�.���ɃDD�!�#	B��q~�m�}2�����L�'�G�p��펗<�Chb���d-���f�r�~���l�彆�
3�fw �u�L��{�jث]�!���#�w��/��mf���&444#--�zC�z�c��2��lw���M��+��:B�&��ܯmDzZ�/{����2ġꭩm�����2��6�k"�W>���ն^�>����Ëi���i73�
3TV�"#=�}U��Iðn��]�#�܏�^hjP�}���̈��i��Ͳ�F���n���z��^���1Ԡ�=��
Y�PY��_�*�p�Y��SJT��{:��ee5�ʌ����|��׫	���eeU��@���=�C�q�fw4�N�볎MoU��U�Ί��I%Cd�B�zUsϞ���u|Ca�H�U&�-vgܩ���j��� Os�G�����{*.Z�|p��w٥g~�.ye�1 ����q�m=>��p��Ρ3���*���$"":����9.�&�����c48S½䄛6�4���;��B}�!//\|{ڒ2n���N�oxx������^M�!�4�jx�4���Ua�Ʀ��!*�0c�H7ġK��m��Efq�����!].�Ms?�m�O��L�ڦG�0��~H��6���X�aZ����~���PCk�M��(�!j{uܔ���m�zl�Us��2��~H�G[��s�Gg�G����hk�c}�3�D_���G{��F����h�ң魚��֫B�5��i�!�g���C�z�����B�86ۨ����M�!�g���R�&����S��h��a��
M�WфBz6�˫��h��J��M[�W��D�����JE����,MO{�޷���wOƂ5]�Ȧ��^���W��B����"[�����K��N�>d�d���BCS3�WԹ�Qt�1`��w����֡Ƿ�����1�3��Q�刌�_z���!�qZ.���g�|ii��ɞϟe����>]���YΠp�v�tK���]�s�߃��_��iK?5�s���}�gZ�a��p�ΔydG����u>|:;��g���hj���FYouM�f���!hj�+oyc����U�MQ��N)�wZ�������3�**�b�qC������hjjw�šަ&u������܁��:7|[����*Ƿ������ឩ���z��p���z�Թ�X�(��-�e���C--�(�W��X��!h]g��5/km�BYY�V�i|���mQ�z;���މ�eU�H��X�G�+x��6YjY�?�z'�)F����������Y5C3�c�	r���n����Mﶎ.��fƫ^�7��;�ع�B���,����6�=���hb׮ʘ��у�&��^o�w��ݾ����Vo1��,�/���=�}-�z����;*ܰY,��3�Tx;��zǏ(��AO�{�Yݼ`(�}��q�^a��u�<�����^�yc�ӃE�>Z�SD����0�C�Ý�A�w�`����u_�P�b"���@D	t�\J�q�a�"}d�\���@ �fg��V�i�kz�Bt����h8�Qg��־w�\��OCsO.x����n�z�1l4r���L�ή�傔����%U|������T�w��*�m,w�T���
wI�7U�K�X���]R��-�*6ʱݘB�yk�����۫�%Ul�^�.�b�jwI[wV�K�ؾ��]RE�ջkO����d�w�HwO����������ro����j�#�f-��{_1K~�hF��|<j�ѱ�BYYY��""�>˲��ڊ���s���Gyd����CA5�8BBͺp��/�kj	��c�-�������9:����N�s�Z��^�P�V��#���$� �8I�h?a�u;Y�u�X�Ӆ������H�._��]Ö~��k̑���)"Y��Հ�����|1\������i����8��ӟ�t�����߳����8�1�kP�!++k㑾e��)F�S����]ԡ�y�s�E�W=��y>#P�hI�ӏ�qN���B��qr��A��� """""""""5��^'�-��>���G�D����y%"��D#?P�"�n�b��|3���� �DDzJKKs�ekll�s�^FF��kQ������s��vӺx>x�鷯)}I��+��K>��'|#/�Tf���&'ir%DDDDDDDDDQ�:�^o�u�Kj�}�f��K��8��]��ɥ'��<������L?�$=_AT�òl���""�Sn��@�'?��G�������u���N�F���Y��z$�gs�Mon��b�CS�4����������a"y���	�/��fܼ�I��?6y��k.3���4��9��mA{{|��_��iGb��� oSg����k.�p222>}��D{ɉ�p/91Y���+N�U��4#IU��`˫K��'S�w'4����P""""""""�T7Y�@��+7�t�#���^�W���)i���x�Ȇ��ό��	�nEZF��x����pDJƍy�m�hkkSӈ����aY����sT�!33���g�z��hghH��%��h���[�X7�HrO�-?�m4~w��͂Ǎ�;�DDDDDDDDD��qV5;�;N���]�x��K�z�9l<N�F�Llw�9�od�9���,�@ �W ""oS�쎎8��П�.3���y��7��b_��.� @r�����V�㎻���Fk�k���g��{<n�\Ͳ�*�NKEDDDDDDDD�m����I�UV���<�*R�*��Ƴ������]Z���h������.DDD>�/�����={��|�w�՛����p.91z�d�uZ�%u�~���f��;o`�F��(-�C�?�E&�;� """"""""Jec49ֺѮ�R��E�|oٗ6�#����Fk���3���DDD�\�=iii�r�kSS�n�馎H�?��p����N�jܼ&u⁲�KO~{��y<n��b����������RZ� [x��$�6�����D
ل�{��Ǎ22��O���"""қi�*�������I./�����O}�2��L�^�`��SW�������M�������B+�`"""""""""J�����z��e�q��������Q�w��-�=Fd��aC��DDD9�4+���~iY�q��|>_�"(��$�O�ogee徛o�9�	$6Ѐx�N��s��?����G�����:G!+ +i """"""""Je�����i���;�˾�v��:6H�C���{�Q��A���'}�����RWx?lذ��<���x饗��/��@��h���)j�ղm�������!""""""""J�bή/w��g>�O��
�?#?x:���|�Q�N�K1�q��=?W]]���������Hݧ��Y~�C<~��
��O�w�;)�����S���@C!��%R��Yw9��q��R�r![͖?t:��*4�eE"�DDD�`0����N��~b����@���*'�y���-�HQUAY��o�����!""""""""�D�Eb�C:�E�Zu������}����T9�X+�8ADDDq�8�߹HX�8�|po'R�� ��RwG�i���O;A'[�<* ף4�u %��DDDDDDDDD��44;�;Ha�vW���ay���#"""��%,Р��N{-���d핏�ڞ��x�z�V�t���������(�p����|)�]��OrT0��34��p�r�gZZ��'YQ��'�&���Є`R\��UO�`���������(U�y|&� l�x)�����lxX��ף��f�Z��***B  %���~�	%(��� �Vx���"Q��=~�O�c;kN�CRXP�Zx����h�kh���f~�u	�� 8M�.�7��a�Hq�m�z�0�_��p�������H;�k]�N455��'L>U~����DDD��Lx?�imHq��z}�|4Q
3���u	�B����G�Q_W����'�p`��>j*���@DDD�+a����?R��9,��A�|DDDDDDDDD��R�[��O��"���}�0���Z���eBa�ʚQ�KX�A�&t@YHq>����A'h """""""����FtL}�e� &D<�zM�ay�Y�]Vy��[�f ""J!	4tiЄ�9")�����LcA���DDDDDDDDD���Ft�0=~�1�|�����8�\�l���۲��{ ""��IX�����NE��@�˅���^�a""""""""�x����c>�N��&�r�=�����h��8���'""":\����"���5K��F����KDDDDDDDDD�Ҥ���.#8G~H�@C����@C#�@DDD���Za��l�M�zU���=�ѿ���]HA���W�e����:�z����������(�58]�z�<]�S�? E���@�(a�G�ir��x�ϺR��� ��z9<N��>����������I�Ft�8)�//ߞ^X�τۤ�L���ې��q�g33�PUՀ��vQ�KX�A�E'���@C��)h�u�+���q:@DDDDDDDD��j�Nx�p#}"RԦ���1z�H�\��ӱV�5M���8��'L�<n�"J.۶m�k����{��qdgg#''yyy���=�Z�����Q$4�P�t`��v0u0�f EA���r��������(�U��g���?��iw\z�H1�0��:a�V�`L��/��߉�9p�!_���DGc&�LD��"J�W��?��O7�����.�����{��BK���
=���EB�N�n���{�c�w�U�ڎ�үMjd�����iÈ�������(�U8z#�;�e����a"�Tx\�\��c����� ��P^^��0C8����HL�tC���
C���w%v���2 ��t�)o^����#�h��Y#""""""""J]N�.� �w>���í�\x\9O#"{��7#3�˲,444�ˑ�|���P���gff�����v;-��(�u)R�H'�"h�h�e"""""""""J��M"'��sc6��.���/�|�U��R����.߾�n�ץ�����#Z���@Q���ʎ������s�#Q�����0`���C�ڎQ�%tx�&���"#��K�z��ܻ)�G˾�`����?���h%�.�Ӎ<x]�����p.R���=�Ұ�@���c���(u��z��B555�r$�@���Ch����=��Qdhh@jщx�ə/�~-?�D�����@��)w�� """"""""Ju;т��~�a��=�O|g�mW�r?���9������G;΄KD�h������r�#	]�"??���s��*,,DZZ���>G�6�'�x�X#{�O~s��߽I�˾q��u4��i�ce��A�a
�
�'o^�$�����b�	肍��	��<L��'�^�"z(((p�jQ�C�=p�J%	4lp�4��8����9I�@��M�wADDDDDDDDDz+�"r.�{�w�~s��w I-/���� -N���4�6���*���zر���Ҍ�7���Ԭ~���)၆����6���F������>����gf7��m�����RQP�>
������DPPDQ�G<@��C��Z(�һM��>w�lvg��tb����l���~޼��n6��ff7��������W��[
��CW|o��=���@���l���� �7'�5���;�.����g��*1:��l4��������^dz��B�Mm!��H��H��ڨ���ð�H��d�����Ú574�C����3���A!D��SN�L�-F�����Z��<��~�����Odj)j�| �8FD�Ʀ��pB��߻�$� ��d�}Y��4h��z�����X�M�
򐚺���u� x�i��_�r������~��ga�Cu{�l��P#� 晹���W�pٚ��G���oݰ@�YED`bGh "������^5��@KK�����x��g��0T�!++D�i�b�р>5b�������ŷ�����[��W��ܥP�z�=dde� 5A����0::#p���T��Ĥ�::�Vͬ�M�=w�"���f�)HKML�*����U�/!��F��[�����='S����uE��������ׯ
�7��M��M��9��M����l�]]ڂ]p�t�ތի��e����mc����f՛��z�a���_y�^9�
�<�"WKIi�w����[�f��?tE�W_~�,d)3
���lA �~rD"�o&�P���gڴi������/755��`�733�>�T�4���e��@��@�[f.��d����[�֫W��󇠰�?x����@1��3�8����
uX�GvP��1���ftt��Y>���މ����W�z#V�#]����(�lr�˦Y; !�ޑ�8H��UM���Y>��9⦊*����S����zG�~��;PV��zW,�]#m���Z����������Ȉ�os��~+]_EH�#^�-��(���jK#5�D���r�u��]Plm˦U����ͪ����.�7	���M��qZ��W����y�܉������H�����]`�ߜLR�#�7н=�����s&bB����C�W���Y���M�_7F�8��.�(���3��i�k#�9J�{��]�=K��S��G�=�]�W��zg������ޑ�_��� \ͮw�U琵=7���r�����T-���e������s���<t�d���4�R�7g��
������t��r�Jlذ�&	=����KEEŀ����v��Y
=�B4�1	4�1��1;1YK�*R4]����o}��_~�-/CA�z��3��w?t�v��CY)�sT���q������mq7������fѐz�=r^���A�M-jԫ[�s�B�����ׯ4����zk�	G/�K�n�;� ��+U�"�$����ׯԫBxT�=^֯l�q6�%�P�(i[^�V����z��w�[�u�jlϲ�p���os[j뛠�-��_� /��-��+����F@�i�V� k_�w�A��5�j�+��qV��X��j��o��~5�t��qG[���w�A꭪��U`ZQ9��c�[�wgܡ	3TK����gyɭ:z>^]�3�& �^�*�~1�z%�PYӠ�'U��o�A���U�jlϖ㎲^�o�;���z��U�����j��~E�J�v�~�58��2��*k{~�ڞ�5tt����z�4�q�6*Y��}��W�v�9�|
z��eU�ߛ�efC1o���(yM�>|0�}�]�7��a466��`����Lg�{�	;���!%e�gǐ��$�`Z��b��m:T��o�/���?�ݣ�x��7B!�{컇�}ϧk�ERך5pi���3��4�uE>���tl|�i�J��B1��29���BN�[W�^��OX_�A�z��9�z��_�ج�뷻����vs_�z�5�Hu�I�~��_[�]��1Z)z��Eq��0�J����]g��3H�
m�Row�!����ܷvYTY����j��~U����jp���W�����x��Ns_֯�A'�^EV�M^��Z�__����/���
,����٠c�;�{�Ns�ޞZ��d�����_C��g���3������p���F���
4��Z�W~���W������>so[ݻ3��"(f�D���EbTS�-��%R�|��+���&��p�Q�#%E�)�hp��~::::�m�6Pr���Dmm��&##�Ѓ�UB�UF� o�5��Q�st�")�>S{�W����s�P�m�|礉a��Y�_ɘ��Z�Q<�'̠)5FF�xB�H*�O�A��#�PC���T�Rs�O���@�zc5H���!y�o��b�	5��֫Y���чT38�iz�3�&�P����)�=Ǿ~{�����߻�����n��#A��1�л��"�;���}u�~c����Q��{�|�fիGYow��ε�n1[P�L�:�N��o�6��=|լ����A<u}A}0��L=k&��K��F���
����W3l�^��+?�@�GH��/�ƍ��o���
���(g4vdz"Y����OVV�r�x�=�8E�Z�,а�lC�فbM�m����������o�kg��'�د���/�4�~���J~�.3����԰4�� ��u;�ְv�U38zB�o�p��ʎ���n������ۥ�a�ߠx��6qܱ�M�h�Um�������.��׬��pΪ�v��X�Z��hF���k���pN��%y��\�Ф��g�;��뷺�Q��+�{���t@9�ݯp����+{�FQ���nGw�2��vks�b�֨_��?�����T�6�_�1���0�8]��F�ׯ4	_�>/Q��]Q���z_��5����Z�ׯ8��yv(Ɉb{�a�U�W��rO�z��`$��4Tn�;b�W�±Gw��ᎇSZQ���gw�Q�s<yLB�Ko{誉�
2�9��\6�����5C��S��<(�eS�@�l-'�*܈�ξ��q��[K��y�Z�r���B!477���mmmhii���u�����vJ.�@�^*++��lg���z�������@��h?kT�Ӿ�PQ����Y��#�>��+c͚57��"/�x�����]��K4��a}Ƭ���S�(,�����r��1�PCa~����J�ԛo�;���Ҁ�p��:,	qDS��B��~��3�:0�z��2�:�Z^�I�� Oޯ�ߞ�*�<�7�ڞ�	fx��	QH/���l}���^����®7�ڿ�%��W>�E����R�摰띐�Y��P�]o�l�IT��~�Y�ٞ'D�=Wz�l�d�777�����;��QL��B�OUJ����K�e��u�/>�w�e~��U�OC��Z��cVo5[�)'�f}����@]cK��[��f J����4i��E�z/��������m���z?��"??��A���<;� a�]�k����T1�;dOո�7��\%(0�gV�����C�}�s��]��_��{C�/�r�@aax6�"�(�F�f3�j��)ZfQ�+��w�^������p�g�i�N��s��S��'$���� SUHsY��8�����A�r[$���(98�[F����̴�N��	;8��cLu��[f��
��"dL�h�;�}�ۏ�
?}�YW��ǿ�Ǯ�,�
ܞ��^��t�_oX�F#��#""""""""�4����4�,͟�e�o���|;��������g��o�hY�P\;"x٨�W��i`;A���2��4��m~q������`*���:CC�!�3*p�O�@��Y[�l-��V��掇������N9��X<��\��5��P���B=7��[%""""""""/u��o.& ���g���;�?|�s���_>s�;��yM�����k.��ϊ�1�%<kT��S��(2̀,�MuM𡩩ɞހ�W4�	�8�Z|pnOfchx�hB��l-^����[�Um�֯���U��F�N=�{�F㹞z�������6j�'� +��l�F�	DDDDDDDDD4�"��Q�O��2�\d}4�7����_�1So�����7ܐ�S`ej�=��/����}k*�&C�g0�H�^���U�g��D|�fv ���UFvp��A�m��d:�
E�����b	�"��Lm!۠|��14��e�ҷ^��\-�Rƥz���B����{O=�F�O>��e{Á�ӡ�4�s�lxуF)���������(z�G*�F��Tu�ed�Y�Z�,;$�v���~t��uW(d��f�q�W�ܣ?**3�w�:���gjY�����Y�Jt�L�DKK 9�}n���@SS �M�24Q�d�i4�l��C0<`���#>�u����B�jkk�e ���8���h����14��|Z���Z�F�����ϴ�\�=����z?��S�)o�M4u��7����TMk�N���kȫ�B�>����Z�2�@�l��Y��l�Z��FDDDDDDDD�&t��
��S�E�H���R/���})Z䮇���	cc
�����u��34�u���3n����y���覙݆Вj�kL���2���x2��MN&| �^ ��Zk��=�a�iغ�DD^ ��h��3�e�����*�{�X�z5N:�$x͸�֎�}�>|ݷ ^���dd#�����y�Mv��]]��\m���e�f�Y�@YE�@����-D�7V""""""""�X�ه��"��/K�e�eYΗ�"�KN� O=�Ct��L�i�F�X�hv�׍z�0��Y�B����J��ξ��BKKV2���ј�h ~�?��Y�[֮]���|z��q	4�g�j�)����U�v{�"""""""""�]Bx¨�Y�4P���f�W�O�o/DD�X��C��ttxc*�d���b���HMM�W�[�!���*�bP�����6:�޲��|�c���9�9hmS;ᶯ4�zs�z[T��Z��R�6||?7'-�-PYYE#Ru_T�-N��mV��r�^��Z�ï�	9�z�����&�DYo~^������*�^�ژ���-ȟ`ի�����o��w�z&��I�z+�[�o���w��=7(�=WI���#-��;1?M��[���Z�66Beյ-��U4�N�X�������~y{և��9Y�mT��ںVk�X����Ʌ�����j�ۢ�wR�u��o}C ~-�z�_��VocS>M>�_���Q]����1�[l�[�z��֮�]�S&���*��(�)���:n�{i��d�a� Q�$� g��2�h�r{gg'h���۷o�C^1�{�/�8C��EZ.(�|`6c��և���FDB!deF�j:h�tl�Z�lӻ�����]�x���wuF_��ix+�m�U4!�ف�����\�z��o�ڡʎr�._<u�j6�+�Z�숺�e���r�Oͦ�4���vk{��ީز]S��-��`0�z�.��ݡ��I�&��hX�st�WK��y��=�+�=Ks��ͪ7���d�k�j�_��5�z�c�N�^E����mi���"l�e��RoSS+r�Ң���j�[_@c�Uovt�wѼ��(�5�6������b��h�-����jӻΪ���%��+��^	�ԩYoSs55��͎��j��I0�^E��Rouu�Ι�Z���5�M���;{����V��F3��"���7�|B����=P]VV22⟒Y�'"��Kd𡹹�P4����hH��n��?Z2MfF����ֽ���f���޸�8�}?9�#M�M[M�(6���:Cq��Bf��?�>R�4�7m���Y%�a����U1���bݞ�C�r�J�!"%%�z�.(���4+�=K�!�@jJl��EC��o��^k�~��Pn���V�����]�h��i�ǳ~��0�q�Դ�W��"k�ʍLa7�Z��ہօs�1�\�C�fwzZl;��m��LU�^	3�74�\��y���E��8$�P_���U3��4��c|���䯏�ޅs�C���4�3ңO:Ι�z�Rm��������;o�D��j�	3TU5X���~5w�D��Y�>o�3U�CFN�c�o����}�|$a""��@O�A�J�Ans�J�E�F"P|d�/�1ȶ�-�H'�A��I��Mu��vSt�4���m5j�'���jh��4�'���]�jU�7�0��w�!خH�q�*�O��!SS,_$!ͪW�&a<aGw��;�lW��O���]�T���*5��x��ɿŪ��J�&a<a�␑)ʪ�؞%����w����j�o�A�q�R�=RAa���#S�U���7����@���7�0�c���TY���䗐NY�Mo����)���	5��~�38���ԩ�#�0�CB�=�V�j讷>�zgB
�W�F�ak[�+���-%	2�#R
"""UȈ<�y?i��>4ꃄ � �e��P�q4��Ev�0=y�����!��Pg���V��L�|#Ed��B�7�0:�NE������ީE��k�Zݝ���MO@�ӊ
P_/��{�����t͞�x$�X�W�z�L��{s�7��F��+7kh���~�H�o>�d���^9�^a�;��o�<�@�e���܎�����9�Oʷ^�=�{nU��Ԫ7E���)�4���~�]o��߲���"ٞ�ׯ���[V׽~G��Z���Wmp�������a���t��Uc��~�_����`{W܏3� �z��_���mt&��B��Fٞ��nmaמj;�4�z'�X�W�~�]o[��=����L��}����cW�U����p܏3� g����G��z��N�z��!l�Q��T::㯷 ?Ͳ=�;$��z��P���z�uxU��*m"(9�ىN��CDD�##��2iҤ!������"�Ђ.�!�W����vk]����k����K��bպ��z֖�5��,��VN�v��K�ؾ��^�����׳v���K�H�zw[��N�z��m��d�l���6�K�()m��d����^�E��[Z�l/�"�����N��C��C�4�^4j��H���DDD�7����dOm��������^����筝�i�q�^ �׌z�5��9ADDDDDDDD4�dt�?�q�o!Ȼ��e�|LDDD��|صk>��������3f�@ZZRRR���|>ttt؁	;�R__o�$Ac�5�qKd��C>RA��h��k#�N�&""""""""OU8L����$������l�CDDD�]]]�"&O��ߏ��l{��MӠ��Ө�4z���Fee�~�����auF�w;Wd��v��_#���Ev�al�CDDDDDDDDD4�~e��-��4���˨�TDDD�D���D"=�eT��3gڋ���G]](1\h��<fT�L}�;4��w�����������D��ύm��ot�<��� ���P�#9�577�>��G� u�!�� ""5����k�l.��B� R߻F����������Ǝ��J�?�9 �IH���!/
�B�/�+�]�1�=E���>�8�W�0�ccn�V��C�)���ď#[�]lDDDDDDDDD4�d��Z6��'��%GWjlE��"""r7��JWD��-�ٿ��JWQ��#�ь�1}�P:�ځ�N�>̤hH	&G`$��]sZI!b�C�ӬzH
��-w��HkCR��o����$y�Zʻ25�'I��Uo(˪�%I굶��, �IA�og�f՛$�W���r5d6%G���~�s`Ջ� �}�Ո� �7`՛�$�ᙲ~�5d�'���В�^Y�� �I�Ԥ^ͪ7I֯SoM�����N�z���c�|��F�c���y�`W՟�=I5�o��7��T�z�D����PWZ[�1Mw⧐�"���]���Q]]J��V��>����e��M1��A駑��a�}g��K�8��a�7�éV��aX���Po$M�[���ʑ�D<�$�X���O���ת��M3	����{�qO-�4	�l�����$��ڞ����Ɔ�zs���#��M~��5~s���@Y�^��X������fv���N�qăV�u�W���st
un՛��z����y~��[�WY�z�Ih�����o���ιV��V�G<���=Ǫw2��&T&O���3��
o�+����qj��{п#(���z5��3����1,�|/�>~�_��W9OUx R�dbDZ���hn�̦���[���U4������Ձ��h���|Q�R��]xݬ��[[���{�	ܕa�x�����R����2J��f����'}�n�:a��z�ڏ�Ϫ�)9� �����y�Bk{����U����N�c��}C�g7��p�E��!����#{|�$�:'�"�}������v�f��}���=^���u�=���&�Αz󺯯�z=��	��w__omχ<A^erԻ�|����v8�\��Ͳ����&aO8����;g'W���v�=���s����'�^ê׀���������Ի��
�yx���w�5 ��G��-������´�[f~فd4!/���}���l�R��α���(Z)))��Qb���Hr��E�L����؋Ǎ�q�7�D�6�CVm��&�C��jX���S��զhW�f��U�]�>O��?�#�_��l���t�6��ףM��pNV�ui��=��α��MQ/�댜��o{����U�ǚ��#�X�W��2�ц|=����&p�p�c�G����9�6E��s�MQ���3rN2��+�㰛�ODPX�z��sR�g"��3Y�ձ�E^��_8Ǳ�4�<���4�;#�V�X+1�.�>~�_�N��z[d��D��,23�P]�w>�ֶv���������H	RL������F9��x�	ܑ�f0x�z�	ܕ�٣1�3��`ST��C�{���Z���Й���zx�	l��>�7��C�ޙ��sz�o{��N����3c��9����XS���9�m�d���9�x�):`8���M�^j���Ů�Y�vx�L��#��z	�86��Ò�L��Dx�p�c��V�z�ԻŪ��#(��&�`�ǖ���7��&G�cM��7�7���H�,�J�� �yߞ.����(�)hw{���8M�
r�G�r�.���&p{�U�E�zx�	,s�Ksa�z�qf�O/��h��Bx�pN�ۙ��O�=�;M�!�H�x�L�!�9�x�)���EY���#4r�@��2�ӋW��1�끦�p��WΌ.���JSt�p�c�Gu,���&mU��G
�ԻX3�o�ql��n�w��j�_�q$[�[?��˧oR���p��֓��9��ޱ��l�[p�	C.��l�w#��f�ADDD��
4���Ev�a\��'\�H)�h�+9M`��G�kx�Q}��@8�z���������n��M��9����*�Ӌ�M�x�]a��BU�o4�^ToG�q�><��sވ"��P�	m8ǡzxȑs�zxȑs����ц��7E��:߈a�~p���R�&5�pZ�!H�H���u�ۏ�ah�V��(�9�^��j�{j�m8Ǳs����wڻ��e8�!��Z3�Ss2�z��f=�o��ː��abO�n���3	%�T�)���D�_2���>�a���T9X���5>��W�	��}k��b+X�3c��[�q�_����U�6��W�&pG�U��7��>�f8�p�C�&pgNws0�zU9�p��n[e*Wo����M�x�U�	��9��zf��xA�&p�������U�	l�s>_��Q�	k8ǱӪ7�jb��^�ю�����zSԫw�i��c��.�50�-���hG��o�q>Dҭ���Z���[�X�d6�������`�a��m6⇑��i&z�	_��)>���(y(��zOd/j�|÷�*�â��0L�"�/5P�jMі������AWmx��"΍�^�Ό�o�Vq���7��&�R��̙��s�5���9Z��W�3�yV���׫X8�p�C�3cc9�?Ն��7��P��X	��Vq���7��P��ب���jM�XG���nKSt��s���jM�XG
��(ٿ20G�z��8Ԭw���Q�yS�z��8J�N�1���w�m6[pEx#n��@�������v��+u��#hi +��v)׃�(��y���!;y�f'��/e�x���m�~�l�jT93��H���<m���ȉ�W�3cZ�M���s���)�o�4��P�)�:٪����*��3�5ן�V �_�q��4���H�s�4��9�?U��#�8Ti��4�㰛�)��9G��#��>36�p}x�a$�*M�xG�����MѷTX�	�W�&p���{Dw���M�xG��Ϯ�������iɱ�p��t��F���g�#��Wvp���BY�IP�X�g���;�����ؑp�n���#����͈DP�ЄHd����3&�������)��f�a�l߷��('�)E;n�l�?���g�6N����:���#7Y�nL`�no7M��=3����	������M�D���9r_��όMx�.o'*��p����
�8��NT8�����HG
�ϮWwoS��#%��	vqS4Qa$�ۛ��
�8z�}՝M���&p��x�n[o^6���HG
����n�7Qa$G�r]~�_pg�#9�����s?����F�����o>NыA���َ��ZP_��܂Vh�MO��H$���vL�dff�����M�����v|3�W�a�64z�c�����0՟�ͭMѺ9��x��s뙱�U�[ό���c��?M�[����8��Nt8���&p��993>�͑��0�íM�Q�ץgƎf�nl�V�nm�&:��pkS4���[ό�4^�qkS4Q#����zG:��`��Nt�Q��z�Jq_8Q#�gכ�a�sW՛�p��z�������ٰ�ޟ5rNՋ��'�>o$E�c-�n�o3[�e�|����7�1m9i�D��FSFV��)���_�f�qx�ҧ�R��"��d�~������F�D��������kj����E���ČwMW�[�P�G�-rf��j��v����Ӱ��ѫ�n[��Y�c���հ���۞�	]ì��X����(ֻ�	,!W�;{t�H�#7����U�����4l:u��&�����K�a�{�(�{��=�h��.�z%����W�4�����qнy���vSTsO��y�UX�r�z�1o�;�m��a�Y�W������0���o�U�;�Y������wC�m��>{��Mѱ�?aW�?�I��ѫ�n[�W��㎿�m����Q�� M`X��EϹ���4:�+G���ڴ|��x�'jX�(�;�Z���q��^	�|}��Y�=���猤�w<<aTb��վ�(��A���Q�یz�1"""���@��9�1ʱ�l�5�%��)(b�����V�C��:F��d���� i�>R�O��IB%G!iHӻ���Y���%Y���K�(]��K��w�f-����P�lH���%Y�/��%Y�/�%y^��Kt{I��dI��+M~�џ$��]=?y֯4�eI5�4kI��[7O���g���-f�~_�������I��7�<oԀ���sgq����HDD�L<�~��7���ӾY8G��F�K2���>t�]�$��jG����;f�웇|����hį��6;AKM��EDDD�d�A�|owE���w]�[��Z(z�� ~نf���������(y�5j�ш�����z14�@�63�?{�Qe�0L�1M�7""�M$�i�ɳ��L�pyx#Nӧ�S�Y���J�م�{�y��`��m�h/�5��<�ӲA��c�b��Qbs%u��:@DD�@  J����G���G�r�h���PȜo���/�^�q�3�کa"""""""""��6����6>��3�9�C
��w�&���e�lG�'#0���p{(����y�-Ŧ���8Ihp�����ăF).�g�;�z�d�W�:�ރr�����������h(rLQFxѬ��T����ȸ�mf�5�a�� RKff样5��9��	�Qb$�^f��i��O���ga�>1�Fl�^6�p���]fADDDDDDDDD�3�"��w�g���pC��|#6l5[p�DDDD�")�}f7E����T�ꛂ����l��J��3F52�Pcv����������h$�S��o��}.���d��d��7�z�Ө�;F#���ԀP�9�}"�n���O��!�-�E�q���}�^�eZ.�d�ن'�J�h�ڡ"""""""""�Dꂁ�j<o-���8U��c�B�=4:�K~.R�'�*T������#���k:����߅@D�<4M�����H$���N444���������@ss3(qh�E�O��2O�Ƈ��X�M�d-*��5^6k��Q�=f DDDDDDDDDD�M��Qd��R�!m��'a��M�p�7~�l�K�Z���F`�����%--���HII��p�(�A����!���F{	�wK4b�ن]�6܉=���*��k���e��v��7�Y�mf�����������K��#f91��ǎ�&�H��!7:�JFb�`4�u�뭯!	��3�O�%�1�5|�S�^"""�K�	mmmv8A�J0����ZZZ�Ђa$�o>��0����-�i������ô|�����b-}\�}f6��x�Z$\o}@ """""""""r���ex�(C|8X��!Z�j�����q��a| �Y��m6`���������Ć:r��>!���(�d$'� �'� ���dzR1��v��2�����Z*i9��,�ֲ0W�FҬ_lbwD�0Pev`���{�6l5�#` """""""""��#�uF=֡޾�����s�g�c-3�iߞh�f'J��m(1��n���l� C��ք��0!%���TDDDC,��{�B!�J�����^3����ok?�N"���HK�����`��5K��g�K�7ف�X��3륇�k��C5:Pgʠf��������������Ì�]�	��yHA���b-ͺ�jgͅ9r�:�;�Y�4�0��kE�}���첏��qV9�:�G�c�c��������M_"""Utuu�	(�W	&�,���~�cAGFA&j���k�"""""""""��4�Mf��8k��������3�O�3e��U��Mw���h<Ȕ�`��Q��� �M��GSf����b��������������
Rs��E���B�/������Mw⅚� ""���}FT��BSS�
.5m�4x	DDDDDDDDDDD.��K����k_����۷����������P�DD���
�GT�� ��5��222�`�x	DDDDDDDDDDD.��|�ܜ������Ԍ�k;��-�ov>��Q�p�OH���񀠂�.�D���|��HMM��0�@�0S+������>������>�h���˰0gz�mm�v;��-��5%��A��!gD�P(J>�{,V�\	�a��<�7�%���oG�@DDDDDD�0�6Ӫ�?�&��f��?��U����q���2¸��i|���Q��""�	*����
MMM�:::@�_AA>��c����"���������(n��NBQ��_�C�2/����`�,J�c������O������f�&*_�������"iЕ��Bs��)))��| "�>8�(
�GW�˝�� ��g���"''&L@^^^����B{�2u?eѸӭ�� ��E�):'�4\�Y2��#M�Zfe�K.���
�������~�w�vCU�ī���Cn���e7���FBFTpB	�����n��D��������|{��Bvv�}Y�V�e	0����4шHsP�G"�F�uuuR��үW~���R���_[�	׼w^���I�A�{n3�@ `e����;��L��?� �*P4���d�p�T��e�]�A�c�����������Fl���(++Sj(wi��ݻD��K�N�O�n`����eۃx�r�}���q=f[��ZK1��0��NN�AKD����wH���񀠂�Q0�I�C�
L��BAA�}Y��d�#���������h�d\	5TWWC�wﶛD�-ǟ�,��^F╺�����1Zd4	Cy-A9�T��MC�������5��A�����dinn�_�D����v(���
NXAFVHM�tec��"""""""""J���4ttt؍�s�D�EӐ��1����ӱl�2xɄTNGC4^���쀂J����O!�#��$� �N�E����awa������������h�=X�r����ڲDD*�ѓ֭[���R����(V2�B�p�\��6	��:h """"""""""c������i�xꩧ��o�h0>��&H(�	'�-deqd�a����������������͋/��0C��4�g�	)8#*��";;۾%�����������<��鈘��TRWW��kׂ�M��GT�}Y��뉝�����"""""""""u2vSS233��D�8��/��~33'��k�""��_�ޞr�ԕ���'�������lKS|��Ѩ�����]�`�g�O�> �����'�ss>��&̵o{��}�����^iiiv A�p�~�V��V��ĭ����������FUeeeO�ATTT��9�0QltMÇ'��Gc8k�H���U�o6lC�/s��wE�0"}�����	��y퇎��\����2r����[AD�+�Ƈ�O��J	4�'����������IQgXpe���=��*/��q�22񭋿�s�������-p�p8����>�I�����5��dO�ųN¥�O������G�˸���Q�w�u��~"�D�z����|�T_2�B~~��5;;۾�����܌�""""""""�q�7�i�{�Z�Uo��q��+��8��R��Ph�y�;;;AD�K����)Gۣ1�T��6���k�p�+����ӴDD�\222z�	�HPT�˨
T��+�0�@DDDDDDDD�EEEq���N�_�]��^C�G�T�	qbe$�v���9S/�eig��s������r%�хK���3>�ܔ�S;�iO;!�x��2y�@a'� ��t����DDDDDDDDD.��DО��!K�m��Z-D�~J���EȜ�n����1�\:�3�+?5�O?_�w:ɛw��74��_�>���z<p��@44Hk���t|$���$� A�����,rYn��BjjlS"/sק""""""""�$VSS�ϵ����䀼.��� 󉒙�����+�)%Μz,R����eJ���}w�y;ںG9ɺ?�XIh��#�C�g�Rk�=D�_zz�=���d�=��s��B�Dn�W�81;#X�n]����~1?��ݻ�<NGs�����dh������$� g"%�=��33'��-��C�kqw�3x��]{�	""�KKKC ��I��BgJgaAD�X4����=z*++G�8���[{���(�kL�2�`�����|�={6��ݴ��=�eJ����7���"Z�A%�O�}��$�'���=A��a粦i ���@�8��5��/�s���YS�ȍ���8���>����͆�1?��ӏG"mk-�{ͻAD4�:ҭ�FWf���$7{��ݔ�7�Q�ϟo��,L�L�W�/������1�@DI��C��͛G��%� ����>�W�
Bn��YYY "w�'""""�qtR�J���������b�n�{&���c��綿�}o�{���c���ĝs����{4�ث/��s��Ky�~d���5�, ������,w�}yi�,ܴ��q�g�D՛��OT�����͛7�v6l�����������ʑ���@�8�h�8{�qQ߿���+�� �;��i�n�a_'"���]b4�V0�a��4Y��`5ިߊ-�{9�3�,��hm_��	��a�?)�gN=�^Cm�G�K�����J�� "��N;x�W�)���P��� #*�+�"��D�]4���sF<l�i��Z��Þ'�@�Kh�t��h('L:�t��C��{���6�������b'��]�ᗸ���a͌��ê�����v�����]�4�:AD�E2�ªU�p�Ǣ��پMFV�4UD�w""""�ɐ�r�K�,��[�s�X�DD�iBJ�4�t{�sϓ����w�����b�n��<e/�sf��|�������_>a6~~�e}~F���D�Al����4�3�!G�(�/+3���n�}mb���z����<�\fg��o�76���|DDc��s>�����/]����������͟���<ۑ��ۗ;�jfc�!cV`TWb��w��s-f;�ikk)�z���fӝ8q�!�gM=֞����O��xݞ���ʷ6# """������*oE�j�|_8�>��u��4��y::;p�f��㾳�b���5�R�05����Y9K���
����H�� "��*;�^�/�9(N/�����c�n�	��bБӴ��-N�49�2d3�L���gBf� bFPo���-"���߶����̬�q�S� �;@$#f�(���{���?�}ƞ������+h """r�W���i�\7�}�}�8�`�=��3O�O��|_Bw�<S��C�QTn��~��!�#��Ӧ�+�o���a���e�����`5
=DDDD	��d��"�\2j�'g~�����2&�[�>�хK����ADDD�4��t�`0�P(���Ԟo��׍���pݤ��H/�n��;w?�GV� ���}�#s�~eޙ�y�� "J���ܹ�I�u�s��ʯ�sO=�>_�w:~�����@DDDD##�R]����gM]e���CADDD�E4��w'�~�m\{�<y2���QWW��H8'Aϣu?φp�u�aҤI=��	$�y����m�o�s'�|�|��<��"J�N��>�>)mΚ����2|i�ܜ�;�Q�{����[��d����}>�o�
�/{�����#���*J��S�Ȩ
)�P>yf5k�	>�)���*��~�Y������H54!����7d�Οή��~��Q,^�و'*��'�����&��Ĵ	��lQ"����x;N��wR��O����""Eeii������L(O�m˶�U�م�J��d�@	�D£O���}����U���65��7�}3�d�D��������i��@  �4�+u]ǜ	s0u�TP��ӧ���Lj�� ""JF4y�?�^> � eW��ǳ�F��r���ܙ����	)Y�mM]ԇZ�������T�^�E9ӑ���t�{z��H��7��$P���:��E�3���D�?!#l=g���U�ð�4�e=��,�/���Q�Ş@%���?[G�NI/��G���s�t6Y�_5桙��{}L�(��j����b{kY܏99-�sg�(-߾�t�����6F���3��qڔ���~L�R�5�fDD����.�C�بoD$��{�m~�����УX)Q��X����/�/OL��Ϙ��.J1u,Z��������!#e�X��-7����T���()1�@DDD��x�ĴܘKק�O^��'����)v8b ���M��\�۸}翰7����j�y/�s
N):S3
���4��n܁u�[�x�:�T����J�?<�[}n�ش?�ro�uips�9���cV�C����wwⷻ��<5�s�눂E�b�v�X���uDBx��-�|�?�j��>���Y����㌩�`^��gI��A���W��c׿�
yHX��ï�s��ӛ���s]j���O�bk}�̟��g���O�\��OV�O��<S�w�y�續`�yg����"��R�>V�x9Ο~<ΟqB��=V�Z\C����'ۣ�v߾�p�+P�˵�4Ȱ���{OuGc���5uۡ_����ᶝ�����������?����<���e��S�4�_�wN.>�>�:2D�������%O��w��p;�!#!�q�7��#���4=�>#\���k�5>���324�{˱�݁�O�:	�^�U�d��P�����|��}�f{��D�����e|a�C+�;k�*�9�X�f�c�fӝ�;F��"�����M_=찵������ϳ��u�C1��/��������P�6��<T���&�Zw����	��}Y���aױ�Һ�ǒ�O�����'A�,�������U���x��E�?А�O?����\�DDDDn4C����iO	�hs���3BQo4y�`�X�b������%!9����%8����3�c�b�<���"FB��k_x����9�`16|����5�Y�#%��'V�'L:(ꟑ��W矉U����|+�@d���k����X�T7�?iּ��	iV_6�4�~��%ġ#���7.�,�[r��s�����^���q�Ϟj�)#���ɇfx�~3���*�d�c��|��L��>$o����KGK8�������U��z��(����b`�D]]���G%�0}�t��""""�(N����PkB_��M]m��iz�:���rp�\<s�Oq�s_�z� i�?s�M����0J��h�
�g�K�2���)�H�53N��W|�۫:���m�̜<��B��q7�a��M�F���0���wP�^��P�=�ƴ�B{^��d�Ǐ�_;\��q{��ո��k�Ȩ�����d}�o�)�Z������� �:uʑ�͡_6� �(�#$tM��~�^�S�a�}�ss>6�@���r�mw�y
*,�Ҙ���h��,�>��a�'ۣL����Ӛ�{1�@DDD��N\6��[[�;ӻ$P����bm�&�ݴ���ѻ(g:N�r�2��͚����sf���/����Q=��^��~�i����Y���i���2���_�?-:gM]e��/�A��p���|���~��	l�5��L��Ѣ���Ekp��C�<�L_��1�Ǌg��Y�2$�<����?��o���?v���s]0�C�~٧v7q9n:����;���y�Y����s@�A$�,��ݼo{�'������SN�&��H�~����w��Wڿo�<�}�/�պͨ��#,R�����c�}�ٙ��̬����x����V�6{J
�Z�D^��OM��dOQ!�P8γ֕���� 5��f{����/A%Krgx�o�H�7��&�#����oIX������������""""��gf}�ۥ���eoԏ#��U��M[ﳇח�C�wkk���f���/<��}�L�[�=�m�C>����������\�g�7���4}��m{���;�Qdڅx����r]g3N�������/bx��-�߶�Y|�w��}�?/{*���"|�����w�3<_�.x�l�������`�˸�����{��3��g�!���%� #3H�����:������0�C����v����������ǣ���X���i��ҷ~f?V����w[�GF|p���So܄�u��_eG�7n�s��6rϾ�y���&�r\8�D{=���'!ݗ���K_��*9���ijd�4���d,�=m��9���N�N��0�@DDD����D�f������4���[?����!ܯx��v�ኅ���.Ai����rT�b�l��~��Æ"g��d
 !������z3L?�r�Sspe���U����]��GW�צ�=8���lE�r��'ފ�&��]F6�����S`G�2�Foe�8���ۡ�������f?��K?�s�Lq�O�Ե�"^R�G_�vT��hIM�{�����~���}B���'� �U�wמ'���j�{�v㐁��$#w�6#�]�(������`�d��~��_��������h�I�u�i�z���Ot����gD5""""�1�@DDD�89���|��%�p���cz�x��]���pδ՘�U�sۧf}W���!������u/���`L#
|g�]8c�1X�=��6���Y�G������g�-Ær��y�����z��2b�L�1T�V���o�i}n���9��U��7	5�Z|$�(X�s��g�>�ۨ�?�?���v�g�Ea�@�*�Rf�@(���;)P�.-��eC�{� a�L�"{z�N��-����J��$��������i�T����ga�C{�e�/���u��8̠����p|~s�&Ȕ�T�Z���qfŎu	l+�0�U����hyr�o[����t���JK|-��o�ͥi���#�L�J���f�/G����F�=�6�ql�  �4\�S{�y��:��p����	  @A�  ����Q�丄�r���[�:Zݲ��[=�Z��N���Xn��c�:�1X�U䶹_kW���L�z�4���m/�-�����WW������{Bv�*��Î���pâ����-O������+�����������v�,o}�}�(_�r�ܶ�����,S�H�@|����Ã_{���K�J_�*�8m�ju������KG�YF���2*���ϻ�1<��]yt��&��h������n�M�� ?��v�#S�I?���� �@V$R�T��>u� �@e_e�F)l*�x���=�?��h��.�%^p�+  t   �̙�����u�ڮ�o;���Y�����;��@Cy��H4��=���Y�vUG��4!ǲ�Z�A+�*���x�f.oh��1Р��j/�pQ�I.�ڻX��^�S�V�76G�O��X�f,3Ҿ�t�k��d}!�M����l�)�5�s��K�%X.~��:���O�'i�Q�[�M� �E���1rV����&����˶��z:�ڍz�OC�Մ�6����C����Xۉܷ�u9PsH `��e����Y��,.}]Fc�\Y� ݥ��\,-B��E�	����X}p��Xe t1�� ���7����Y�fI\\�X,��������[6���]�'�8���Mx�`�!���'���":#���eݘ�!��5�p��䣃�t���[9+�گ��^�?�F~4|���ٱ�<4�!?�������Z�	&F����l�q�^t[V���k/�3����� y�}ݼ���R���}M}I�_�t���j�z��u	��r������;��C���@�$�殒��R�I��C3uƿ��-/d~*��Ҽ���M��G\�^ۯ�tԙr���  ��%�۹߽     ��xx�m�ԩr饗:�T[W+���@C;�SS[#l�� ����<-�}G���>?~Rp�L�m�ގ	
7��m\I�.������A����~ӂ���/�j�TM���m����=����q�}�'�-I��
w�O�?6a�}���_fƌ1�t[��:��H+cx�&�QZ��n��&6�Gy5�nC�eo�[�goE�O�ZӶ���h�B�}��Dk�|�Ϟw<j���K{߄Z��95y�     �^�@  @?�ႛ']*�%�.�o3-z�)�A�	2<,�SǊq*�F�����y��N�5H��{����k����fvz��5�ͯ�'�-m)MwY�Qu
w��������h-�05z��:�hK�Έ
sY���mJ�M��K�+���8��T��i0|A�l�(����OCA'%MwZ�U�/K��I_��,C~����ٗh���y|��9�?2~�9�+D     ��h  ����PIII��pT[_���i�~�|�=������L+��@� 3�6&b��0��;Җ���;s�g�;^߿Wf�k����:r玗���Z`���I3�tϴ�ʡ�r38�i�F���:�]����-T��߲�@�<����Z������k���≮P��1�H["q�}Y+a\��@���b��\9r���Ꙍ����I2�Q�%k��>����n�$��hIb�Ç�J%      �Y  ha��F�U)����okq���A���~&5I�����=zU��w���6:�v��c��?���D�z(���k$��H������=6b�|q�}2$4^�[eC����O��Q5���� ��C�2��V�M��L޶jP��.k�tY�Au�֔7Tw�qԻ>���~�h�*!m��]yLm%��ǖX�pNkD4�p��N�4��tF�h7�J�������Vi���
)����U�]�������MZ�]I� �fX���ɳ����;ټ6�5?�Y�#<�ooS��6u��7    �#�  @M~~R�����A��-^߿�p��Q��i��Y���E�%����cje��O���0����Ȩ<h* h ���ZM$>8J9��^=/mGp���+S�/�����oV�X3�q��r͆ˇ����k����R�����>N窴��8Z��x��.�n7��c��Wʫ�_���F[J��4�ժڒ�1��>�����ʓ�`ki��^h�kJ$5<�i]b�
8 0�\x����'6�o��*}�`�h�<���wk�bYg�    �G�  ��`��W�,�Nyش�����G������/n�Ω�dhh��:�vp��������G���8?���<�񑜘8ݴ>8%�����rz��{����G�_{�����<��}K���By��W�vO��⣭�U��'�l���Y�k����Ѷ���(��V�F.tY����Q�a ����k�      �<   }ܞ��a�����:��ސyrB�4��`s��Ы�u֑�N���U�������R���o2�J�5����Y��y���~�~~r��_���,Y��ޣ��
��cw��h�~OE�r�N?���GQm�˺�󾑻v�,�VB��S�S���v�\�1��O�����oQ]����R�s����Z*�+      �<   ��#�ޓ�G�)�cF9���ԫ���:n�p��y&�H+3xfP�����x-�K3)m�����G�%�B����s����{h�`8��l�ZȢ����㤴x>�ؿ�`EQ+��a���aO�/�͸ƾj	����d>�6��/A�����b�RK%�5-f����
kK      =�@  @?�����iy��۝�?I�r��������O��e^=�iѣ�;�(˒;�^��~S:�:�"u���GĎ�	�)��<��c�F�jYU�^=���#]��Z;N�GY�cw�~�us����|�2�� �͢��9�y��~���y�jI۰���      @�#�   �O���F��ٱ���eҥ��9-�76�./�4Dѝt��'��9q�drT��mG'L�(Р��O�:Р�����n�������P�h��x_ݯe�A� l.Mku�5�vH��NB,A�uZ�cHh��V	:V\W!o�_!���o_��C}�-I��q�ZR�o�j�=A���ʵc�qY��`3�3 �ꎒ_L:��T[_'w>|�466z|�y�g�Y'�5X�=7���    ���  �~��/��G��NV�-\��~-�DTZk�j���|�t7kS�iEq��T���Bb=>��ookቨ�0Y�<�e��L<���r����=�W�s'��%iR�����f�PÉ�������#��v�,p��8Ԣ���כ��F��=�z�}�&ɭ|G|t���� 1Q����QC%##����b?��j�&m+�];-    �i   ���9�dki����7M�Q���ʆ�娀p	���*埌:]�B�'�)vY����Sg>ҫ���8�%H�W�{[���Qgxh��Zz+gE������)Р~;�<���w��1}U��T�6'6?1_n���\�r�ӶZU�����9g�1��x�dV�y��vn��c��3]n+o���2�k� �����U�!22R    �� �   ЏhU����#���؄)rB�4��`s��Ԗ:-���ɉI��A���,7O�Tz��$�u�5��L��퓯������>�a򗉮�����?9i��1x�,9����>h���QC�U��X��~�e,�['��TذI���g��\��.A����D�sտ�V>yn�L�G�g)e�U��`��ڼ�������s[[Dh�w��L��������/�" �45QU    4   �3�f!�N�\�DqZ�U�
4�=�C�7d�Ӻ&\"���K�L���׏���{��ϒ-�鲲p�W��Y���'���P�ǫ�]9ra�s��V�<3�.��uP��,�+,8zb�o�Ϯs��CJX�<9��.���Y)j��oI}���Ǵ���_<�$ɮΗ?o��[�Ak����W�Ko�U�ze�]S��&6��%�Mt^���xĩfʫ)����U�J�ɷ͓Vk)���Jk�	���9q�dA�l9m��m����w�� �E~�w��YZZ*��ƺOB���M�-=S�˗*�VVZ=���Pc�    �   ��R��n��|�7A��鲏V�cʕN�O�*μV�����ʿ-��ⅹ��1�̲|�5`ؖ���#G�Z�l���ޗŹ�\�`�E�~��dd� ������NO�U�~��ӐB�@���u���Yי+�[�q�SfP��ǡ�/>>�n9�m��H[�=�@�n�H[�a��n��?w�)�;Μ#��8�B�=R~���K��L~6�,����������T��Y��b��+
�
|G�D��E'oi���5w��] ]�$�P���K3���(;w�4?=�q�F���w1��?D��&>P�y��5�Y2\����R��n�    �=4   �C�g.��N��\���Ɖ?��W��e��%{M5�S�g9������Q����o�'y�W�kE�9��傔��z��̓{ߑ�ƞ�����NfXr�kYU�M��]��r���^V>:0\&G�������h�ciUO�@��D�Ы쟝�G3(�x��U�Ӛ#��b�[�;��՘sL���44��o����\:b�	5L�L�o�?$O�/���>��%i&��U)�Ō2���gH�%��8�oA2*�ܺO���Ě��������6A��}u�vs|Qm�[�U�I�12#f�̊+�g��g Ҷ��:C�PB�7y+g�\��~ڀ �q�����Kw�8k֬1�:t����/u��#    �7 �   ��56�=�^��������i�[�\��o5�����u�������7WC���wsW�����:�`����aǛɑ8�6߷c��5O�h)=�A�˾�[>;�^S�A-4�L��Z׼>��
��U�zݢAix"��P��p�Y����1�I�����?v����fW��/� K���K���o*Q�V���y����"ץ���O{?���r�'��	�<��T �7(����x�}��ÊW����=�"�A��� 	���R{


d�ڵb�Z�4r�H������IJJ�����A���$--MrssM���c��!K�H�  0 h   �tP�Ɖ��r�6z����.X}�����@�_�w�}0�%��Q��k��5wJ|p�tm/ё�.�_oz���XY�M.]�7y��?��m9l4�`��L���eŠ�8�"u��m���Y)W|s�W�����2��_�ss��R��3l�5�;���d��{�O\nӪ#��r��z��&8uڠ9rB�4�7�� Ik��ʪ�m�\�2Sqd��� ��5SJD�����:�N���.48p�L6pشi��		�!C����N#F�����/4����c�w���t���w��СCRk�.  H   ��jk����4���'��ˎ�,�}t ��/~'/yC��ں�۷�h���`�x��̥&<�`�,��8�К�e�f�S[ct����KnM�<3�n�>���	R�U�/ha�7�ʖ�t�c��A�Ai��?n~B��^����������(�x�9_���m��L�ǲ�|�z��퓯p�$�����Y�gں�Z�h�1C%5,ل���KD@���W�v5:�w�@:  ����3د�MTT�<���N���(�Yuu�=���4Ȑ��m�0  ��h   �A��4s����}v|�.�w`oop|u�v��rوS��؄).j�eݡ��ށ��T�G�g�������W�������:3�ʑ�����2/~�L�a([k1��A��픗�?�U��;5�ߒVj���Urq�Ir����вG~m�y܏�} +
�zu?_lqy�t���s��7L����>K�r�L�N5�l4���<۴�xt�����@|A����啬/��I� y���<SfŎ3�SKMVI�8 ��2�9�4o�l.Iw�=)o�vy:�Y��V�c�vW�p����.��H><���z^����C���~k�\ޓ=9�>�~�����   ��UVVf�]�����V�HHH�����$66V����O���TTT��
Zi����&��!���b  �#�   Ѓ�z �����{����t�0ARp��E�VՁC��R��^ݧҐ��-f�	�+��j눀���ט��������Jz��2��ɿ��M0��>���<���v�>�ŃN�ъ	�l{�L��"%4Ѵ�� Ɂ�ۺ�u�@��;t��g�:���#1��&�P^_eޏ�N<�k���M[����1������őV!��Go�^��_o��   ��h����|3��a��`7�Om[n������П����L�UUU%���f�j���&XQ^^n���d�6�Ep������֋�G� Х4   �]:X��z���};�J�Uf�I:��+�;C��+���z�U#OwZ�� 0P�`@@����T��4�a��������[�%�	  ]����    �g�'#�9��<�[��A�  ��J�v�s_`�Z[��   @�@�    |�7�~��}�	  ���
h��"}�СC���Ԕ�   ��h     8>q�����<6��H�  ����0�����ѣG����   @�C�    :iPH�<5��.������76  �]qq�����>ꡡ�2l�0ɒb   лh     7�5���<Ӿ<$$^�D�ʕ�%!8�iۜ�By,� �����Kee��v�W%%%I~��� �   �&    �M�~~��������j+�� ��Wc�$rH��3cUp�    �]��i    @/�����v�J ` �
ml��    |�@    �HC�U���e�e�s      �s4   `@jlj���N��Б��My}��Tʪ�m�\�2ɮ*       �G�   RI}��^�c<amj�      �	�       �6D�d�e��ojj���v{u��p9̾��u��I�}y������eC�/�'��~�ڗ��o�F�&   �{h       �i'Վ�[�����@�-��"eeeg޼�r�ڗ���
�_�ᔚqr�ы��s��7KEE���s�1����о<cկ�"�A    �       ������;V֯_�񾉉��Ϙ1cdӦM]z?    z�       >��~����r?aaa   �w#�       ��*++�گ��ޣ�������:   лh       �s����j���"�������~
  ��;��U�$++K%**�LZ�IFFF��CBB��@�      @��=(Ol}��755ɖ-[�`���/_nX,	Ji�q�BQ�7W�����ٶm����������'8U���  z��ݻ���_w���^�1((H���ͤAۼmY������#�       ���j�O>��qrssͤ%p��0�������ߏV��U�HNN����  ݫ��L�x���Ni먂�3�%44�Tsht���m���R       ��5�L�u(q�����W\(��KQL��Q���)���H  ��믿6_���6S^^^��DDD���� l�����I       tZfR�HR���sՄ���d���󿞷�   �����c�]QQa������[Z8[]h(B��54          �UUU�[555��:��b��[Xت<�lu. �C� �n4!3Bf��Ic�/�IS$:&�e?����)      �'ԇ�l9���mb�tVcc߮�d�Z����LYYY�n`��)66�����y� �"�  @7*N˓�_g�d�@&N�貍�'[��N�i �      ����$���fR@���KCC���-�Ѓc��V�A�qqq"�@C�          zPgBv�y��.((H���@          �r�BCCME8h�A�m4�,� }�  �������gii�455�6�|�����
        ����6SAA�����ܮ��Us�p�m^+=��5 ��wk�'h  �;��%���R��y���dРA�G]�a���r�>�A$T       �_		���2A�Ћ���n�5�
aaaN�-4�`���� ��@� �TQQ!{��uZ�/�       ���$����V��\x�Snnn�����mj|��:�@         �1u�Tٺu��oѶ����fjKPP�ia������Vy�=          �q��Ijj�ddd����:)((0S[BCCM[��6�?m�V���Ż         �Gh���;O�}�Y),,,���f���ks���p��-���b��'          z�T_}���駟�ƍ���^ ���J3�EC1j��l�-t�6���v�{4          �Q���r�g�)��"���RVVf���r���p�ohh����ɜ:�E+8h�A���m���B+A��!�          �W

����v���!��W��O�z�i�ZPz.����)++��m�m,�Z8��		t/          ����P3%&&���Vrp��P\\l�mW�����|)**2S[4���k;h[���8B>F�  ����*K1}����#IA    �[t�Y�uj���c��e𡴴T��4�S[l�=�l�=h�A��V"�{4   ��е%�Y- �ީnd�    ��ܭ�@��p'���VtЀ�t�V�A�Z��b�4          @�||())���&����N�����6z����`kmaku���'��          �w�V�U*++ME���[���^CUUU���zh�VpЊ�ƍ�y���CD�          ��F���:�G�jhY�e�]������Vx�iÆr�y�ɘ1c��!�           ��l-����`��'�00�{��+��W\!Æ���@          �a>>��� �����/�k��F����� �     @�<u���% ���4��(�*   }�'�����J����F�{h����t5j��  �a���f��+�W  �E����S �w�56h   ��bcc��w�����V�=4   �5�M��/�P�Ν+!!!����������V�K�        �[�|Ћ�l�[��1���+++M@���kB� �n�t8�`~�KLLt
3���@>|�D���{       ��U*ֿ��������N���*h]cc��'           =�ӊ� ��?h           ��V|p'�PZZ���'  �F�#e�%����N֕�q����_�  ��K%�*_  =��rl�  @��V�a߾}�s�N�Z[C[,3iE��� ���7A@��Cee���h  ��U�<e}��%   �y:�c��`�  zN� �  �~H�2h��?ބd_���o����L555RRR"iii&�PWW'UUU�"�          'A�~2���v�� 2Q �����c[
7����i�С��tX�d�:tH�         ��R/2$���6�a~ ���� S��C�           �:           @�C�           HJJ���B�oh           �bcc�C�    �>ꧣδ�p`��T��e#N�PK���4���u{� ?�\9r��5�S�%�v��V�="v�̎'�RZ_)�f!}��^�cF����2#f��GJ|P��56HI}�dV����ݲ�p�[�ǰ�D9c��6o/��2�WZ��]�_����g\�091q���l���>u���9qt�$9m�1T�Cbͺ��Rɮ*h>�6Ȳ�R�P-�!�;���B�'Re�u�nJt�?پ���3K������k��|�����b	��8U|iɁ�eu��?6a�L���q�T�����\��9��Nk��(o~��3��,Ӽ�8w�1���c}*�#ih��y��A�eDX�}��ϛg�t���_f57�'F���(�k�<�5f�yo*�'_5Wmk�8�>g��p�l+�   �/AAA�!�     @��_�C�.��G��{���:�����Q����s��Y�g_��a�_����Y���['_.����}-Р��?Y�2�R3��v�iK�ٌ�m�N�!����[�+l~o^��T���U9Ps��m���d?���h����F�*wL���Ar��1g���}�^��zͧ��!!	N�û��[4h���8��������}����{c4�[B�~ܵp���@���O�kF���q��\�j���c �g�ul��<|d�{n?n�x�W��3?�k�繆F^>�F\�ilj�'�?oh��ǩ���͟GǐDK��dT�5O����笮�� �   �     �G�L=�i9�?@~4|�<��-�3��u�_�*�hP��������92n���0�|9��ߚ� ��-�����}:o����`�tVd@�yn�$�^�W^M������l�@j������_� �ʳ���4�G�l�RS��&G�ʿf\c*�h��P]y�?�s��fPZ!ƛ@�~�9�V�?��jk�ՕIt`�9�mRÓ�   �gh      n�j�������:��Z���k�`Mq���S�
[=���l(����B��>H�8�>�d_��4]���|���T����qL�P95��>��if������0�`mj�����~Dx��p��&�4ذ���d�ҟKfU���-*0L>;�^�;־nE�V�w���q�:��֙uZAD+?�l��fP\��uYq�?��/�`^��48$N�s��m��^�_i������m�%���P����n��,���K�ʣ��w��9�_mY��J^�t���o��1cLU���	f�V xu�M�����G�qk���?,j�n��}�h@hB�gc�����������f}�yp�;�4o��V�ׇ��v��ja߅r:�V�
���:����    �>     �mzu}���?'<��LNL�n
�E�2���w;m��x���s���J�4,�� o��ʧ�����i'��$���KwЀ�G�l3h���6>d:(ے��]��Lx�ۻ�]%�%Lu�������y��i�����7mFTL`��u�e��{�[q�S��-O��;_1����ZU��L/e}&o}��`�����V�Ct��*�U��p�<����Ux|n<��A��� �-АS]���mI�<���m�Y���y�r��r���{t��f�V�89i�|�J��|}hg��~~�'� ��!��՘ß�+R��[�t�8ZE�գn��4 ��4 ��UZ�C�	:ݶ�y�������Fvx?�x�    �h      n�2�WK?��L��䦉?:|�ȅ.����I?�#���Ӌ���QPC '}�{�ӄM��4Ԡ���9�,kՀ���ov=���ǚ#6w�xɭ
:8|ު[e�qw�J����S���}��t�5E;�U�рǟ�_����@Q�P-W|��8�E{�����w�py�{�W���'Җ�Z9᦭O����a�%�*%f߯�n��8PsH�X�V�   ��h  ����ȑ��$e�p9묳�n�k�����q�X���]2n�x��|��
�K��;<ƙ��$�)H�=�<I�Op��郟��V  ��6'n�L�N5�ڮ�˂o%��Pn�x���8�d38mk70P� �5c�g_~2�C��Nh��޵Bh����1j��]�췹~�E�ymq�����W[<���\5�t���Qg�;^��:Bg�5�ZUB[��kǞ#����S�4��Dm��.�.�f�e�t�N�"u�}���e��4M6��1�M����f����P�V���ρ�a    =�@  =���R�����Q2bH��m5�5"�������X�2}�4�c����v|����)�1	�����"��0  �q�RO��렠�M�^�~T�$��0=�_��\2���3��ȝ��!���rbp�ǁ��]�-6����76xti,y���*	W6�W��~C�ۗ��Ã_���
7O�T~��_gy5������n�_mg3*|���}Ϩg3�ʌ�0�zuh�l�)�Ii���w�     �     �C��`�h���e�Z��ٌe&Р���@4�O�i��*��7�9-{SI���Y�ymI�V�
������
���SͲ^���u㖧ea���@;��zC�T��'.(�>�+X8��q����
��v���Y��`�V�h��9��&4   �� �  @O��lZZ��X�B�&���RXX(;�v�����kϞ=�z�j:t�X,)((�����:�_�㩩���k�Jyy����Iee�dff�����'  ` ;w�1�M��+�_���<0�f����#$%,Q��
d ҁ�c�ؗWm��bv�8�em�c&����jk�W�eE��G'L2��V��nK�������� �mS.����%8L+���J���Q�arް�̼�Z�&��D>:�N�7d�5�g?>_��V���* ��Ǖ��   @�B� ��r8� 999��o:��n�,����ty�ל�U'����zY�|��\��i}��  ��~2�t&p����D[WK��
y7w�\�r���|��cǋ2�Eكjsi���~�j�9�e�>Ps��㌋f�������m�>���^I��rЋ��7o}V�z�	4\0�D�G�k&���L�J�����������Օy}?T����v�d�������Yh˟���ۑL���*'�UyN��w��V�i+�n*8�l*�']I�sl`����Z#�m��   �     ����e��,''n�P�X/��2���hPW�.�;w��2H9�9fjأ�i��ٿ�1C�����W�rl?P�N����l���@��;���H~6�,ȹs�r�W7Jo���&\���O�/�0Р���ۗ�-!�cF�գ�p���̆�=n��	����4��^�J���ZՕ��fZ�(�8�bHKqAQN˺OW:1q��ܡ��   �c     @�4���]���s״:(���uf@zPH���b�	|Y�Y��W���Wv��+�n�9q�ۼ]�*?oխ�C���8��r�#�ɔ����O�*�&�],�������UYC�x�������]I�<�T	���暁��p�j�C���76���ߔ�>�-�ib�p�?��W6�ț�W�lcV�b��̲Vih-��p���z��Y    =�@     ��5�-_����K������mс�+:�ZZ54Y�Ŭ��w�~h��<�[�?9�2����
��󗵻�VHz��^?-#�(���>CB㝮�o)����ch���a�w�ݛ������o�=�7j�uf�_��w�����u�j����[]$����]S�1��Fz���7�6?�����
:}�(���[di�z��}p�by&���kY�eQ�i���rVHy��.�.N9Y~��c��tTeu>�B,�ҕ���y6c�[��w&   ����F��h     �в��=(�W]�C˧��'�y����7mn�\�2{�ἡ�ɵ��+�[���nq�xkv��0K�Ӻ���ǳ�2W���3?�(����14�p�A�x+6�9L�Qk����]���F�i�l?Y�r����Zz���
�>��X�|>|���}Y8#���Yb����&篾]�?�ƣc�Tz�x�,r����TJ��]��2>2�T�8g�1�J��N۴�&Ӳ���y�  ��TWW|�@     h�VZ�YQ�U�E�lw�̪<�lB/v�<��a�>��{�����mfǍ3�zE���mkJ�hў��Rs?:0���FG�^w�˺ߎ���7�gn߯�g��IW�JCC̼${k|�0��>��ڎ�Pt5��g�kr�EfY� ~c�W_����<�>>(J���[9w�1&���Q7ɜO~%��2���1x�i[����Ӭرmn��I��p�ȅ��I����c#�
   ������C�     �J��`��e���]�׾���D��|u�?�؄)������ԥ�GO�
�#�&��q�?Y]�]�|����z���8�.����
�)����j�928$N�D�ʏ��7�-��qњ;LK����6#��������]�ҡ��~�|=�A����t�K���|�:�D�͡]��:s�   �\P�4     �V]�r�������";˳e Y^��hX�<G_�*k��zE�uc�5�)a�rT�$r�DD@����EeC�ܱ�Ey�k��/�W�������A~��߲i������c��ʳK����Cb���Gz�����\��@n������[쁆��fKT`؀k� �j�3��6e��� �Z     @��͇���%�n��3bFۏ��O�@�W��~�����/6(�?�����X+���m��s�ǁ��SO�Ȁ03����. ���K�w�(�����A�QgIy�� ����@~9�l�|������L���.>_���2�򀼞�ܭ�F�'��"u�	��ye�\�2�~�E&�a���8  �j��3���fT�U  �J     ���Q��*:8x͆KF�{}@��׎�������<-M��[J�eɁ��W��m�U���Zɮ*����Z+��{On�t�Y�h���T�G�I���'�O�Ҿ��m.M��D�ܼ�Yy�����/��w� �];_��F�&!� ��aQ����|�qP�9v����/< D�7�(�SC('$N�/
��߾�<[��]%�|�.��)W4/���ʃ   t�������KII�TUUIMM��	�!�      \8.�*��v�A�U�Z�]K�����i^�F��}���8�T"�*w�����~1�zϮ����'�؈��
ū�n��_�A6��kw?}�w���4�M�Ho�r�g��	ȴ�Q��V��r��L�
�kpÄK��􏥶�^|E�S�R�MM�J�n�mB��])?>�,�w�c�A�~��rR��7�ɏ��[N[�gS	�Z�   C@@���j�JCC�	)TWW����̄����СCft-     ���}����A�R�g��o�0�ߕ0�@�^��u��+�n4����˺S6W�?����U������\a~A�	�[U4T��k�'=`�ڏ���'�o*q<����@�>��ϑ���������6=*��2�7�Au}>�{�Y�"=-��si����)HI}����;_��G�a�DS�A�(��c��˂oe�g�L�;�h����ڍ�P�;�\Y�ͽ��Q7����ϣV�Ж���펎�,�p��1x�[�#���{T�h5�'   t���_�+**����"##����^UAו���ڵk��     �D[%�U�J�￶�K���b֧�@�Y��Ibp�Ԗ�@�Z��f`��90��u�����L���%{eGY�ՕI��^b��%5l�;ּV6�˫�{���{d���e�1��\����3i�۲���U�/��:3�}b�tӪ����(�m|HK�}�_�Ί­rl���st��o����[	����}��Ҡ��O��*�(�$���*���z��������]�r�<���iY���6y����6z��3�rהE��h��̕��c�guhh�	38~���I���]�5͊   ���4���&h[x�6�z**�=  �)z�T��'�\ ���Uee�d�/4>��O�.�{���ƚ�]�ۮ�}�t��Wө���r�������%<<\jkkM٬�~,�E  ��pe����^����y���Mr��i9�W�����yK�7�/���Y���Wۯ��*�cǙ�-d�,�ܸ�i���N鍾*�"G}v�<0����Ғ�z�|[�"ï7=,��m����-O�����W��4\5�tyx߻�>��k���7s���MV �嘳Ͳ~��4(5���:�w�O���Yf�V���0:�%��H���   �_ˠBː�NZUA+-�"�  @O9�A0A�ѣG�WGDDHtL��6Ϗ���,#F���֒Y�A��w�f%ߠ� IMM����W�i�!..N�Wn�h  ��y={�	1���b��}��� �^Mo���I����f��VݡW�߾�ӷ^�E����9+�U�j�g���aWh+����4�\����'�fʌ��f �ѡ�rY{h��*�n�RO�<��q6?'��dm��UF���+�-skm�q�W7��d,L�-�#�8m���O�7���U�mh��Qe��ǭj���!sOE�}��%in[C�n��9�)����m)M�����yOl,����<Q^_����
�Hi}����+��P���rt�d�<����4���|����;��:�>m�c�ȓ�K$)$ƾ�jˍͥi���1��㼡�ɂA�dB�p4���/��./�,�g~bB�O����u|Ξ��  `�ҠBuu�KXA'���V�v�4     �G]�����z]�W��56�%k�_xd�{f���_�C���۞��`]�n3�D�IBP�y�ՕI����oK��շ���}Y��L��W�Z�?��b� tu�$�����A����)���x�FA=����|�/z��VYi�Ҋ7��}��_�T�ϣ����mf�oE���%G��)��.�v;6hhKg�  ��F[:TUU�Tp����M�U�oi%���@  =$4.R��&yR&o����6��ѣc�$�Ȉ�Q�UW�r�2?��ɳFIDm�,O_/a���n�Ҙ%b   �PY}���έ.��hj���/��   $ZQ�Lh�DII	A���� �	�  zH��zy{ha�N-J�z�g��1�͓�g�i�W�����~S>r��0       �K��A����mJKK����?\��Y,�0a��'          ����
)؂
uuu��a���%�	�     z��I3ehh�*	 }ͤ�  ЛhPA�?8���C˰BM�{��?����)��"��     z��L�T     ��j���*��
-++�rSS� ���Of̘!��~�JC�          ���
m�����-�E"##MK	����%>>^F�%111�_h           /h���P\\�Np��PZZ*����'44TbccMhA')hp!""¬� ����4          ��-��VH�T����#V�`����̼N:�a.h�"�          `@РBuu�SX����%�PSS#�;LPA�	-�
�^++	�C�    ��I�ɩ. @߱�,C  @�a�Z���ʥ�B��
����$�;�
�����BHH���h     ��ݾ�    ����c(�Th����R OhXA�'�ǟ:ix��B�#�          ��i(a�ƍ���#���TT��l��ɶ&��4          �Q[�n�w�}W���h����i�в��cpAoG�@�         @�ٱc����Tb������
�
111f�\�y��          =����Tf �00���۫(8t^��b��@         ��a�j@�j��`-��`x��         �#���#�����L ��D˰�n��          =���Tг�jB�p�-�`k"@O �          �GX�VAױX,f�	����gDD��נ��kh���O�ވ@          �A������cE[h���:          ��hXA�	T���s	+h[�3          ЍZ�t^'��uV

`�#�           >`B	m��������`�1          zD``��%�x5�`��`���� ��          =B�Io�����m�l��S[E �>          �)S���ݻ��~,����N�ɱ�Bxx� �]4          �S�N�6HFF�����󓈈NА�c�[�Ao�� �-          �\xᅲx�bٹsg��h��D�v`��� ��          =&44T.��")((�����TПi�~          =.11�L `C�           �:           @�C�           �:           @�C�     t�0K�X�,�����_���w�U����?w'7��fP�Rq�BT�:۪U��J]�O[gk�Uk���v��Z���'�ߺ7(��!���������D.��@�%$���>��<��$&p�'�'�     �     �ᖜ�g� t=E�r�y�R    p�h            ��           ��h            ��        ��eff*##C����z�VKKK���:v8JII��n���㱮7�f�)
Y�0���F�Ѩ���T__ߨ�}���V>�O�`P  �m4     �N�.PԈ
�-�Hs� ���dgg+''G={��ڮ���,k�t&�岚�A������Ruuu���jjjTYYi53(  #�      :�	oߨ�5[���OJ�
�{^  t���T0@T߾}���g�]��Ƭa�޽{7;�3�������jEEE*,,��R�  8Th         ����2n������էO�=�Z����0d�M�8Q6�M��c۫W/���\&ckI����n p("�       $Qj�M�� ࠈ:��4#yF�$η���L~���c�:áf�3��#-C  t��
ᙕ��m2�{j�       �&��Q�2n�88���?�/  ��2�6�ym�sYYY���ZgZZZ�f�Ec�7$�5h            {+����k�fu�P(TgF�%�\<�/�@           h$�������#�<bVd0�Ng$�Ķ�v�}k�}ks�O��a{^�           �&�a�B���=p���ض_�k������)))�^u�Uo�vn            �B��;֎���}���sIJJ���O��\K�'�         ��f���tZ[ @��F��%�J�y�~n��}�̙w�~6�~�ז��         H:3Ȑ��.��. @�f�|>��������#b?#����=�k��|_c	4          �̊� ��0�_�߷+++;����p���[4s��Q�_����h      �&d�q9#���R Ԧ�b�������-�#?%[�����9�vg�&T���;��b�V�l  @G1�3f �����m~��*�H$�mވ��͍!�      ������iX[��5�9:��r#�O4��������M
f���g��K��7�E������e3�6����9�t��i��{�lJ�>���mzbë����U	    �����~��O?}�i�>H�O�     t	�U�:�V�膽�����k�qf*�֮�̖ϒ������u������VTmR�3Ug��3zO���\�L�WW�P�9n�u��������4o�R-�X��@�2\^�������7*�@�.��   $�{ð��  t�hԬ�?������o�Ώ�}_
�2����d�۝���@     �A�?C/��faҼ[�Y��eC^�/�r쵺{ķ4mЙzp�?�*{�v�=2�Fk���q�c�^_��y̪��=V��.��!  �ͼA������	5 @��������^1cƌKwϞ={Tl������aʞ�&
:D��nhnw��5nWx���c�{]     @�2"JKKS�~���*ٿ%��Ǔ�5�o�V����a�k����K�vy���V���5�Q������|�-���E����L��R&�u��������#  �B��*++�r�5 @'f�}������W_r�%�b��^x�Ŷ/&�%����iS�N�ݻ�@     �jsl:o�y	��̙����y�֔)S�=U�2��ġ�D���-�$��)�ewZU�t���)�FD�/~��0C����v�b  $Îh�>��������+��it�.X�r_U����h��T/ F�2�j�[�.�f��Lt��v�[��j���ڣc��{wh      ]�-ũ#�<2a�ҥK�lٲy�ƍk�u���V鼾�����r۝
F��?��h+�`�>)_ݨ����[[���ֺ  t���-Z�"���AO(Օ��\yy�6�n�����DO������.��cu�sN�������d�i�ۇ�@     ��a���Ç'm��׽�i�����z昻t��'���Dv�M����o�{��9�R��c����9���o�J    Бl6����b�%:I�     ty=z���1�i���&m>_�^'̻E���+NѥNUE�'��#�ݥ/k�jƢ�����7�.��S����3�     @Ij�0�&:O�     ty����<�Z�I�����rܙ�8\�q�;}��9����m�E��߯	'^�j��O�]¾c�~O���[�    ��lM�d6�-/�y     ��s8�<Ngr�J�s����z���ߵ�z�ҝ):5�H����٨+uR��:s�]�Q�:�!�4GJ¹�v�O듰oWu     �"�������a���h      ]^mmm�<OUU��&���D2<>��V��tч�ʈ=L����l[��*��3g괼q�>hj|��@�5�{�M�I8��E��ŏO�5F/M�_     $AM���Ht�@     �+����bu5�����HD555���T{��F�!�?��3�i�o��������X�k�5�:��ڬ1=鸜�	��*����/�     I��0�9I�ϗ�$�     ���'t��'����`�JJJ:�֬Y���>����M�]Y��_����}�����z�'V���c���C��*    ������\r���@     �3�̜p����$]��w�Z�qA��ؾ}{�=תU��h(V��GdԂ����9���T6:���/薡_W�í���AW}�k    Нh      qw��|�4��{�U�ᖥ�3��VgP�Լ��&���W�j2\�:�������[^�¬���r�����z������B���\��M�5���xI��m�%���3\Yp��#ݾ�	k9�D2��    �+!�      �~��y�\�P�x�&f���ܩo<U3=_��`���w��J�9�#_I�^o�u�2Sq���ʉXUVM}J��{A+�6)Õ����k���ָu�B�e�kM�tͿ��+n~��s�׬�/l�P�+�Z��tg�����ɹc5%�(��`���     ��4     �FVUo�	�n�mÿiUk8;������Z�=��U!y^/�DW|�K���oj�~9��&c>,]�o�K�EM�����O�ò�z`��V0���ζ��� �ӛ�҃���ʐO  �D�<���[e�������  h�     �D؈X�^�񱞞x�����n�齏�o���H��9��e��/Z������
����9V㳆(ǝi}��֕轒eZX��~�0�2�s�c�U�a�7�Zb�A�>�����/� @k�9����J���  h�     �,s��c�~O?y�~2�
]��d��˽+���W=+��<��m���*jZZ��j  $K�mWyUEC��]E�خ���+++�j�
�ÊD"J�?|Kh0��pUxRO�K��N �-h      ��;��H���  8�T�J?�}��=���O�{Z+t�A��� �"�      �uR���5�vN�k�e��z���
G�_r�"č   �����~�  Mh      M�8ܺw�U�}��r��*���ŏ�    y�+����|]_pN��. �8     ��c�G�o�ܩ��9���ŏ�,X-    �w߶�5�b�t��f ��     �˱���XU���a�cza��   p`}X�Z���G������f���W�6WҞ{�Q! �4     ���G|�ښUnZ�{��   ��+�  �      �`n^��fo�ߦ�s==4(-_��)     �� �      �Ƽ5�Zj��� ���/�̓/�C_�&�      ڍ@     ��3̐�L�@o�BѰ6�+����~�n|�5      Y4     �F�S��ظ�ta�Ir��:���ĆWu�����]?�M�3�r�p�Yc*C>=���zl�     �^     @���ѼS��́�Χ9S��a�P����_��^��s��{�շ+�����*T+     �d �      �n|^<��[�՛E�6"��;N���+
NS��k��J���z��d      IG�     �]��k��/���O���}�\}Q�E����x��5u��Z\�V      �     7*���>��?M����E�r�r���ʧ	3@f�^��~M�N%��]g.2���M�QW�j�~m�/�Ҋu��     ]	�     g�DC�^_ڤ�	Z���5�d�p`�m6�~҃:!g�u����uݢ��y�D��o�~'�mo�v�{,,�BOnxM�n~�ZF    �Ύ@     �3�/���o� O�.��e�j���ސ�a�����t=y�䱻5}Z��U�QE�'�ӣA��:-o���e�c�G��%�	    �Ύ@     @'18��~1���ZKD��}9���z��;e�=�|nVUon2�ewꊁ�駣��B     t     @#f���{��/͙bmO���`M�1|;��v��:f(��	߷�Y��~4��}�7���Ć0������wY˅$����Mo���?��y�?�     t6     @#fh����1���f��]��~��Y�u��5M���n|C�v~��@���U�;�Zf�O�l�aOա:+�     @W@�     � ��ӯ��P��\w,�E�\��Dk;o�R��
    ��@     ��~�v�Q	
�3s­�ty5c���.屧�[G�b�P�B     tG     @\E�'t�郦���zu�ǚ�u~����ɒ���Ά�    �;"�      p��I��Aա:ݰ��_gVs���O8�oj�^�t¾3�բJ  �V�b��[�-O�GC�Ӥ��r-�o  @Kh      ��;����,w����ʂ�*T	��ǣ����޴���V_����"��~�Óp��9��54a߮�  $[`�O[�Ա��i�oҿyY��F4  ���o�      �4g�����N������]����o/џֽ�Ek���րɺ��$}P�B37�ҪkK�2b[�aM�VW���]?>.g��;��    �� �      ���7N�s����jvL��\M4�js�-�w=�ʐOh�s�km�
o���&��{��g���O�����Z�1�%*��l���:&{x���FDjwď�z ����t:��	�Jv  ��     ЈY5`��?���p����՚�s�VWoUM�NN�C}SstT�P���x����Oր�\���NՆ�Bˍ�d��k��R����7�Y��s���4U�7�  8��6k�r�J�s�=�۷�233UUU��۷��)_   -B�     ���G�8�GV�aY�]��w�\N"����/�OF^a-i��q7���5ؿ_��?�m�[����V��7�>�����:g.5��ck����\`-���kt�� @g�i�&  ��     ���Ӭ��Y����w����x$��W�]+�6�_'�TW�j�|_U�Yط���ٚS�����K�N�&��r|�~6�J�4�|�Bý+�Q0N8���     ]	�     `��]����2b��>��0Þ���=�y��]0E����[E��#ܷ�Y��i������t���������b���:<�r����N������    @gG�     XF���W�����[Z}���߶�f�:F�0tͧ�Շ�+�J�޺s��	ǚ�4��}�~��iU}    ��#�      ,y���v�o{��_��fm{�d	��Ț���[��˚�����������ܱ:��X��)ݙ��HPE�r}R����\B�    Хh      �P4lm�vW�����֖�����j| �q�x��     �4      K���ڎ�9�M�ﺮ��L      �E�     XVWo��'��Og�O�E���Z[�q����J�	     ��4      �{<��m�5�R=u�m�<�v���֢k{�N�5V�p����}     ��     �������j�>���t�Ӛ��MՄ���s�~1v���?�:~���*      �E�     �U�j�&�[  ��IDATu�����S�w�w�s�>)_��5[U����P���5D�3į���M�f�l     $�     ���U5�����oә�'(͙��y㬖���g�_��u/[�V      $�     ��ֺM]p�����N�	9�U��[���#A����r���\��o���      mE�     4kQ��  ��WŚ���t�X[��-�߯��R��?�vm  @Kh         �a4$���SN9�I��e����  �2           @�C�     �]���vϱ�z�V�  8�d��:��r�\*+/k�_�  ��4     �������sܻ��|ճ  ��M#"�V۫���9h���H����}%����6�sT��:�G�<E�r=��  �@        �V�����1�Y�eee�z~E��v�d�1���r�:=SN� ��D�     4���D��2OOn|M�}�  �rrr�������V_���-  p�h      q�Y���t�N���F\�;�_��%�4kӛ���Tf�k  ������)А��"  p�h      qOnx�j�2���iZ����7�j3#����jn�R�  @WPUUզ��~�U�       @kj��ޕ��U�괼��}��I����V�R�S���fnxEk�  �Y�ܹSuuum����Hyyy  �     Ь�a��%V��?��iڠ3tL����sw.ѷ�B��  tޜ����������`B[̚5KYYY־3�-�.  Ё4     ������/Ymt� �b�t]����{�z��	4�������#uD��5ț�T�[;��_��
�����p��::k�N�;R�R{��+M�a��՗hI�:�W�L�HP  
�~mZ�e��),,����  :�     �b�M�K�����rF[���#*���	�����(˝ޤ�kE�&]��/��j�>�1�����1��1ա:=��m=��?��  ���qe
Ik8�Ś�ֶ����U�p��B  �ch      �d�٬��늁S��L��o�+�?��ӓ_��b��.p�YY�I���D�k��mw����v���1H�N}H޾)���{<<��:�����@����-�X��`��N�K�3{OФ^���!(��մO~#  ������;�s֨eU�  @�h      	������
��ai��9sɂ9���jn�R���.�}��6��w��4:���_�_c����3��QWhƢ��\��o���R w.�Zfbo������q�~s�    �Uh      q�o�_�w�U�aJ��V �⊵V��[�UM�NH��>�l����[0�:S��դ�7O����z�[�y���|.sي������d�o    @�@�     ��7[���o.q�̦���淵�W(t��՛�mOwZ����P.�S���n[6�E�5�V�     ]�     �+̰�W��J��wJ��~I��x�p�^ٱPh�!�}����&}g��hm_��ʂ�    ��!�      �0o�ﺙ�Z��e� ?%[�8�ڟ�u~���W�2����W    ��@     ���mA��صL��a��oSW������^h��˓)[�a2$     tG     @�%�/|�;����ѐ._�K�����ӝ���ڈ?���zk�9Oؗ��%*�W    �Ό@     @'����e�E�Q]���߲�M�T����{�     �N4      t?y��y�f��_7�HI��c.M1Л�p̦�b��?��7N�NyH     t     @܄��2b�%k�t턬aZ\�&�Z�������1W+j�n���-�[	�����|R��    �;"�      ���'�7����ڤ���԰��:s��Z�+l�^����QW�ޕ�hh%s����������%��o����5/��
4��{�
�����X     t'     @��O���i}��vB2�<�|=2�F+��?K��'6�ڢ����%��C�ӫ�n��>��
�     �]�     �A�ÿ���W�����WX�b��-V�ŏ�c���G�I��%�o�R��>    �+!�      p�;S��n���hHW�b����m����ǖy�qg��q7�>�h������kq��k�u��OJ�N����k��
U    �Ύ@     �A`�٬f��]��5t��6{��{A˿�}�����GkJ�x��mU�fk9��]���     ��#�      pԆ�:���Z<~��{���K�������C'������ty����/�'嫵��H     t%      ���⊵I��4P��l�P  t�Tå�����
Fí��ishHF����h��l~ �C�        �.����̤;����f͚V�3p�@}��ߏ���!��]/  ph"�      ��l���뚜�Oɲ�?�M������k�   LC�mS�!77W   �h      ��b��F\�l�u��-  �}�ٳg��KMM  �.     @܆�힣"�  8���׷�p8,  �]4     ����]%  ��ھ}{��+++  ��fΜ����;"�s���s��ɓ��M�aRQ�rnuu/       ��$X���O?�h4j/]�TUUU��g���5k��o��J��  �d�����~V/J�%%%�M����&�ptIO^�UWG�       ���Q-\�P��������7ް����"  �)e$y���_\���nh         ��܀�#"�{�c���湌�am��}|  ���f�J�5�9��Oh      qw����s|P�B��  8tT���${l/ٕ��  :�0���C%q��kUh      q�{]��w�3     ��l6��$Ϸ!�y     ��"��"�6][�44     �ܨ$Ϸ&�I     ���4�_�BOlxUs��ʐ!   `On9�mK `߲lޞ������=���t�O����6�y      nꂻu������$]��d�����o��MoiK�N   ������s�  �u�a7��={��K.��y��w�M���a�ْ�<v�}Y��     @�[ŋ�fVh���	���tM�=^����{G]���VY���Um�/   `_<���v�  �[$Q}}���p�cfϞ�^UU���f�o� �&��a=�yl�`0��[�h�vղ)y	  ���  :FU��
.�mx� ]6p��t�&�m�����^,���ϒ   H$55�j �����\.UWW�jpϚ5���Y�H�������aX7fw�+%%���o,O�G��µ�Y    _�lս+��������'Z����oUo0ۚ�m:���kg�R   ��,CN� �&��wMM���}����|.����4     ��Q���c��zz�ɣ`-K1,��ҝ�   � �u9�{���#�|?j��@     h����4mЙ�����Z�|�z�!   �$�9 ��E"�{.�������75�O�     �S�˫�N�����{�l����⊵zbë�ǖyV�m���h\����5T�S�"s�ͷ>�-������Mҩ�G�_j/e�RU	j[]�5��;>Ҋ�M  ��a����e' �2�w��ψ����g̘��     �	�ͦrF[!�+NQ�3�:���D�m��'7����B�}��֋��Ө�9m�Kz���Ң@����������^(��Ӥ����F�����k�Q�*ݶl��  8��bf���� �əA4�2���W8>��e�ٌ����g̘1��n��X      nXF]>�4kI����s�HPs�-��1�-^*#�@rd:�tD�í���O�+�hr�89l-{�?���+'>�)y��%����o[A�ʐϪ�`~��mS����K�  t�@ `5  L���۝N��]wݢ��'�      �<k��5C�~��mzKs�.PM�NH��2]��+�������8�����Za������_7��d̪��zu�Ǻ��Y���ˬ�)     �(���x<+SRR~8mڴWZs-�     �Ħ�b"!]6`��Z��o�����W�����t���Ct�ag[�?_�l�0Þ�P�?J�<=    ��b����]�p8V������'�?��6���     Є�L��%'Z�����Z۲`�~�fN��+T	    ��HOO7+*8t��fF��f�p�݅N�s}����/�|c�\R֫$�      ���j��0�O��g.5az�p����     H�����l�Hk�y��7�b��d<?�     w��G��/۝���<k	    ����0v[���Uuu��n����e�ٚ\�ܝ�''�      ���3��%�,!�;5��a	��WmT(     �a��Ѩ�~���RRR��h      �b<W|?M��D��-:�O	��_�D��
    �f�!���B�     ������=\i	��a-�c9�g��e�     ]�     �.�$P)$���ِBa}��~����q�w�C    �� �      �Ř���Ss��     ��     �.����Ya��sFib�p}Z��     �N4      tA���~8�2��i���u�?Py�F     t      � $�K>���>�љ���i��m�f굢�5�Fcsܙ:;�     �J4 �^n]=A�5W�h$a��kv�:�0dD��}n�K�O<E��T    :�S��	{�5���r�{�i~��Fc�}���֜��a����[U�V���^�G}R�5�� y�.����P�     ��4 �^zڼ��Du��ZS�ط�L�W    ���J�i����a���O�ai���7��3�0g�����>(]!     � �������   tcޜ��9��W̲�@o����*��Umد�2��퐡��    �@     @���n��  �Hy�tMK=)~�֦��ֵz�T�G_;|R�xv�BmvT  �4 �^|���ի���h�~�߯��u&iii�z/+�t:U__/      �@����/�{Uhٲe��gȐ]��y}�F��  8Th ��ؼ.�u�Y��������Sgr�1Ǩ����W��      t��?�M����l  �B� �2x�M�pR��>�OK�,�at��g�N�����f�W�_#U�'      �#�E����  ` �J�����ʲ*5t�R      �YTW��bh �CSE��W��l{D�aC�^�r�lꕦX�ǚ�:Ή��M  �����iC���n      �Ylڴ�M�	��g]iT��P�we��U�f�{�R^�]9ކ�Cn��
<�xm�~n�\�K � ��,(      �`
�衇R0��ׯ_/����y����_�"~T/��n�2􋹍��K[+��fE�Is۬�CnzCu+��&����n��! �� hs���"//O      ��d�ڰaC���F"-_���w8���m���Jk[fh�ڠkҖ��+=dx�X�"}W����.vUpz * �����,���      L��k�i��ޫ�ۤ�.qi��i3'ȯ��mYaDKM�lQm�G�g���,���v�l�䴷���!�  m`�O������      ppէDU?��s'y� to������D��g�u�Q����}�Y��=��̥-�wWx0��Rm"� �� h���:u��    �u�ST�o_�j$G��   p�E;w�a�̗_^gXM%��'�=6�g�Z���4�x�K'� $B� ڠ��^�E{�%   :��FO   �Cǡr�0�.�|z�i�2S��vk)3�g�w�Mdp�!�  mP[[��b۶m       �+bU����J�J�	ǸR�wW�{��CV��
A4,o���	� h���2u+W��a�?��'       @��{�-�HE5�դġ��fUw�3�`.o���v�iW�[@�A� Z)�v�@���Ӗ-[TPP         �;y��
F����z0����3�ކ���o���J��v�: ���-���lqq�U��r��0�vX����       ��:^m�lQm�h~L�Ǧ�T5Ty�4�*<��9�s�iR��4
<Irĉ'�ɓ�=�y)�&�~���i�K�1���W,o��<P�5�ԙl�V�n��*T+   �3��u����]Oe�'    Y
��Z�9"t.��kҖ���0�CK[ؕ;��aW�4�I	���$�x���i�1�	�e����,26k��u��-��%���   �*~��i   �I�94{YH�!t1�=�Y��Cn��,b��~���)�k���          �Y��!�]K���&jHeu��bG	ǘ��R��f����K7�=S�<�4        �v���w�gď_Y=_���/S�����ѻ�w�囯u�R��n8ޣ⚀Vj8Ԅ��v�~\��5_�����
f�᫰CC准���"�         �%/��K'�4�?۩E��z�a���ѻ�y��4 ���t�Y�Y�˫ª	��vE���X�u�i����,ڵ��U�!aU~0�{m���h         IUPPЦ@CVV� ��v��.]|�S�������V����ڨ*��!X@#����ʈ��|��Wx�/ma.uᕵ���y�ç        $UJJJ��s��phs�m�k6�ȑp�?d��N_�V�!�UY�|E��5 ��=ԇ�-�F�5z��ؚ,g�P��e/��jTz�H        @RUVV��:��/ ؟�M�{(����f�#����U��>(vl�ѢV0�.�h`.wb�M͏I�ؔ�*e{���4�mʊ5s?'v�\���Erh         I�q��6]WXX( H�7��3k�>�����F����C3?��Ѓ�u��mh��m�I�++��z�[K_8����4        �v	m����߯��z�x�֭
�B�����X��v��o��>�#� P�>�4����Z)��á�=���� Q��<n>ؔ;�S�@        h��P]����]�D"m۶��w8J=j� ��hi����m���Bᇆ0�첿Ѓ�nSf����Y�!۫��-�=��w���        �.���k۹���p���Ҷ�a�4��1o�=� ]�����i@O�Wg	ǵ$�PRk(Af��k�к��_ini|?��1֥!�����#�suņ��\�:l���        h��+�`�FJ�o��~5��+����>C|8���6F��戦��Ec\�n4t=Tgt�s9���W         �`�	>�Vء��a[nv��X#����U<��IH�n��ֽ" �뿦����P~~~�<�����         t?f�a�g����Q���U�a_��رA��y�㠎+p(��}��h��<O�<Y���         ��]��ڬ�/��T ���ԇ���Gtި��>�%          �vs9Z|F�J|(�6CQ���j�BYU�y��k�F�I�!h           ���a�����Y9�6T�EUZk��/+�`���|�#B;����-�&k.          �&�%��a�5�>Ǚ���U��hl�FK\����Z�
H ����3��ɚ�@          �3+>�g(�̊��oI�a�ϐ?,tq           ]Fk�E5�������ڈ���*�s��V
w��h�@  �A�u+�� �YE=I��     :���î�.�;v�ТE��Hsȓ�����Q؞"gz�B�TU��*������l��3D��h   8�*��O       ���DTWW۫�������b9����v������c��o��ic�]�A�*��a~1"�4           ��h���l
)%v�␲Ҥ�f�a��q�V�Вb��         Є3l��Q^��	 ��u)��@C�r�ʚt ��?|         ��K�m����wK� ��@C�v�;,�`�h          ��Hu	ID���$�Q������+,          @��mׇۅ$!����N��U          t^9iv!y4           �n��D           @�C�           t:           @�C����Ք���vg��_��;���U
��q�3]�匔/\��k���ze�BE��5�3���>�*���f♸���Ro��B��Xt)lq(Ztqw��ŵPJK�����6Mڸϼ97�4D�L���swfνs���؞�<�.l;N''U���g��[�?��M���v�KH+������zM߳��         ��4 �X��S/��Z�9B�⏃��[��c���^�"�?\�[��V��%{�^���
\E�C��ڙ��O�M/ަy�~��v���d�m�<W���ۨ�雋��XۧԵ�����w8^�?�9g�{��'5;e�          T�/�%#R���� ��9.Q�������,����L��� e�*�7X�V��(�P����
�k�z]Rf��V#u{ڹ�s�[��g����n�Y��4y�����V��OI�{�kw���6c�׼��^q(�*CEz���oc�����
�	�_�y�]���N�{���-�          ��@�h������\��nQ�44�8|e
%���O�N���� �>,���~����/hyZ�S�o��F���Yש!��}�`�~-Z����1�u��g�ב�*���L          ������0'�����K��S��ox'k���W��>��}T�o��(��uP�&�zD�BZ���͑�v��Y;5e�"��ǂ��         4G���2����t:�d���)	�����6��:c��el׈�^��+�=�ᖩJ�֨��5>��'P���s�<�϶MWC��Дя��3�V��
���_��C�z�ٿ*}�椮��%������B:��e����K^V��P         @sB��Bv�Ma�����Q����wʷ*2���m�^�̺K#����G�6c%Nly�z�t����ז�r`�3wZm�a���!���A
p��]����2}��R��_w������о�L���]�0�	���k]��D��}��}��Y�Fu�*b�,m��N�������}:��
�En�u�V�1�����q��W����|�o         @SG��"�Guפ��[B}�j<��]��ꏬ
��;Y���}����=�x�o���Z�,}�ZԿ��9V[Su��u����+�`�KtC�3��uq���)��֣�\�	�Z^$�Y�=��I�c<>-a�U���ߪ.���ܮ�my쎜�������]:mֽj��:�f�ef��OꓭӬ�紹ʺ5-!&-[?$�=�|S-Ä?S�az�R븅�[ZA�^��:9[V�s1�i��*tiyZ�^���>1�        ���@�%.�p�^p������w�
�wt� m�ڥ/x����\pz����'��h0r�������V�z�ץ�1i�5n�o\�榮�ۃnV�+���B���D}3���V\��Y+16�o��5�ᯗ�_�>a��MՆ�2U"�7�n��áܿ�=�mv���<�	q�0�N+�a��a*O�8s��Jb�w7��_w/�K���]���p�����Ϸ�з;�(� �7�gѸ��3��i���ZT��VX����褖Cu�̻hG        �&�@�L���]�0�y���f��,���f�Tb0�����9m��O��ܮ�Wdm�ٛ��+>Sf�LE�V�1Z!�ܳB�O�/��賋ru�����[a�ʌ�x��0aӚ��NI����� ��ݾ�M=��C=��R���5:z��V�TT�~�K���sܕ���s��>��y����r�{����t�
��3;e��(޶_�����:Ą+��q�!_���
���D         h|5�.�C���=�zg~U���s�Ui`gn�20��MK^�G������L�U���س�̘i�p���������ͺG?�zDC�zT:�i��^�m�	�cTLo}r��V(�P_�f0��>Sg���g�u ̰�3�P]1פ�O�ie��
��[�t=��s���8         "+_�C /�!�E�1��WQ���m6���B�_�L����<-Mۨ�f�t��be於��[�"a��g�]��{�Պ���'L�E{���6�\�s��ѧC�*7�`�+��ܦ�ѽ�Ǧ��ĥ��o����
]�'�,���[���U[�����n�Q��         ����W G�4 ^ ��v3���R�n�a�=yi�ǌ;�PC�_�nZ򊎎�G���s_p�U�`Ezb��p��V�!�?��>�0���
4�JY���=V&�Q�a��0�!Lˋ�� ��q/�kH�c��        �gض�@C]"� x���6�3m>��~ݽX�fm�6�:�n=��?V����
:�\�8���Ơ5��kU������0$�[��Bw�Μ}��H�KӚ��:e��Vo4�������}�         �P7߱��|�m���{��>��L��W\��&�[9Ey�6ӓ�i����r��Z�n���Iâz�:�L��u_�;�i�p_����w�����Ɩ�����^y��>�ts�3ˌ�_�/         �"^���Gr.�H��k�Q����x'gK]��zz���F��0.����R����qw�������2s<��b9�ˌ�NY��V}Xj�[��{],_{�_�v?�       ��ԓs+}��a~�:^ �<���_�veش5ͦ�l�2�ڞ�|]�jz9��9����QOtO��W����]N�s뿬�%��ؐ�C�-~I���Ը��o�z�n]�z���uv�1e��,��s�ZN4�C��-�����ޗ���3���       ϕRy��\;��46��Z�5o4�R�ˮ�"�2lJ˳ko�M{�J�tkg�ݺ-���9�G���q'�{ײ9W����.&��K�[��6A��KӒ��)xc�:��h��Pjܴ�xt��J��80vg��[Ud��pDSaBUOi��Z�'[�	         ��sko�[;���EY�@��+9/@{r���*��.�*[05k6,�6^`�{��p��'�V��-\n�\�>6���ĖC�h�u*> B�3��ݲ�uyT�R��}����ë?���rR�ae����K/m�F�ȴ���L��{u�_\�!�0[!>A����H�        4[�En�f�
+�d��oU��}��Ҟ������~�[��BH�h <�i�P�?_��)
�	Ү��՚s_A���>���I
t��mӴ5;Y�bѾ��x�o:������5UL��ʎ'�
<�w׊���*��p��:2��F���>�Ϸ�n���5���Q��`*U<�g|��}�         x3T��+	'��JnS������BJ�,:s7Y �)+����3�������nҞ��ͻ;o�^��U����.W�_�^�����>K��"5�I+���F���ׯ)�^��ט�g��j=��s��m��[��$F���봄���?��U�)��fMM5���R���쟲k�         �EAQ�j
)VQ0U���OՄ�@��X����wu��Q1���a��K^����3w��9jpd7+��l����M?赍�k[N�Um�P��>�:M�=���9���)p�*0��s�Woh,&hrTl�zĸ�za�W��ڛ�Y��|����w+��Yj|z�2���Z         � 3��gH�ϰB�K�2ݥZ@�-ވ*ԏ`_5:��:�K <����m�iHd�R��w9ݪ�0q�k�>�����ۍ:��(+(qG������V�b�j�l��L�����ZM���m��19�uq�ct]�ӭ�_l���&�[�v���&���ȇ4(�k�qS��ʅ�        ���T��?d�ϊ
n%g�U�Q�H{c��������@���.��{I�@�qs׳����V������l�t}�s�n�r�n�v�NM�Y)+���O�ՎYZ����{��������Ǖ9��m3j�ҡ�b��5��ɺ��I����D5m��쮻m���͈��;�}�}�s�hU�        �T~QI(a��w��,��EMo0��CM	��Kׯ�}�;�Z\?i�:	�`��>�ۉ���a��6c���{�6c�_��5^Pቪ0U"��|j�1[�_��윭�bB�u?G�j{�~J��ЄE���Y3�J����������R���        ���T0Un�`�
�3��m�%4��}�1��+4�%^ >7X��i�s�KQ��:0�(�Pf�TS0U̂��}���Z/�S��?�Z^���Z�
k�W\oUn��{zw�/u��_�_w/*h�;�eiz�2�7s�o�~�.k���>�y������.��~�~!�#u�u�"m��Du���.��	*��        4]&���WNH�(?���-e�SQ�9ii�U�|��h�]�F���j�{�U��@�'Z��I�C۔�M=�L��9�zn����/WZm(&�8�j�栛t[�su��w�ᖩV[���p��C�.c��
�T_�"uk�stE�X���5~�3�}O�)��ۨ�g�k�7�F��xb���Eyڐ�C        ��Iy%����
�~�q�-�@P�o�;�h�P?���!������0'�	����֣K��	��+���(�j�ɴ�xx�G�x�oz���:.~�:;���[5��ٺa���e��:?ﶜd��� Ay6f�T}t�[!�[��-�O�5�S����z_���Ԫ��b���ސ�d���};�'��         �U�rk_��'�ܺ�����N�����:��`�����`�b�vŇ�uX��B��"/�/�����9���~�{���[�FD�*5~^��J�MՍK^i�ױ)+I��~��n=F���`-��k��G=�ow��MK^՚��uz������t]���f��}��oZ�R]:�	m�l��!>A�n���lYj�Tgxb�g        �'3�m�R�KB	%�T����vg��"��Cp��b�B
�ARD`��`�u߄��J.����󏇴h�ˊ�)5~C�3���5q�k�^�a?S���,^p�NKa����p7P/n�Fw�x���@�s��ag@Dg=��j����	ܾ�=��K�:7�p_�~��Ev-���E��[e
        ������*��;�`X!2�d�s�*�
0���P�ْ�[7.yYo��̾���i�H0�j؝�O�Ϻתa�5�����G�v>Ug��	ů���3k}�h��J�G�վ%K�O�������~����b�JY���=���Ԑ����ȇ�?�s�}?%�כ�~        �����P�	'�o���g뇒ͥ�YRn%P5&�(E�j��J�+ߏ*�u��Ϫ|�q� /Sٟ��t:I�?]6��5l�ժ�`�������Ű{�������9��I��ܦՂ�ݷ�c��w��D��s6����ת}p���Bw�&-[���DEW����я�WX�r�7��       ��U%���xv>AT��CVE��6WW(	-$���+�#���9ʌm�ޥ�W��r��,mS���ۙ���~�]����{^dUj0NM���}uӒW����=���~�<&�?\���ki��j��lU����Q����<w΃���R�!5?C�/xR�c�'��/�8��        MY~�i�PHH�v�X(	.���DJ6P}�6��Ct���P|�i�,��<`5���% ���-e����C�ExSY��� �#�?ִ��p�jg����ko��ů���O*%?�J�Wt�G�����d�{�SU~�#�{�!�Z��`�o����?����j,�:�IY�m�{�ۘ��T�X��U        45�yn���H�v))�eUV��Pm~�L�6�+�Pr߄��L�x>��1��3wX�vF�Q
�3g߯��\5&���<^��MǷ|`�Tk�U������^t�yNN����t�ۍ��k?�ڌm�g*\�������R�L�T�xf��=B�ꇑ�MPl�q�ۭ��L        M��.=�[��r������M�'D�P�uڭJ�~x a���@�e��.]2�q�6�	�m�?X��<�����
=4�}�:q�z�ץ������5y�#z|�'�c�[V�h��\_��*����S�QvQ^�ǘp�'����Vjܴx0��]�	����ܮ?g�}ϯ�R�R�       ��b�.���9W�W�¬|E�UE����,]]��'��|h ���{��O��Zf*,�����9���5&SM��e�ki�F�>�:��qĘ��l��j	�䥕z�	3|?�AE��U�|��u�W�����SZAV�}�c������W�o��3�j� �a���z��;���LX��b�L�R|=       h*
]���34�r�	&�J
%�h��@��T^0��4 ^��M?X��ts�}!>A�����踁�Ϣg�^������_�)+Iߎ��"�B�����G��SgޣE��[c�bz��!w�e`T��uT\�8�i]0�a-޷����)z�����g�!'͸˪&�غ���;�'j�ߪG��C�\�9�>�B        M���"�Τ�DS��������Bt��|lWT�}?aT�/`����×
e�H�\f,�(On����ڒ�[��O0;e�F�v�~�p��B۠8���n\�G��ymƪ���z�����^�+�U�#@�jwt�c��1Ǫ�SA{���U��w��]�>8^�lsd���ҷf        49�Q���H1NV(	&���b�fB��P�X%����
WCpy��7�fC�k��a���f�:���u�_RFa�Vf���i�1�:�<�ut�<0n^�����s�krUǓ�����)�x�cV�O�5;Y/n��j��͈���7�        ���,�346S5�TR��3�`���(���'�Qh����Z��� �*� �&����k���\j�<�}�3�h�c��w�<�i=q䴉�����:(����ٶ�hޣW��T�����z��x�e���
s����       ��)���or|�6�H�A6Ň؋o��@sߦ�`�u?.������C��Lq������֥o舘�
p����m�9G>�g�}�{W����,y��ٻt��>�I�D4�yL����ǅz�����֘�>��p�ڝ�O         s���L`�lq��AYSa�NZ^�@�喦m�e��ۃo���Qj�i�p}��ua�qzhՇza���-ʗ'X��M��PO�����y���*��h�{z^�ێ+�6�`�l���W$        м��Bd���`W|��o+��ZRm����!��&�@���e�����aw�iW`D����>W�.�������M?��]��vt��=�?Zт����"�B4��ٺ��)
t�Wx���q����r�?       �����W������q��J.@�h*&�Z�a�^��|���w*��Teؑ����\��S�����՘L�����7�9�k3V�]�~��>�
���D����Qw�2_�k��w'       ˸�dwW���6-����o���CIˇҭ JB-Bm
���P�&�,�3�V%���춿��;|�c�<ݲ�ue��L�z����+�kHk��z�>�2U�iK�n�g�s�V�z�tS�0�q۲73       ht��6�*y��gt8���wȫ��
1N���Jnc�ME���6�~t0a�.h ���4�߻F�#�3�Wu<I�%����+���k,��	��㉍r����X���C��W��T�0�?�i}D�P���㇤�       �9hj���>vYU���5�dݷ�
Β�BX a�!h ��g�}����Zf<> R���Hwt?O?횯϶M�7;�(� ��^�Y�������Wc��B�����}�A�k�C��jd�6�j1Q����Ҧ�$       �����W��y�6Y�bC�LE{�mIh!��v6�
�G!��B��*7�Aε# S.�����):6~��o{d��~:��0k�shr�=��SMK^Z���a���50��Ӆm�Y��{V�_���?�N�NP���<61k��Z����  �.۾|���^���*y��͡���      ���g��|4u}�B&����*��Vp���h���ct���r��{/T���Sp��{T�v�n���^񏺿�W1�a�^�Tdxc��V�Opw������o��]���m����7y�]<�1��M���!���UPPP'�EDDh�8�k�#       M�����#���p�{�J	�����	)�-�V�h�4x4��(��d�E��W��77���;���Z�V렘2ǽ��ݴ�U�+Ȭ���-���f�_x'y�[�����u�'�-'�^�1k�J]6�	=���2�&�����ιzq���u�bM���V�=�.�-**��ի�=��fS��9???m��      ��Ǆ����ժ�.��ME��`�b�6�V �-^��t*..�aNFc�&gs�.ݴ�ݼ�U����E�,�����邶�4+e��]�Y;�j�s�hO^z�f����p_�n�z�n�z�������Zu���������YX�wۋn��*> Ҫv�:0V�-�1���F�P\@D��2��~���+c ���ک�Ͻ���I�&)3�z��-Zh�ĉϘyW���_�
      @�2�X'� ��F u�,���8�L��0a�11}���
�E�e�B����!�ui�cuE��$O��	�ý/���n�κNk3�U�-"�����R�sNٵ�0�����jڶm+        �|h ���6��s[�#b�V�9��"k��2!>A�[�c���~�Y�(�/T�u;�ږ�m�o��hj�MO^����r��37UO��L����6{��c�{\��͉iQ]�B        h�4 ͈��p�̻�d���1�U^�)�0[w-G)��7@��
�	PX�i�P�V��:�$r.osXXk���VuӂcC�Nm�کĬ$e�_��m�N�k����?d�a��u�x�cZ��E@s��S�v.iii        �����,�ѿ<��W���N�)	��#������S}�TcY��YsRViI�Fm�ک�ܽr�]�>�H�VGgK��ѽ�
��V��*0��L��ړ�������5u�b͍��Vrr�l6[���n�:       ��@�L��w,S�m����C]BZ�l�ܡ�7~�O�N���]Uz�ck$�ͦ���tz����ݱj#O��*ԝ��֫��*= ��Ҡ$������ֺ��`�=Z���Ơ}��       ��@�L9�uO�u}��=�]�OI��̺/�Ӯy��gu��,K�dm��|O���5�O�Ze4&?��^p��ms�Ucm�6�A��5�p�_5���        �Y!� 4C�#����oW����R�.s��[����9���,r����9�vl� =���V���dZU,��n]���]�%�         �C � 43:��'���*T���=��g�U�`Ez��?N��(�J������jqj�v�q:���CL��TRxx�G�s����4O?�Z��;��G����wVa����)+I9E��-�r������-�?\��	
p�U����<��*���K�?���,         (����	�o�٭��XS5��M?ZU��m����vjv�J����}zm�������<�ɻ�!�����>׬�����;�6(��1k2��i�h[N�!�s����LЀ��V�c�ZA��:��H�	��g�[��         47�f �7Hߍx@#�{Uzܔ݋����ˮ��j�pr°
���ܡq�'*1k�������U�r��e��	=T%̰�X�0�[~��fӑ��uU�ubˡV��P:9[j�O��oל�U         P�/����9������.�M#ҠȮ�2}�n^��U������Z^�9):z�-�f��T�0!�ɣ�Ш�{���I-�����=����Z�ʹ�x��%V%[�Ge�}���8q�$MK^*          !�����Te5ȹ\�xW><O��S��~\}�;���Taxnݗ���5�
j}�0�`�6��r������oӦ�$5����2�n�?�E��90��a���Sd�֚2�߹s�Sk?כ�nT��v����G>�fܩ��         @	^�K�"=P�����ӡwUf�*��y<X��y}���lYV�ei��)v��ӿ<�F>x`�KH+���]<�Z�o�[�e���3^�;�P�A�o����5Z��U          4 M�C�/Ց���ݗ��aU������w{�suF�Q��ے�[���X��Ǥy�u�b���{`�vGkƞ�zc����T��r�3Z��A/��Fv[�-(L5�/�߫��\e�M����r�Tp�~Rl��l���]Ri(6$R����M'%        ���	7@7t9��}��:r��Z�oC�����G꿽.�p����^'--��k�/h0^����4e��:9���վ�,����V匊ti���^���?)��i�;XI���D\� ��*�VJ�u�@�� �����!�΢�     @c!� 41�}�+��Me��\�v��9�i�ᨸ�zc�M�o�m9{䩦�YZf�����[#�^��i�ur���NU�o�^pm��]��X}��WMݽX@s��Ӯ�ʺ���������s$$$h̘1����"}i�D� �'X-�# �>�6�   ��lθ|�U�Fz�x P4 M�m��U���r�ݽ�}��:;׈�^�rؽV �2��T�s��;n�?�|H��Q2w�ɹ^�������u�O��y����|�
�E��и�:ںo�����\.W��8p�F�.�#?���l/���^�Wh      �V{�*�7�4{��� ��"� 4!��a.�/ܻN������58����}y����b�+ܗ�)�ը�7hK��:9�ĥ�iLL��X�1=B��m��;��4G�CN�S����z^ll�        @�A�hBn�r��>�e�M��K�?^g����
3��U��~�4*���'/��1�ʴ�Ӕя��nҶ��Z���U�K�=��G=/�JJ����zw��r�yw9�����j?��     @��d;FC"�Z����?~��<�6R���9OF�n�����  �3h ���.o_~��O�NӒ}��<���a�T�2����w���z��
s�)L{��;�r��:9[��#�Ҹ����O,ڷ^/o�V:�\�9�����
hn


��[��;w�     �]|�ԯm�~טv���5zs��cSǶ%�K����  T�@���JEK5ȹ��Xَ�:��U`�:8��k�є݋��uj����ߙw�?��:9�i�����ۭ�Du�k�O���g�Ug�"jk|�txT�*�.8�
53�6-M�}8������Wz-�]��@����}Z�y�u?%s��:��$�j��{�*���ź_XT(��p    @}

RDD�RR��F  @Uh��]����R�~����~z���^��5�|>;ƺ�W�y�q��Z��]g;_�;g�]��O��iEzb�翨��z}����cM�b��r�����+5��j���7�Zω��oc��?fܡ�)+ku��9{��ue�+<���e�z�dh��]����Z�Y6뫔g�zX�<     �??�=��p  ��4x���P�jժaNf�_����j��.|�Mւo�#@���؟�*���պ�����UJ~�P{�?��}�o����_��4=�w�բ���j=ڪ�p֜��<-Q�|��t���3�F�?�~��N�u�~޵�V���M?Th0�������&      �S��n�����YYYTi   UF�u�,����Zef����Ь������vQ���1G������/��joT�*��g� |�����,����BM�q��R��6�{��za��zt��J�KSC��l��\�#b��j�`� }3�~�7�A}�}F��Y�w�VglU���sl�       ht��ڱc�u?99Y���5�g��ղ�J�8��w�   *C�u�,������/Za�]N�MYI�m��h�n��Y���=Kk���$�t��n=F��`n�z��w<Aϯ�Jo%������\ã{��Χ�Ԅ���MI;S=ᓡ�t�����/k<�	+���
���      4��Sg�덟X����S�y�y��*Z�j)�$  �
h@�ic��IYU�q�Y�m�_�P7�U��=sϊ�ת�k���{�?����'P�v;���[�O�NӏI�"}�
\�5�3��QѽuL�@�e��QLˊg���j�1a�sVK�ꚞ������-��PCU�       ʓ�S������j������=�oɛ�  @�4����[��~���ə`ݦ�gu�Wh�r�kh�C��[��jh��;Y�C�/U��@K�m��}묪)y�J�/�LՉp_���
v(�7�j'�%���8[�sH�UA��\��xui�3f�[�����������_Ǧ�G�����{�      ����Q)�QQu:�"�  @e4�Θw������Z��*�s�V��[���ڋ�s*. ��}+��5׿��W\נa����0(���՗�ٻ�"m�v�ho~�Վ"�7Hm�b���J��<�i��Ǒ���wiYڦ*?τ3��U��Қ@         ��3+�7[.iw�u�鵟��o���|����-ػN�S�
�����ߙ��V0_�G�L7t9�V���vkK�n��ܮ���(�V�o���B���:(F���=����)�v���I��ؖ�Q�Wg��c�2��>8^��>���xX_�U�״1kg����|�        ���@��%���#�֓}���n�(� Kv�Mߏ|@�"�*�?L�ٺx�c�Vo@��WP����mP��r��G����w��էۦ매���g�����������F���*l�P~޵@�.{C����sL������+;���;��X��
���	�����W���V��"����|��Uc�� �_�M�����5��i���K���Ȯ�0�        ��"Ѐ:�6c��r���{��`��������k¢�*}�P7b��4T�:�	�>�F�mEu�j���ĪtP�E{cO�k�p�TkK�֍]�ЄN'�k�ao~��X������t+��Ժ��n��.�+��_�&�sW��uDl�󏇴5;�ҹ�"�.���4F�S���|m۶՗g���        �RP�Le��fݣH���d���k�ږ�,ԭh��r�܅>�T0����Y��-OK�K^�*����=�<�n�No��!��Tז�ۨSfݥĬ]u6�i�q���N�d�;��J_����Z4�e]���Jf��D��	h�Rǎ�����ڱcG�����WBBI���)�2$�       �4�ޤ�gh��EB�
���;^�**3f+�8��=��J�UЪ�"�Bݻ�]=��c��TWVglը���>�jue^����V����.s�F�z��}�n�zf�Ǚ��'C'���3����))7��1���_M]B�N��������ӽ��[�9��飋.�Ⱥ������]+        �4x���@EDTo��߸���]��V�kyT\k�}`D�j�ôL8}��VH�>�
u��筶w�����m�ܡ�~������`��K_Պ�D�:��J[g��cb�Xm+^\���\���He�+� MUxx��J�Ѿ}{       ���@����r8�	x5�xa�q
p�l����3�;o�P;!>�厏���z�K~v_��j�:9[�h�?RW딙w�[Y��ݳ����Ե�O��9Ey:e��V8����8Y�����;*5��+O�o}~O���>�:ͺ�]BZU:��'@v�M.7���|���U;�`�L        ���@���k�/��AΕ��j�d��VI��X���@C-E�9u~ۣ���o�դ��j�{�����PFa��MK^Q��۷FϿo�{Z����fZJ�?�a+�`Z{T�mP���{��f#��g > �������6G��Ϳh.�f023�*        hX�@�
��y����R�oP�����p�o����O�]��an�j�mCfa�~�6��\ˎ~M�
�OTd}�=��35�O�NSgg�����*oڂ*̰����mӕ[T������Ҕ�_���u��i���        M��ʥ��� pu�Stu�S�e��ٻt�̻<̰_b�.=��C=���j=�����U��d^���.:%ax���&(V�>I��\{��45?����%�[�s�r��j�@*��g��9����F�        ���˘6�]������]�:mֽJ�MUczn������V���0�K>�:U��]�q���4$��ZT��BU���p-��Ξ�_�ДlU���{�j?���-E�l      ԕ|U�{F�F�H� @�!ЀZK�����ZP�����@��x뾩 P�v	��*0F?�|P�����9&-[��Sc3�K�m�^�u;�J����F�ΰ���0a�s�߰��|Q�y�#:�����      ���a�O����  ��@j�KH+-?�5m�ک��L��X�������+;��	������uP�f��z���K]���~"O�v��*��1[����3�ˮ�:*����)�+��k�*(Z�[Tzl��O��K�}�
r h222���+ h��v����     ���@j��.g����,|V�ه<�楯괄���9zy÷Ti��H��8�C�>�6�Z�nob��^���vk¢�[O�6c�V�oV�ж��]��Y{V�Ә����^���Tfu�V��v���$����-���]=.����_��]o�٪1y�h���󕕕% h�4      4Pcf�ք̂�W�9Y��z+�'+�08��f��*g��vo���V��E��㭿�)i�����U:�G[�jn�jy��w-<d�ay�&�
�i�۠v���-Wx��\��?��F��H��@�옣���Vi{x�l�]2�j�J�"         �)!���i��k�4ȹ��B���*kZ D����mӫu���ˬ@C��N����jTL�
��kx�{�+wo�q4yf�ֵ>�����L�CY���������@�iK�p�2�K�6j��k���{tdl�
������
5��         @SA��8�S�w�ז�ǚ6��}�:Ǯ����h�P�rG���ZGTļ���9��Z.�����U
4|�s�V�'�U�u�n��~۽D����>8�����W$� [��~��<Q�>���z��ד}��ʅ��VcEk߯�{l��[�T��gۜ�	���YYrU�        �(�@XX�Z�j�0'�/��}��X�S�?~��Q>��^���,�}�e�.���բ�"k2�j{�%FWz�76� O�%{�!�I�ϐ�2�/����&�8���S�+oג�*��<�0�`_q��+:�C��gV�
�(8�.��\.�����=���PPP�u?�7@6w��O!        �N��y��Y��4;sS�����ݪ��A�]�۪,T7g�t;[]B����g�.��X�a���%/�ym�V�߄����<վ�L���
�F^Q�<��Is�4�
�<-��/r�tΜ4�g�+�]��؊?^���rU��/ O۳�.>m�u?==]/��B���ڵ�N;�4�~aa�>M~H        �{h@�e�菔��S":k��u�|��:0��	��o�K���D�
ZEl�ک�fݫ<W���en�t��]�uOe�W�?� �_����=/�s�y�k����6-���M��
Ua�O�:�n-9�U9�oA�'�����h���T�7�O-[���h�ª����_�9�u�v`빞ۍ        T��ʳ뿰��K�ߢ�;*<6�᯷ݤ�Ζz�%�	廱��.Z����{B{�q�eW���S�|y:��^�~�O�<�	-,ػV���ߚ]�����?_���?=z��s[�s�N�d�4����D�4���        4P+�m��/���)	õx��zy÷�r�L�H�l�
0!�v�q:2����|�:;�#'E��&�/�/TWv<��}ol��ڕ-�_���IY%Of�z��+�U�2 Z�nѾ�e{j�yj���"}�;�����ms����� oV�0����+        �th@��v ��}Xo�Qg�����imY��U�Ϻ�
5�|�'�O`���l�R� HvQ�|�m���m�d-�y�	�x���Ie�
jPE�T^�o��|�=c1�Ͳ��jNؼy�F�!        �4h@�e��9�ğuu�5*�0����_�o�����^������]��r�M�����j�W�x�|SV�J�dm�V��Z�'ٖS��D���Fs}�c�V�oQ��6�����g���l�D=��C�~f~���rU{�D������=.y��7        P9�3?$͵6��zW�i�`* ��M�B8����;�}��<W��j�&
�/�����i��w8�1	�����'W�H+�*3f�>5aB(ϯ�J/����c���hݺ�u�b�c���w�<�-���d���9���Цf-$$D��� O�.�o�����8      4�s�$����ֆ�9�Őr�J�����5��^Ɋ޾�,y�]�tܸ�z'q�<Ua9�%�dR]�o����M��V�����C4 ͜����N� �ӹ\.      (��Z��_�w9]'���0e�hj�b=���/�7WG�,w�,^�T�oP��*���	l�G���ұ����@��f/3��	��|I�?[3S�kdt�r��m�V�1^Q�    ��y���( 4
��  �����k���Q�hxt�R�M���Fi�	�����iHT�2㦽�7;f�bފ��[d�$}�;�E@d��=���
�RzA�<Q�_H���Z�)�Uh0����[�?	    аr�n  �z
]n���HKv��Ȧ�@�b�Rt�]QA6�:�ǂlͽ�,��h������**__���o�2
��Ěϴ,m�Z��.g�MP���y�.���ph������Qf|m�6��g�x�P��
�����I�k3��ǚJ!g���6~/O�" ��Xm���}�*��?�3�       ��K�v�ޟ�1�U�q>vt�b�6E���:KB�~x ��)!��|||�PCC�U���	íۓfܥߒ��x�4�9�-�R����O�-ޙp(�Bۗ;�`��Z��Q��*V?h&�q~�#���k;���7����o=BۖK��՜���t�r�	       �'1�����C�S�!9K�[�� ~���K*;D�?ح�C̟�?��[h�S\��j��r�lT���!	ڔ�T*�`$��]��]�)��B�z��+w|yZb��M��p_א�VU���Ӝ�fL�=C���a�r�Ly�~�ʌ9}��Ծ���iڹ�
��/��Y��        �bvb��&:�PU�En�LW�VT�1��Lez�1�-�eݚ����E/�K�Z��D�� ���R�m���m�o ��*hYA�`W��Z��*(��}�MC'g���?{��v]�q���ܾ��ޥ��ZF�R6
�E�?KEE�% �� E@p� ��L��ZhK���������땎ۗ���y�o��o'�ܵ����T�V$1�n��m{��+�J�by�^E���x�9��eC�TYճ@��DQ�X��k'�=��tI�        �xW��]���׮J3�_'��R�!'ٶ��ŧ�.LŇ�j B�@z�����}���������~[����I[��r���@�i5a�-���[c?��n~A���ܣ�j�������a�B�;��1����^��        ���������vt�Ӵx�og��lWf���o���܏�s���5�	�t�����.�6͙�����z>9~���-uކ�ӄIL[��|f�,�~�ˊ��/���W��k��z)��J$�l��.��:�:מ2-C:b^W       �Į�^�:�X�Έ�ш.^�^�j0ç-e�^�׼��6L1ᆖ�k*>$ٕ���|����a�vh@��Κ��Ͻ���O�x���ǿs���Z���6��HOIȲ%9+��5Aqc�"�	3tTq�+R��zf�͚3���_���/�#�ru�c�]>)uD����릕�Ώy       =������б�F�����z0S�!=��~K����ꡣ��J!j<�m���uG&��ts��k�?���������ͱ�e_&h���膕��/�2�C��=�HJ\B��M%        �ZCy�mH3�.�ƷTx0��֊�UZ�m��z@"Ѐ^�z�BpT{�ڜ����}�6�K�}�/����n��at� �y�̌�y\�w뱭��/�H��F���:�{�;���~�9������^P        D�O*��[��Ѓ�a��;���8<�0(ծ$���C���͵m�����}�9�K�e�Ru����V>��0����O����iA���3��zo�����Ʉ�t��;mb�;*}l�گ�6:
�x��>�        ��h��UX��0�-�=�@CV�]9�6e&��6k���L���&DQ`JE��������yj����۰wg���&��>���Z�����럻��G�Ni�$�~�=��:"$�w��zr�J�s��-���������ti��3'�(�05mt��7W����    "�y�e+�c��c�)%%�ey�"���0$��.u��U�J�O������U�*�g�,  ����ʰ�m2ç��)#A-UR�tK;3����p�=C�r���W9 ,ǊfW�� �������c3'�hC�4,1������f�}��+��4�r�ݚ�ѳ��Uv�M����O�W���\J?�|��yV��?!s��׿�}�]Gֵ�    �ߞ6(--M�̻J#F��x�*��"4��Ʋ:���TӦM��:��VU�=�  �w�������u5����vV�'��/��d��[�:dYUZ��V���N�	��(����������O���v��6�N���*l(�����L��9��9�:{�-�l�Q(MNi���4P�b�P�����/�W��`3��_O�F�;������Vk��-N�>���k	4        "�q#zim��~����_�p����>>�[s?3�%�`�]A�!
���)>>><�gG�1��/i�����ܣ�􎷺��s���y�1Ao����_x{�C]a|];�\�;�Z%�u�u��v�YW��u��n�W��IN�C)�DKȶBN{�~��9Q+�xL�l�������M
�A��˱��Ԝ���v�3Y'dM҂��]�fdR��N��:     r�|>���6��:����_OCC�5�?&s.U�5�C   }f�@������4�
�O*��[c}qەᝎ�`�v�|�Y�0�)n.\�@1�E��,��#�<l���ܭ@��p��c�SǤ��g�^�,���+Y�`��:BL��U��#������O��z�t��Ul�0x`�LI����꜁3�W<h�	R�=�J]3�\ݻ�9=��u�zz��n}{��Ѥ/+%.Q=����v+�p�Г�pH{��k��    "��fSmm�~�a�gFF�<�


�kx�߼ǅ���j������n�����b��9�ʓ<�p  ��Nv�WT\���f�T���s��㴿�E���Ņ	;�N'8�G�� ��h83�e��T�Xե���5E���^���8�Μ{� ŭ����^Tk�2L?�E]xl�E�Ƕ��G���m��]޿iհ�r�5����\�c]?�BK�nw;�b�����O�\��w��gw��Eek;��`�G��ռ�st��sz�\;E����l��f��y�p��}    "Oyy�5>�O��j&�`  @$1�}^�~��I�RZ4z�]���h�s�k#�e�^?��CVrk���i��d�\T$�j��z�RU{��������|Vw�{�K��l�A9s��.>׺������a�:y��N�Mw%�A��+�O��G[�jO��Y�o���bos�z�?L�6��kG��O���Ёi�p��s�a�ei�&��ީ��h���q	�r�jJ�(�q��&�B��iz�xE��^8�D�K��:����        ��6�q�[;+}Z��Sa�_�u>��˺-�����Q��Ǝ���I�o	:��Cξ�Ck��k/�.D(@1a�'�����]xز��~N�nz������iQLn�ӪaFY�^�_�Zk�n׎�"�����éA�օvs�ZژC���o�e�R��w+�L���彤��|G����6��m�c��5��v�ȳ;4�
�O���uv��=       �h3|��m�m2�O�e�>�~E�t}`�Nj�Һ��j�[ck;����􄖐��쐕$e'����rR��r{x
����P޿����v���	_�mk��p�K��~X��`2�.2��uߦ�u�ǭ
�T�T��߭7����[/"�������֖��v��Ƙ�5m����p�B��       nI�����h���	4��I�~+�PQ����D���@�f�n୯�M%�W)Ov�40�fUt0#7��~fRK��T �|�yU���j��r�����[�����oic��6��w�t��/+������C�����z�?m{�
�{�]Js&)�8�q�s��Y+�26y�~:��a�|�q۫       ��r9̅fY���{	|0m.̴�gU���V���� ��ѯ���_�mEj|K�a`�ie�R���[�۬�6B�B��@7�z\��uX%����H���z�y��1�հ�lE2�������E��%+u�����I�(9.A����O�B+o-?h�i%��	?�4��uQES�      =lM>��רaZ�  �������m�����ooqh��/o��G?��}Z�!�����!e&�Vy����� +�`�J�� �
l~A7��wز�i�����ץK~!����33���)W*��x��}fh��t����g�����#T�|+��a�:�+V�ݡQIu�cuԀ���s��z���4��oikm�5/��ֿO�KG������͋     @�0a��?�;�VUT�� Ds�9٭N[]|@g���*��!��Bp^^�Vy���EfRK����6%��O�@�~������48!�e_6���cZx�^M0F/�p��r"��Z�Dw���"�9���=��&_��4���-/�[������n_��x�;����k��t�j�i����u�����iv��N�u�'��G�/     �h�?̰�ֺ��b�uK� �SW�&�P�`Z\����0�>���u��u-�+�is�_5�=x�]Ǵ��J2�����1qr���}X���t*111,ǲӴ%bT{�t�ǿ�k'������su\�D�4V�����3m�^�����������x����M��7�����=��6ڃ�¥:���i��(�=����Nӯ�^����~��z�h�      3X��  �9�--�茩�`.l|�޿���&9W^.{���Z���m�?V4�ƹnM̱+�h�.�+l��7�/��7o-밊�iY`FG꼍�_�R�w���V)q���c�!�m�ܶ�6+�%S���e�����M�{�/�ؤ�~|�VUm��6��J�����Y7w�x�o��V�^      �m�Zj  �c*>�uw|���k��]^G�?3�Ln�A?;ۭ�9�Q��N=��0,�j��#�i�p|�$�=pf��3~��=���z�\gf�x]>�L��C�+E����H�o{M�hy�f=��}}q��A���^�7�?�F_s�����w���WtR9PyS��-�i��     ���0�ЊP ����RF��i�JՍ]>��I>D�F�t߂&=�����"v>�N�!
�����B�dZ4�V���{��i�6��nҒ��g>�oƍ���P�L�D���W�o�sV�Hu����:�`�=�*	��{���0��?n��~~�U]��'랱#      �|]
3�"�  "��k��&�_5��4�`"O�^�>���I�b�J� 
�/����Nԥ�MU�����6��՟��fU�v̹Ak�`��ם�S$��2Ϫ�0#}\��7���ܥ�?���<���t�rغ�����5     @��V��� @��&��.��/������Oe���&!̖���y�����D� J|X��K�����W	(i��7�?���?Пg�P9��7�����F�����Q���S��ޮ�%+�r��ZU�UG�麦�Ȫʭ    D�ө�O?]&LPRR�<���ݫ�ū�DCs�}�����E]�A�Y���ب��254�������Q��� @2���)
sݺ�i�5��`�	<X�u��jM^!HJ"ಜ��K
־4 Q��2��N�{f��V��7L��io^�gfݤ�sg�j_o-S4x�h�~�����y�?��m��lmP�ea�.�Vl�Z]     "���W||��:�(�1�eM�lRE���DCNN�fϞ}Т�c�j�z�C��^�Zj  D�D���:�mW*>���U�,t�٧>����V"�@%�-�Z�`V
8��[�����գ���~>(]�h`�"��Iq�]Zߴ�8oᏂf0��շ�^��z��      "WP��5  bXW+>t|(�����/O\�Gph �ĺ�;����Ӷ�������t����pÏ&~�����~m�ޥh`�uC�\��B�	S���w��>�	Wt�+�    ��ƍ���Tum�J��ZV����I�x�3P�x�a�5j��A3�"�  ��|�ilms�zh	?��!����(����h��E��"�,���M5*j��1�����<���*=0���ڶ��Ju�FE�uE���aB/�.L�__��:�Z^AIPĐ��m&fm=���ɠ�   z���g������z~����
=��6���Zj  �S�n[`H���G���a\\\�u����t��p�c�W�߭Zo`(I��.�W�UT#U��E��h��khn�����݁7,5X"��?�0�P��Ot<��E��%��)Wvy���:E������y������7B~���x%�� b�Y�sT�����m��%L_bc�ȑzi^�|�     a�0C+B  ���Uuuu`��������1c���h�7�Wm�;��h����s��١�&����*��kM�TTk����O�#����d_00,�Z��/�4D���+�
���m.e������)�=@�wa��o�{M�}��/�ؤ�y2,��P�q�C�]��]��{�_����tSS�������ө��k:55U6���     ��0C+B��k��$�.��� b������4�H0#N�
�1&�%}v���l����h��żm�p
�A�!
$$$(==]aa#9�<~��������6�����p���נ��6��uME�h��LlwY��^_Yr��:	=K����e��_�R@,<}������޽{u��v{S�LѼy�i��}f�     \�fhE�!6�8�:�o�C�4 �Le���f���4�%�,����>i�"��w��n�!Õ��6�,�_�eN��Ĝ�5�c����S}�=?\�Gm���sq;��E��]��맒
b�������ܚ�}�RCw�3f�>��-     ��'a�V�  @#� D�J�i{m�F&��,���KUs�.]��?�>+�О�[#s���P�`b��6�o�ޥ?n�oX�%��jw��w�+ ����w;���     ��0C+B  D�8�D�(c*$�s�|�p�Ň-Kq&(��R�7��L~�t�����3��כ>`LT��i���沛V=n����*4�0˒�b]ccc�������8    �KfhE� ��02î�"��X� � D�gw�h�����֒��\��ɺgt��3��Ljw��rf��=��Nϝ���E�k�R�a=�ͮtgr����k�jbYMMM�[�n��'�,     �!���5  ���P�!�4 QhE��x��pزc2�[����Z�o��~<��v�9wб��'������:���w�{F�6,1[N{�?�����u�i�'���z-?���}l�[��}���}��     4"2�ЊP  }*�+�A��	D!X�w�feL8l�1���z.�o���=�e���]?2)W��L���?Q��LօCf6?�&_o-��LJ���U�Ģ��bm��ܱFVO�ҨM��>�k     A�a�V�  @� � D�5U��4��5%�籷�N�nyE�M�r��|k��":���Qg+��>l�c[_��3�	���zGm�      �7�"�ЊP  ��(�a�:]5����I����'�ya;�?oS�N�D�v>��!'hF�8-�جHc�v�4�K��o�6����'gOms����ߺ      VEU���  �4 Q�Z!|q��a4l��c,NȜ��rt���o��ߗ�Y�o��e����Z��*m�
���9�ڭ��f�R      ��2�ЊP  �b�(���H��w눔��-���9�u�a=�?o��@�qR֑�����Ȗ�(R�>N7qQ��^/�X}��!�崷����      B#���5  �(E�!
8�\������L��^��&~���c�kN�T�W�*l��Z�G��sߴk��|��E@�W��;���m.�@�5��ms���]ZU�U      ��3�"�   ���(���԰��%�M���V���	��5а��D�j5*i`���;\z�t���κb�s�G��n�>9��Y�u|�6��
      ��
3�"�   ���(��_����a9V��B�0-'>([�f������<�����0�`K���s~����=��
7��i���Low���k�~6�6�7�<zf��     @x�d���  E4D����z������z�sz��m.�y4�ß��\>([��G���z㒇��SԹo��m
�,wZ���N̚��z�w)��o��V���<�k�vח      ��a�V�  @� � D�����{�kr��Ö}a�I:#�h�U�,,粣����J�N�����a=��M��IYG��Y7idRn��ns�aHB��~]�����_n��      z�"�ЊP  ��(���uǚ?�_'�y�2�ͦgfݤio]������KA}y��O�Kԓ3o�Cf��jkmA��)ݕ�;']�o���6{���X�[������n�γ-���X     @h��0C+B   �h b�{�ş贜�[��n]0?k��j�yBze=��s�O��g�-�������ڮWzh�	|}��������J�ֶ�={=qϑ_m�F��^?\�G      ��e���  �4 1�;�<�eg<"��yزS����ܠ+>���� Tj==�֜���.�7�~V�|�gw��W�������4���3]_v��0�$%�%t�<��S�mR8|u�9��/�������=��     @���0C+B  M���O�a��h͓���k�\~و3T�P�W�!d��p�zq6��|�5�~�VVnђ�ʫ����B���Y!�ԸD%ƹ5,!Gc����#4+c|����r�!�faߣG�:^[���}��      B�0�5  �����h b�o6=�s�ҩ9��\���_T�ݡV<�J�2��?�ͮ��N�T6��l�&����n��m�l�����
t       43��P  �VT���`"�r�4�*+,�ڐR&��B(�������w����Ȥ�6����k`|����>�{�z�ɩ#�H�@�W���'g�@N{�?~M��ˋ����      43t�P  ����@C0h�+�u���a9�o��T����J���Ewh���(͙��:_6Wc��%?ז�������'dNւ��Aݧ�6q��+uӄ��m3a�� �~$      �a�. Ԁ}�{e��3�ə\��Cy��T����Rrrrxfb����:��z��{��p���̌�Zqƣ��������Z�zÄ'���Xp�S���Z[�������봜�:\������%      �a�n Ԁ��Nm�py��Y  ���(���������F�!V�_�Z�-��^<���VjH�K�cGWW�:�
6�mz�#����Dł����!����ڏi+�1���)Wt�ܘ0í��      B�0Cj  �K<>���n6�!� ��[�B'��=����ihBv��j�E�	4<��E���X���%kM+�['~ٺpK�x��P�K������.{�U���I�il�����}�����Ȗ�      �A��5  �!��&���5h�W5z�j�:T�dSU�]E56U4ص�J�SmS��.�� ƭ�ڦ����{��5%md�랔u�5ʛ��߂��v�r-��l]�o�y����J��:1k��y��%	�y6�kKM�v�YcO}i��j�5���pк��Đ�,����S�[�d�=��J������^��������tfF�8]4�$�9��?�꽍�d���R�     @hfB ��9���-\���V�/^U�ʛ��`k���l�����+�1@?����
5�?����s:]�\̿t�i�hUִWU͵ֲ�䠞������5ZP�ZK+6jY�f�ח�j�	�&���tF�њ�3��-1�>n�x�n��%-._�%e��6_e����y�+Y#s��ȱ40����[U�U_Yr��Tm      B�0Cj  D�&�_5�Ry��
$���UT������M�����"�������꥿�����v
��nmo�2�,�&��g������(\�����~`�f�.�%9�q��=MW�:[�-����}�m6��9�����uߦ�t������      �G�!5  ����P��?(�`n��+���E�)�~ƴ7X��Z�1�R];�<����1�W��G������iU}�2�͢e��r���G\���nz뽒U��?��     @�f!B � �i4A��Χ½���B�D��J�t�'��/����a�(�ٽvݵ��Nw���U-����K��߲�Oz|�kz��tJ����Tdx���v�z�`�      Z�P �&|Pq@ �5��ZY�l_H����
��r���l6O��E��Ƕ���e��+��.�M.�-�l��ХK�QAC�"�y�g.�Y/�p��t\����t������q      z�P �[M^N�
�}-�j}-U���|Vp�4���#����Z_w9��`�@ �y���%�ӳnR�;-h��_�R���|Ab�iEq���jǹU���}�������X��>�F     �_f��  ���

�-a��>��Bq�_�y�����%�v{��, ��z��:꭯���ݪ�������~����7fhU�X�u{w���qA��e��z.     ��� �x]	*���5QQ!ڍʰk��4��(`��L�E@8�/թ�oԏ&}E�N�DN{�L�+Q^�[��cC2{�b�����__&      �a�@� �D�W�nl	%��Zn����*�I.�n��R�7�.Q 11Q��K��Kp��$�x�����Ezr捚>`L����N���T��Y���A�j`|��c��5�aţzr�     @�f� �  h<>ioC�A3�OVSl�i�[#�c�Z/��(P�Q��8,���'�Պ�-���o�	_�m�"W7�5��%�c?��7�K�*���ӯ����,�ח=`U�      @�f�@� �C^�T��Wپ@BKP��/U��_� �]���`Sv�M�R�:Ȯ�G��[�&�#�����|�{A�����O��E/�Y��L��Nϝѭ�6�J�Q�T���P$��ԫ5*i`���^[�[V�I��zW      /��P�~��ф��:_�m����B��gJj�V��H��fU\�Hl��6e&ٕ�`*1ح �#�
1��@�.Y]�Mg,�Ig<F�<�k�6`t��Kp����wh�{?PQC�"ɍ����c/��6�M������wy/E|+     �XD�!
j C��-����-aN(���*�֚6�~@�LX!#A�H�k`���Y��tf�	+H�N��) ��T[x�h�.~�~:�
O��t������9�ҩ�oTqc�"�գ��/�^����Mz(�ߺg��U�T#      �a�(B�@�k/����Y��l#���UQ�TQ8��BKhaH�]	N��4 �6�߯�w��욯KG�����&���p�ɩ#5���t�wjS�n�[��'S.�m�lMw���F�myU潨��2     �of�B� �T�il	'���*�98�P��m�e.�	(h_P�n��80�0(ծ$� ��i��m��m�[�(�}��t������J������Wzq�"�[r\���u�.2��u?����[_�3;�V��N      �;��� A���WM�*
-�ʭ�
>��Bm��=&���$e%����m�tV`���j��A�@��_�~l����k�eV��-��D��;������Oiosx����G����&�p���[�ե�jY�f     ��f�� t��B���TP�Se�TZ�RiaoAt_������pB�]���9�-�\H�"� AU�P�k��VE�}ҥm�cZ=\?�B}q�ݼ�q�
�	E�B�+Y�8�j}m�g:m1aBg-�YeM{     ��G�!�j Љ�j��{�Q�}��\�IO�)'�%�`�
���[f9����(�SZ�;,���l
مe�/w����J���P�1(>C��C+l��ЫK���������^�o�=_�ɝ���t�>��ְU�      @�3� B �Q\��M�6X�$�VZ�=dZ��
�-��Z*0 �h���uk���X�=r���p��?���LL�N.{�?nN̚b���|=��o�y���j��?T����B��8S�W���Ǯ�����T�i      �a�F�@�_�H���Iq�L8���i�UU!�ja��!�@C4������
@�=����ڦ玿ê�Б�Ƀ���o��S��{%+�f�2-.[�UU[۬�`��4<1G��՜�:g�L�O��s��}�e��t���L     !3�� `u�Wk
i3K��*(�$ۭ����}a3��*5���JHNN����s0ʲ L;�c�����y���=���M5�3�q����5*o���M[
�N�{@��0jg]����^���      2f�G5 �g�N�=\Y�L0�ӊ
6e%���0�I.�7"x4 ���2���f}q��zd���r�uk��dk�����ǭ��V�A՞:      2f�5 ȯ��r���˪�`�=��ZZ?d'�TY0#5��@��zn�-(]��'^��G�#���c�[�B��y�jc     ��A��#� �{�h�d�MSl�Hl��-�3��JOh��@1wD ®��B���!�r㳺e�%�b�Jp�Cr,S�a~�Jݵ��W�J      �,�@� zτ2��D����Z�
����*���C�@��UW�o.P7�~\����#��	��e��>����H��xKOF^M�      y3`?B ЮC�
	6�����L4a)�Ii�& ����:=��5kd�RuJ�4�͞��cuD�Pk^G�M�T�[��0�S�B��w      ��0C�@?�r�j�`�(�
"3�%�08զDa�_ D����������*Õ���Jt�5��lͫ�4��[���j�/�ZK       :f@�5 �!N���/�`UWHi�nma�� �G�@�+o��      �at�PЯ8l���EV�J�+3Q�N�);�n���[��N!� ��       @Xf@�j �s�?�8�RF�MYI-�sk�&����d0�  ��       @�f@�j ��c���Mް���[+*��
�}Z�
9��	6��+ �@        �3��5 1o�p�&�ص�����ŷLU��}�����
f^F�~i jh�III���
˱^�        X3��5 1�Dn9խ��ը-e�����@$}�"�j���AX�%�@�<�WSX��       a� �e$�t����`�W늼������BKX!;I�wV �Q�9�2���7      @� ̀�#� �4�]:i�� Њ@        �3 d5  Яh        a��  �       �� ̀�!�  @�@�       �k�v�  �y        �B�}�P  1�@C�l]�Z5���_��9l�'�y      �HD�}�P  1�@C��X���v�       D���  �I        �F��P  1�@       �[3 bj   �h        taD<B  �       �.!̀�A� ��@�       �)��:�  �z        "̀�E� ��F�       �.��z�  ��!��kM�Ņ>n@�       �&���  �����;�����{�:�n���tzX���n���h        �0b�  ����~ּy�}u|       ��f@�"�  @��?���m.��l���7p��p8��v{e`��������k����7�'�        ؏0b�  ����:��^sssZ�f``L�S�:����G�].�k���?�7o^�[Qh        X3�� �  @��|>[cc���������=��j����+��⣮�@       �0�Bac�٬ �\>�/������M���_��㏿�p8>{�W6t��       ��3��"�R&Đ��$��% @d�x<���5-&Bz�߯���3�
�|���W^y����K�al�`�Κ��JVj{m�        ��0�=B!���,��K�� },..N)))����B���Ԕ����=��㯺�]힗�`Db���y�5]�P���k�v�r�U�L�j       ?��>���n�f �(������),��x<	�c����:ao91(>C_z�5       ~��Cj*�n }��󻾾~�SO=u�W\�b[��hX\�^_��.�ɞ�Sr�iJ�(��=���h~�J�/Y�w���K       �@;5�������O� ����9�~bb�����A���!�����x[������g�5���D�9A���ЉYS4+c����S�4H�G�U�ζ�X��͢��^[$       @�f :A�!hjkk�~� ��P__o����>m޼y�;��>jԨ/���pXd7����~kz�����7۶����#�;����0�=uV@�#ݕlNɞ�9�1}�9l-�C+8����+ѫK       �:�@j���fUUU��rQ� "�	��هVg8�]w�e�1��_<�f���c��C�خ�~�E]����}h8TES�^�_l#9.A�eN�_�af�x��Up�<Xc       �u��n"�ЩFyT��x%Ͼ�v%:�rڝ����jln
�9�m~y�>�D�*S_�q����K/�_ i�ݗ�f��o~�v�ndU㩷�7|X�N�3'�����Q�(�������i�d��t��xq5t�����nW\N�Re�/�o���d=��_�6�ޞ�,CN�S���c��xuO�/qv��2�:4K}-#+S��h殓NZ�%{�C�z��������(�'��T%gP_r��; N�.����f��Y�~o9ﭔ�xo��[o     D0�M~7���'�Ipm[�����z����iHJ�A�L��6�������Ɨ T�k��~�a���/�������A����fFT��Tf��5Ys��Zcf�x9��bUs�
�˄�ak�iRc����/�dLL��#��ʓ�u�Y�K�\�=�z`e�iB}���-w;y��ʄ	��РsO=W}���鯖Fw��Y����\9<��N��CcǎU\\��̙��dʧ��U��h�5��eJ �q��K�\���     "��aSŕC���nů��N�l���`�����O �E+#h���y����x�9�j+a*1��}�܇��)i�Ғ��ZX�F�J��7��Gm���|����JHH����ƍ�.�F�w�{Wɮ�.�;|�p+Ѐ�1����->>�K�O�2�
4D����     }�P�E�  ��f������qm�k��� ���S�:�CaC�޷�k���<�B       ��5 � �  @��~�NS�;���53,��I�#���hF�8���5��&�
0�W�RJVkkm�        �C�ha  �����9А��̰�ghVFK)�=��z9�����>        �5 � �  @�������|A۟�fK|��w��Ν�9�8
�!	Y:s��V����D�Q�T;�       /B�>�  ���^����s���������K�ac�n=����3�j?1:i�5�o����|-(Y���@�9o���d��k-㗜vM�1����o۬�x?      "��{�  ���;�0p3&��	K�aw}����C�t�;M�eN���):=w��0Vc�[�Qg[�4�ka��]�\�J�j��򛋪 Bn����}*2�oN=�T�2��n�xK�TE�      �j@�E� ����%�Uz9�5�ZVۉc3'������3�š'[�(j�Ђ��ZT��
:,��#� �He}��J>���p8     ��G��a  "^�����Y��0�W�N̚��9�ur֑�6`�r��
8�j��Ł��[N�]1{�.p���iɒ%���ТE����is?��}>�u���B���Q�C��S����cUU��X��Ҵp�������Ņ�����U^^n=֢�"���)}D����f��tyu���� ;;[.��z�������ޭ��y��������M9ή�����xo     �~��of   *�y��P�M��O���0L��N�X׎>W	�5�a;�b]y|���]`6��HMM�ƍ؍M���L���X#99�&oݚ���"jCC��}SS�u�\�7���F��ժ����gn�W��s�1�̕�u��JvG��	4�\��:������kB���z�N���j
������1�i3jkk���X[�y����L"�Pt�f��
�0���u�>�M`�5�z������=0��=p��������`�߭߃�����L*�Oː&w����j}��zo����}oM(M     ���3  5".А�pkF�8�Κl��0��.!����G�l٢Xfkee�5b��F*s��5 �y�fŲ�[k      ��Pba  �J����5;s��dO����1^N{ۧ�__��%+��t�        �C�1�0"�?� h[�&�p|�$��	2��}������5ThA�j+��00�W��C       PbaD�JO��
 Ж��g�;�>oU`8&���m�W�P�w�W轒UV%�Mջ �lv�t@pȴk(++Sii���������&mڴI[�;      ��D=��pO�O�I�Z �Å%�0)u�n�p�a�� D���ӷ������￯�k�*33S&L���Õ�����4��ũ��A���*,,����e�577k�\���     D?B�Z��-Y�YIc���� p���� � D7S�aѢE�      @�B�Q�0��۟��y�e�<�'�
 �",��UU[5�����z�        щP�aD���/�_���g�����Z՜'����.���o��{O�� "QX%�U�        D7B�x��Le�*?�K�H �0���,w��&���W^M�ʚ�
       ��5 bf   ��-А/���pM5�7>e�:�:��3C��_<�߯�JV�{+���[       �[�q3  s�h��?���Gꃲ����w�\gB�0}p�Jw%4���L��s�ש�o�ҊM       �-B��  �Ia	4$:�:6s�5���7�\��zr����M�z�h�
*tb��~�R��u��u�U�       з5��f   f�%�p|�$��N�{��]��\��):.s�5��f�N��}�חY�M��'S.׏&~ES�FjN�4�[�B       ��G�}�0  1-,��	�ì[�*bos]��\4�����[���a����ڧ5o��2Tg�M�       "��a  b^X��t�vc��v�99k�ukZM�Q����^�O�,��SG
       Y5 l3  �/�%А�`ݚ�mIt�59m�5m*/x��6��YWl�f�R       �<�r�  �7�hh�5[��3�\>3c��lkzY��v�S�\c���       D&B�  �+a	4�/�n����-��|�Ԝ��O�/Y��~2\��m���       "�a  ������n�H����W��_���gX�ō�ZR�����6ʺ�S_*       @d#Ԁ�!�  @��@���5ʫ�����zj捺a�z�h���w'�m�u��/�e;�b;��}i��龯��ek[a�P�2�B�އ�,�˔�t���a��2����t�t!ݛ����q�;^%[��W�I�D��؉lɿ�{����:�ȖTI�:����K?�9�*��c�^R,O�S���gZ�;z
       `�p�3  0eMH����������~M�i����֧/үol8�:.�X���jk���7       ��p�3  0�MH��0!����M�{�߫�S���k�Oz�_�/М��w.�ź��wȪ�        ��0f�  ��&,�`�w���T��<�--�m#���^�4�Y឴��sy� �7��\�v	       �}5`�3   Mp��hu�{�0��Dúkӏ       �n�pR�  �[&<�        ��5 -�  �8h(t��}��邲%*�+Ц�}ְ��V       r�C�  �`BWU���/��*}%Ö}}�'tצ��;        �j��   �	4,*��o/���y)�{�n}k�j	u�g�$       @�#� �   �	4|y�Ca�G���{R{�U�_�k���g�_n�K���������       �}��0�  `hp9����k�T_����Z�����m]�����y�U]�t�_v�^��*       ��@�a
"�   NbBgUg�掇S�y�������2�U2�@       L1��� �1��w�ʼE��פ_6�����q���v���k��j^����>2��D���V[�@�ZC]����s���{�≟�U�Jt����n{ �֞z�ؾY��P�~y.��)]�˖hU�U�J��h����腶z��Yu����6!��
ߑ7$�f*1��ǵ-��5��ro�        S��)�0 d�g�_��j����Gh�{�mV`྽�hp$~���V}aɇ�q�;�|���#�m���IZ2#�L�Xq�I��g0h����[ǉO�ɹ7껫�&�m�+[���^��.��>���z��KB@���.�3�����9���       `j"Ԑ�3 ���0�W�}̚7�k��ܽ_��n��b�\�sƅV���􎸮��6$��^�ʳ*?\X�DŞ}m�_��W�;�ߛ������[�j�65��-�m�I�2���2�b�//���x����iB        ���D� lm�o��Z�ak�	��՟W 2���ׇ^�W��Lˊ�h��9#���O���t�y�z��ohAa��n�M�ή_i�%�����������_���ez��o��t�KK?�V�%�&        ["ԐC3 ��]]��
_�|��0���췦S�7Ф�6�H���Kr&��pI��a�S�a$�"ßZ����uA�!wMh���γ��\T~���ޙ�iqQ]�~?����h~]       ��F�!f ��P�+�o8<�����84�q�Ni�v�2�
�kB&�����O�oI�,kJǔ8y�Y       �)�PC#�  Y�k�oh������{pܶ��x�����Cc�����E�K��5�;��Ő        �#Ԑ�3 @Vy�m�"������Y'�?x��E�3���K�g�n�o�ާW:����Uy��Ɗ۵|��c}e�O��5!��?��)�/�        ��PC!�  Y�`�M���>w�T�)Խg�����o����i�u�B�F5�w�j}���n�8ァ륉u�*�Ԣ�Z���[��W��X<>�zLx�҅r;]��W�y��8���S�O���^K�r �IYY�JJJ���UPP �ө��~k
���R__�      ��@�!f ����M?R�@��y��T�-��5\\�̚>0����~+�0���[S*f��on��ꃭ'ݧU��������B���=����=Bn#�  I<���s$>|�Z�J�^{����T\\|�u�pC}}�~�����5      �D���3 @V�'~�}ׯ��{���*W�3.���W茢Yr9�r&^篮<KW\u�����[��t���t�p�3��uv��X}�~s�W���W�����Pl0�z����_���sy5�_��J��]��2�#�z��������&!7h��2ǧM�6t�aa�Й�^�Wn�[�gh2�M���R<�����s���C���U̥Yf���^���L�}-**Rii���<:S������G�X̺4����5�澚)~��<#�'�}�ٳgkٲe�^G~~�/^��{Iݓh0�#�c�<��c����$//O>���]}��ݛvs;�;�BI���of��33����ݓR�"ϭt��n�-      �P�f ����M�[�Q�.еUg��y7���p��V��U�aC�ޔ�x�m�jH���s��K�f&���cVe�t�ܶiX�٥��e_ג�Y����G�?�Bn"Ѐ����F����QYYi��o����+���G�O�H$bx���w��Fq)���<�Qu7����Ϸ _}������=e������!GD����Ztl���3gj���*//ץ�^j�ML8a�Z��7��ݍ��ܪ���Yg�e�����zn     d�!�  �&�Z�^�ɏ18?^�c_�'���	��C/Z�	 ��ҏZ��;�S�^��1��S�k���7u]�9V���6�ت1Z�:w鋛�����.�X�sJjm���@�&�:Ë�9Cܜ�ozVTTh����� wA�P:8�[ŭq�F��}5g�� �d1�M�"n���SvK���Rm�g�����{��
�����Q�h�ϭ��7s;<�����     �B6@� &U�`��,���o��o�`t�Z��m{H�[�k�U%t�6u��<~�LW}�uL��m������r�       @V#�0�3 ����פ�ʗꌢ:y�n�"i���6wh~wߡSڞY���v�/���5�J����=c���q�P����D�       ��5L�3,����������7]�H�Y<����:S���5�;tQ_]�~�|�j�{�.�Ҵ�oX�n׀6$���s�@M����kW�'( �����u�5�����ׇ^J��uWZ�fx�?�mJZf��Ͱ%�B�L���Ni�Ͷ.)_n͛�ā�ت37�8oh~{/e�s�       @N �0��_���L�
��n�j��ts�Ҕ�ؙ�1hp˙���Jw$.홥������u4F�i����4 S��>��{�'U�-ҷVޡ7�TC���۪��'��h�?�������x�պ�j����m�ٟr[^�[��s�|�#�o|e��k��\�I-�6Ǻ�ۦW�I~������P��
��6a�˗��j���k�뇷��@        gj� ��  ;���Sk���_�E����������u��/2��iz[��z_��r����>���[����ms������������g0�2o��X�����f��:�~}z��u����Ĭ�J-,�i�S�����������g�_�-k��{��B����
����3t��V��PlP�\s�b�W�@v"�  ɕK/��sj�8"��@wo����1�u5��      �h��a ��_6�Y�W�E�q�g� ��-�)e?��_V�����dUfXV<G�.��t~q�}j�w�G��9�l�5�2�����~���Ö"*��/ꮰ�Tv�6�k�6tr� I8�R�z�^2      �,��a ��_5��M�뽵�鲊V5�Bw�U����c�:=ռFq��f��}��?�I��µU�XCB�䕫&��
 ��:��k�5�Ďރ)��l�k��v��!�[��s��a&�7������e���,��WkF^��N�u_������7�L�:*3L        9�PCf �������g��T�����=qJ����?��^�+�XC^�	S������x�\.ר�*�������U�l��v�'�n���Q?ޢѨ���c,ϭp8,      �����0Ê�Px[�é��}E{��n���{���K)��5u�v�ݟ���tb�O��߱�n�z��fhZy�ⱸz]!�� `k0&�|�^�~PJ|��$O�9b��'�'�oW�إ{�ԓ`��+ʗ�G�����Cr��J�yF��aϠ�J��P���'��d+(����T�C/�z�8����!�~�����'���S�"Ϩ��<ǘ�[O��a=����ӚlcznaL�v��\q8��_��T�z��V~I�͊    ���P�ip�ne������G�PHSAӁCrǜr:�r���� ��4`l�m^�Ӯ�5�+i���S܎��f���7�oc�� ��TynaL.�T�};3�ؘ}f���͏5     N��S���a&�񸊊�����r���.c�X���U� `2h  ��f͝���Y�{��U}}��ױd�UUUY�Q��    ��D�a�@��x���VՂ��>+�k��gii�
�ڢ����W  ��)��h�[�j��I�_�*<�@  d�+��RK�	4�^�Z�>�����~Ps�̱�޸Z�l     S��Q�ba��|>��������A������2�p2� ��N)����]=�5��#�{�J ��b>P��I����     C�aS4�p��㱪5�h8��E� `9 @�0c9��	4��      ���x�  ��  �Do�ؿ\1�;;;O��     ��P�q3   "�  ��E1��!k���U�±��{�ޝ:�pՑ���dרQ     �+B"�   l�@  6v���H�ߺRnƾ���~i��     �M�Pa  `c        Sޔ5f   6G�        M�Pa  �4        �)j �   ��        ��ӡ�   �h        �9j �   ��        RȩPa  ��4        �FN�3  �,E� �,�
����8���و�9�u�<�<1    �dYj �   ��  ��u[g���%Im�XL��=c^׺�����     ���Pa  ��4  ��ֵ�P��ے�n��&�y]'o     IV�3  ����,�K��ͥzz�K��8�d'�hL�x�e3˪�7�TϜ�" �g١i��ͭ����q��><�x�E�}p��zmV��	     `"eE��0  ���3.�V�l�c���P���i����`<Uu�iF,_�#>�b�&�g�i_g7�     0)lj �   r��l�]�G͕���WD9�3h��4     `j�e��0  �1        8�
5fȸX,����B!M�6MEEE  �@C�p(�����a�G�Qى����L���r)Ϟ!2�lO����H��pXq=��^�7��#�j��     S�-B���������g�>|X�f�RII�  ��!А%b���n�n�喴}v�ڥ-[��N�������0��`|u����EgkѢEi�<��3C�젠�@�]w݈}b}     ��I5f���þ/3�  L,�"���+�Tuuu�.o��e&���#�e��W���w� �Ge�n���tuuiÆ���K�ꦛF����ɼvtj�s�M�XRۚ5k�P�g��y��Y�r�1�9�o߮�[�jKQ�4C     �LJ��0ø1D�t|U�tՈ ��!АC�Ν+;1�F
3 ���a�@��ŋ�QJ|�>QSS���yk2��uuuV ���Xyyyָ����jiiс�3��U>     ��	5fW愽��J����<�	�  `|h�!����Y�GLM6H��n�x��S�aϞ=�     �߄�3L���*M�6��~�T�4!  0���o1寊���q��`Μ9�̙�v���o��     �ո�3dL<�f*[$����DB��Lx*L(cX �4  Y�@C�����	4p@���.L�ݑb     0�J[r8�u�$w j�dq�pML���؟q	5fȨXm������N�D"ڿ�b�cA�=�	4���U����Rk�T{O�O̅ ��h�1��8l�t�����|5�     ��̻��jjj�ys�����v%��7�s�Gv��Pa��s�\��9S���������.�2�s�0C�����91//OaGL  ؝��m�9���eҪΰ�������&�]^�     @���fZ'F��>�Ov���!9
e7	5f7&�c�[��㘶\������z�@  ـ@C�	��h4j�'f�V��`0h�0�q��     ���K���S~~���=��4�AZ�|���i�3���@X;v�@��.�Uy��t�^���z�V'��7Q�R��z�����5�4���(��� �t4���/����JWM��V��=ɍ�7��/�fК��sx�v��03�����=.�b�x�ơF4n>]���aN��VY��Qo��i�7(t�c�Cἱ�fֻ��Knt�C���w��@sc�OB���¼v      {�D"
�B�
4�a�	VvwJ���j�U�Yi��c�Vfko����~V�ϭ���|s�j�y�|�덻���M��w�;�|Ѿ��j9OB�����u�ުג�*�OM��\�C����(3����;��	  �#Аc�tP���i�������L�v����sN�^\q8#�v�LmذAm��������w�j�+�4�,���]}�7g�oʯK��7�]���r�"=\Q��$|>��kG{{��᰼^�     �}��`>�������H��T�5�b�ŘB��A��= 0Eh�!惄�Jn۶M+W��drE&o������#&��q�$1J�S�8c�4�I:����̄o2���۱c�V�X!     `�\��P�	4��nN���j�v�X;Z�
5f   �h�!����'n˖-��X�rM��S�����v��i��ˤY�f%U�0�ֹ�2�������aR��Q�ᬳβ�����O����7ظq��ɤ�jڴc�|>��zv�Һ����y͚�W�X�dIRyF3�d�Y��`^?�ļ~h     �^\.�5��Q��ݚ;w����9�{����V#�3   !АC8��2ͤ�TWW7i����z�yoOj{����k�)�>�h���Im����f�w���֛�����>@�.s`����lR ���]�^���Z�%W_���������_{��Q&�q��1#y<�߭�+�����u�ީEs�'��}�����P����w�9�,���׉'>�t��Aى��     ���d�+�d&3?Y��l�2�@��VVЦ��a�!g����|��iE�!l{�ǆč8bi�5y��-O��������\�O�M�=\�)�z�'� �lF�!K��/������}6��h�u�s���T*I�|m�^i�����E&���0�L�s�>��-Z4a�4�� �����bUWWk<�*�4���NXIƖҐ~�����q�!j����v�t��	     L,S��RU�5m����c&�\R�aKa���v%����vh�����b�kc���{�D0�5�C  h��O�|��ycU%[�~^������J�`��0�L4s?���&��c~g�d���0F�7��>����z�S�lg�����E     5�E:��fX�f�.Oz����W}}�B�#g����I-=�9�����EG�+���Ɏ�P��k��P茉9   [h��������e:X0Z����$����A*���     ���B]�;wX��.MH���Ѩu�Tf8>�`tuuY'M�IƲ�J�����m�����   R Ѐ)��V�`��!��#h�(�&�o���w0     @�2ðv�|o�껓���	4    �h����������bև������~L�L���Ç5�2@��}     O�J��N�\�[   ��rZ[[3��p8����k޼y�H---]߶m�4Q���3�>�0e�s�L��={�ǎ��     @6�x<֐����I�   N��6G��4Hj�8���̦�_ݿQ���uܑ��G�
�]C��j*�J2w?zեM�����?���9��6E:��vD�2�7xy�Z-�[��6莝Һ���Ք���٪PF�9��v���������      Ȉ��:�|>k�	��m����   ��i�v>�o7=�ܸ�)��דRӓɍ�̭��]�.u��x�2������:?�U�wsB���L�o����9ſ�'�"�8*ƥʸ��?��l      Y�=Q]]mM   @�h            �C�       0d��S�oT6Z]t@*��>����   �8        C��Z�n�>G��/�S��>   7h            �C�          ���q��q)�ؘn7��-04        �8�3�P6r�%W�}w8�|  ���LK��)�hppph
��
�BC�Y~�C�n��=�r��%.�������Vg��So��@       `����ھrX���Kv����T�_7����7g�  ���<�5��F500`���ba����
��f�1�6g�
7��:��R��GM�E�)3�@          `Js�\����TZZ���#�[A���~k2�@���`*8�EK�I���S\�]A5:����M\��x�?xN0����|��c@�          ���xR+�g��S�Rw���*q�U�)T��X~Wވ�7�����x&�p4�`&r0a�)�*�~k:�H���1�������m�x|sb�fڐ�_{�w�)h           ����֤H��Ӝ�����i��B�U�메ב�p��!,�����"f؊��f�
3�B!�ʃ�p8LzbU�r��~��?���D�ZnH\]�X��O|�m�          ����;Ԗ���v�����o�5��Ti�o�jܥr$~Rq�\*,,���c����`�����n�p8f'.f'.o1�#����zp0A�Ĵ���v�m�ui�!�           �q��i_�՚���C�N��y*��b_����)��q��)*vW�!����>��Tr0CX�`��ᘕ���Tr�B���oG��k�i�[�Ul��;���4           0
�XH�C��x�r�R_����j��Vg�jT�&��v��M�f���h4ڟ�`�
9-w$$.�xk�KrHL&�/q�!�x},���x޸����#4        ��Qu�����p�}�v�  0�#���L`�u�KQ�)��L��_��%����Ga�ۻ\������㇫�F�၁�`oo�?x�����(�z+�0/q1/qy���4�1�UJ\#���X�z~~�+����B        C��ZӉ���~U�U�5��������%)�8{" ���[_u߀:�&1m�ۺ������8/���y����KJJ�����u8Α֑��JKK���x<����?����������8�#NJ���ў���=�ܳ���wMSSӖ����HAA��<��@�e  �A>�Os��UMM���ʔ��o�Xo|L����rU���jooWCC�ڔ��L      ����k���sf
 `3yO5���z���$1%l޼ٚ&����!3SRR";ikk;7q�6�2  d�x$6��k��m��&SZj,^ػV�v�P         v@� �l�"j�1�5�`乽        ��y�Bf=�裵�=�������rS�ЭX��     �U�`��Vkߩݲ���jy�K���a�TT/   d�8+z�M��:���}s�W�      WT����w��V�U�]7��� �   ��4            �!�            l�@C)ku�/ޟ���!9��X�Ȕ�G.9�=�+�	��+�t)H���82���1N9�u{�S�z9         �@C�pƤ��y�}�Ѵ}v3$���$Ν;W�E�z���0����ez�����^gFz�)--�ʋ�ҿ���\V�+RM�?��a��         ���,�9@�t:�MF:�f��p��g,�^c�}qGr�5�?�\Ue5�k�ܱW�|��c^WKq?�        �mp� �,�nv�֩3Œ�        �f        Cz��H�e�W�굲�a���A   �h����j�ʕi{��׫��Sv�p�B�\������� �CgW爯1���jjj��̚5K���)�y<��     �M�;�����9��]y�,�   r��,sĵd����i�lڴI/�����nPaaa��ܜ��� L��sg�/J�܄��x�	��5�\�3f�]��ż�l         ���l�,X����]���v�Z�Eqq�.��b9��}�� {����ʥg�]^WW�g�}Vv�t:u�e���������(	        ��4�s0�N/^<b�@v)++���@@v`��)�         ��F�!��{v:ظp�B�-ӧO��k̢E�     2oe�Z�X9��^��}�}�j�놵���֌  ��B�!���`�xW��:��P�ܦ��Kr֤?S;�iG~� �;UD�9s�     @�9?�xvV^u�S�K�y   �:9���@vQ^^>��/n�i�Z�5?g�}�ßN��@k��i�[ N����        ��E�!������n��^�n#����<gj�.�1��\         �<9fppPv�F���pP����2S%!_�9ӂ�KU1�"e?�˩�ÿ�>M�p*vy�1b��         ��4�`0(;0a���~ΠN��׷�3��Tx��ߥe˖��gC���y�N\�!�.���v         �h�1v	4mmm�={��m�y��C{{���ݫ9s���t&ukiiѦ}ۥ��LP�.��5         ��@C1U�t��&,аg�}�{ߓ��See�JJJ�pGGG�����W�x�_% ��n�1�{�     @f*��3�lrFR�{�i�a4  0zrHoo��a�|�زe�.���	�f(����	@�j(va^cn��k�     �9[
Z���k�#��y�fu��   r�����,;ٽ{�U�>??_ F�aU�[�E~���Z�f͚���rkygg�նs�N�?/�ϛ��2�cBCva~MMM���         r��lᐜn�b�X�.�����NZ�[5kf]��<���.SZ4�������\�t:5xn4c����F|�ihl��f�1�m-���N�ܛ�O��$        @V"А%����/K�#t2��%[�U�ץ6����7i�I:��5��}'�g         d%         �����  ��F�i�'N�        d��xT  ٧��3�n�       ����3�ή����ݲ��u.SUcͰ�vwP?�|]   �.        C�1�J"y�FO�}tD'|_�cn��M�l[~��܁���f&�{��k��=�m���P�f�����(���ꇮ�D�tf�:�74�ە\�`��tM��tj���   &�     pZ|�1��
��>}�C��0�����M�J�q 0�E}zw�)���BI��k��"R0��:cR�ay�.�=�߀#�h�,H��o��@�9}5Ve��@�  0�4     ���ǵo�UVVjf�M�6-i�ξ�O      cB�           ��     pzG.��֯_��K����\�`PZwp�T.     �1!�      N��H��}�Q=��cI�.�     0f        #������խx<��Ͻڔ��������ߦD�M��K��WkF�N��D��G����j��yr�\
����
�q~L   ��ˊڢ�e�H�W       ���QxHk�������Aݳ�kO88-q3�C�������m�L�_w�Wuu���  `<�R�!���^�        ��?Qe���#���b�c���t:UVV���.E�Q�2�ۭ��"+�   0r       0"W8u{OO�u@�9k��0�SRR���^��a�"�ϧ�����{,;�/   {h�r��^����<�����;3���ϼP/;7�����o��ǀ      ��)F�-,,�.c�&@ii�B�Фm�D&�`��A�k��8eU�(�  0�4d��h��Ϙ��v��ŪqkF�s�5�m�x�O�
      �cڛ���`�zhoo��{<�'�+oj���W�1�������a�@	  �Mr��ŋ3���ӧ�v���	˖-Smm��A�\7o����ZZZ�3ܘ�C       N�v���@v`����H�7o�Z��� ;  @� А�L*�$���̕�:Z>�V��>��X�B��~{ڮZ�@��p���L�v�ߓ��p:2���	c0.��@���M   @����We��<\_ѣ~WT�|��x0���{��S�?sB�V���OѨ=^�������B  @���O:ƔV3��R� ;�u�<^��:�������'m_*�~5tL�����W�   S����taK��ݞ����q0s���P���v�Vv*���<2hΜ9V5Ü ��۫Xl�!���L�V��	   r��2f0Lɶ\�����U�~�n��f�w�y�6mZR3�Jcc��u�T�j���;r�ñ���0_B�/$     �=�f0�gvs��.r��0����n�/q�81   �h�A---_gww�UJ�xk����<͘1cX��0_,\�P���	>!ꂋ.��W_=t�|y���ft���[o���eB?�C0:�9i�3� �dx���y�n�Ts���Ԧ�}�q$~.�X���ղ��*������HP-��еW�kz�����O�:�U�w'�u��   �h�A;w���:��뭒rv�/*ԊK���B�����rھ-�nȌ�˖���2��^Pkk�*E� ǥ�^��f�Xj�`�>lM  ���|��E_�׷��6m�@4R;��N?=�s:�lq�>��R����x�+�Ěo�=���NQ�}�LeG  �\g�����o��w^�Nҙ����SGGGF����k�ڵIm=�i�&MKUD�W�����.����4̞=[   �^���,�XC�jF^�V_�oVE�?��գ�^Ԗ�:�U4�Bw������z_��zw�Ez��o��?��±�     ##А�q�^�uE��[s�����t������W
@�M/��/���W�0C`dREE�   �EbGB�f���|�3�;w�5��a�����qM�
�4�.��h����H����Z���_��~Ә�r�s�����?ח�ު�.�K+��P��    ��@C��z&oۑI�6�˚�,PQЭ6��C�-G{�j����oW�"�8�9x�   � �׫���0�������R�O���s��)�-���[G3����G�]����� �     �@�!��qn�B�|��ؐr93?|�9�&vl������y[�z�m���3������   L�wĖi���0]��z���SZϊ���l�58ҫj�rY4�._;�]�����q�t��K��r8����yF����\    ���,�V���\曤���;����Օ��?�   ��ֽ\�<�*k���Om�بX,6��|��i�G��o<�6�Z���q���E�:�Զ���x��o�%��������#���6���m{���y��"Ѐ��ڣ;�C�/ѫ�N����]eޢ��v    pr  �%����)��ܷo����~�   0���BUTT����Nd��Ȅp�C���͚D��`�0��f�n��_�.]( �}ף�m��z�o�g���/ks�~u�{�3���i:�t�5��-��j_�Y|^    ��#�  ��6�B-�*�ƣZ{}8�[��v�Dy�c�	�"  @j�t;�׫��/ү�}:g��3<���]j���ʮ�C�a����|^�Ͻ��F��k�����k=    'G� 0&O�6��A���o�)�v   �ROO�)�n``@S�y���<�ѕ�0��}��F��MZ��mzo���<--��2o��=��S�@�6v��o_�ͯ[UB     �C�    �,��ݭÇ��m���5k�,M%�����g�dM    ��!�     @�y�O/��G�85UL0�T<��z��ǭ�<�t�      l�@  @p8r�FW r�y=���U�k�i����ݚ���     �N4   d���2k �xae��
�\1�)=�q)vd���K   �������%�ۭ��
�   �ǻ'     ����1i�'���;�l   a�{�����ӣ�Rq
  `4d��K���Im��[�����n���E:k�⤶_���W��       H��ٙt}``@�`P~�_   Y��Lݼ䪤���z��ƌn����K.Hj۸z�       H��r��   �h�AK�.��O?��uVWW       0:ӧOWww���������   F�@C�����:���d73��t����|II�>���[�Ѩw�}K N߹k�j�m=��!�+�c?ƣq������J�qA@   ��H�{�gެ;�S��3���m�tצkK�~c����+K?��]�Y��-m�.=���>��Gj8, S���ѢE����/��M�  �h�A捱y�|4���u�Mw$�6X�_|�


�������jeG���&|�+V��h   ��{�m�kɇ���8�t��:��O�@�E�X��w香�]��+�_ιN�/�������M�x|X[,S{{���hR��~5���N4��澙`�Q�CQg\   �i����Y�]����H�����rY8V$��:3�>     &Z��P���}����5����7U�-�?/��u �,��7�?�un�"+̰��A�\{��v�Ҝ�j}w����ʳ���o�����P�T�8��B���N�p���R �|B��岖g;s���&�`�~�_,�$*  ��2遆���k��b¶�=tH��$�S��OG__���'.x��fϙ��]7g<���ε�^+�כ��^   ��ZV<G>�G���z��KV[�`�
7\6}�.�8S�X�]z��k�c]b��K>��ݪ�C�b���7}�t577[�J��P��fG���&�`.s�����ڪ��k��#!��   �Ӥ�y�w���::d�Q���>���"q|ɳ�L��;�+ [�wK��C��O8/�v���.H|�tLli�k�y��*+�ڶnݪ����m��>��%}�����v='   �T��WY��ޖ��G���N��30�1e>����jukw_��|���L�j8~�	s�߄r��քL�  `"h�r���#�$�����Y&=��s:p�@R[O�MZ��s�A�����_��,X���J���Z�hS�b�Νj,JW	�
�~�J���y׻ޥe˖��g�`�׵&�_�m�̙4��r���    �(p�Y�����e}�~y�|M���w���4~�2�) ��RCG���%Ǒ�j��n�P�����o�0ԉR�}�c���/�:O������5��Ah<������m  ��ç�,��ԣ/>���k׮������W����rn&�a�a�y�#{l۽C�����˕-
3������     �T��z��i��i)�W���.K��g���i��?5^��H��~���z�|����t-�e=���#�/�=3t}�@�>�z~�m�[����:��nm_���3��m��g���-�O�;lQH   ㍣�Y.3��<�-^�7��3�  ��򫋿���`R��J{
��m�������ݿ����L��9���:�9ղ/m�_O4�. �|  &��,���]g��;��N���7���G�ر�a��z+; F0���29|   p�e�s�.;�tᰶ�[�HǔhO��9*ղrc�   �hh�r�f�H�'�L�Fq�o�"��z{{�ǭ��g�:���=J����et}���   2��O�/��v'Vs ��¦�[���    N�@ �̑�B\���z����?�Auuu*++��wuu����
4���5隚��I;v����<�   �L	�
N@��!k�T��!�d����z���?R�Y����\������^97�x��&o_�m7{������6�?�d�  �d"�  6g�4lݺuX����dx��5M�(��j�3�D&�'���<�b߱��r     �!GD[�GW�rw��Q�k��Z����Qo�8��&   �!�  ������Oh<#���K� �E�ux��_6 �'���{J<����h��a�n�y��v�{��xV���z��K��֟�7T.)����KO{=��.Q�'���m����ٻ������_I����I�E2�d��	��)���G)e�}J'���B�SvK�(�P�e%�!	I����I����4�N�Ķ$GV$����"��ܫ+s,K:��;KWi��Z,J��S��e��ۛ���џ�?�$?D%�Uza�Gzp��rz\�Oeg+kԨ��M���s����r�VVo   ���@  @�e�s�  ��ѩ*:�e�Q�X,���}g��׏�����C��Y��t�'?�۳�0k��6L������X����*�p|�T-:����t�����~9�{�w�ջogD%�îѨ���Ѫ�՟�?^��8���U��m��	4    �     0 ��1�,<���N�m���1߼�w_ԓ���A���:c�3����EK�����aT��Ǯ��gE��I����_���)ZfV�xf����C�П��K[�    ��     0 LJa^~Z��i���54&]�+���uϚ�
��uѲ{��[�in��Ҥ��*j�Զ��N���:RQ�H=���-�]s�1��u����ޫ3�h     h      BfT��Z�U���i�)�3���
>�~Gc�9�<<v���}*��x��s��S�|�i�G�����S    �#     `@0��g�����	��ʍ��W�R�t{���}*�f�o�ѧ���Wmگ}uk�2��S    �     `@��X���hMN�u�;�uF����fՆ�5���&-*A[�tŨ�q��c���6��nL�������-��u�����Ʃ��F    0��n544�Kccc�׷o�^���     ���YE�y�Č��h��U�R��'_nF�������N�"�thB���Е��t��S�����i�c�t��󾷋���~z�٭�s�	    �I[[�>����F�;���}555f��'�����4     �ai��V�3�8��Os��f���ݦ߬~����8�<���5�����a�ٺd�ɺx�I�x$�Ţ��*=�����_=�4�>   �`�m(���V.��3�     0`\�����@?Q�1�P�K���]����k{�U�R�E>�lxc������_F�*��t0���:�_��S��YG���oE�f�⫿�Ә�-!"�l��&W[���W�jӂ֧��]�V�   �P�6�'�б�c����     0`�n[�ws�樏n���bס�)Ay�Uie���4*[���/�ڮ��P��/�'��>���ZE�   }/+%,3gΜ��F۶���b,9 k�G���z,�~�d���n�X�Y,���(�[��|��g)fT�ޛV, ߍ����w{���b�΄���m�016A&�׋ӷ   @p���(333(�e��&����A�S
���   �zJ�����M��WF����n4�_;��q���b/,n�ǥ)����P+���%F+�9^ B����0|�1t}�)�He)I    ��f�):::8fe�y ���^��K  �F�/��B999*//�o�����n�5N�����~��n�	t����;N5Oh�c���@��h߶�`ʉp�c��i	���������d�E��t��p���D��:虥��X��k'   z���uϔ+���/���?n~U��n�p��5���~��/z�h�    ���[���Taa�����n��M�>��v���� C�bC����|�v ����Ыm�����innVkk����r���ln=��O�~��fj�@k�H���p��7�j�v�t[�N-*��     Wbd�F�e��]����ZZTb��TB$�J  �P�q�F�y�栽�F��G}T���B�Y,�4�����N���w�y猳�:��@Cذ��KzJ��X�\-�$..�ې�QE�(��k{�-1�����G��oZZ{~�1�v=�P:��cD7���}F�   ��s;?�k���]�+�>k#tܚ������5:}�r   @pc����_ac�⡇"�`�ej��ۯ���lFyÄ��6��>��n��O֭[�Pr�)�����l��% ��mQ��1EEE�|Q��c�QFFF����V   ���nSK+����b.    ��������o��T�jFtt�5Ţ�;N���ʕ+UPP�PaTM������������o�i�>�n������͛J�9����w{���R�r        �dŊ~o3g��O]L��5j�B�!��c��@%E�i��Ce�H��HUVu���n���
'cǎ5���n����TSScVL�J�v,Æ3�Cej�����   @O"bu���tJ�L���d{�����X�Eek��甆�V����S��ѧ넌�;H	���n�ז�B�_�B����j   @+--�{�3����cp�n���܇�������G����=SV�ig��������iii����5iҤ.�Y,嬹W+];�r\V�U�Raa�B��	   ���i��朻4(*��z�n��9C��p�.��z�h� o.�>Q�~�blQ��}�Єl�5�(�2�"�����z�    ��ތ�c'�;�%�@C?bn) �v�+���п�RҐ�   �Fvl��=�%E�齒�zv�ZS�ݬ��I�#u��������;tԢ�Z� 4z0'}�^8�W���Z���?���<5:��~63e��u�N4]�{�&��6W    ���~�(I*����@�bL�*x�  @o�9�Rs���_=��7�������V���p��y�-�o�5:��_
���ּ�������Q�\����z)o����t�n�~��	    �#��τ�`�Q^%&&F ��P��N`^*   �)���f���3������!�ͩ��SU�\%xg�ق��!�j��6:.K��&�o��z����/�}���O�O��Yy�"##�֧,��    �������NTB�]�T\]&Kn�/�6�M��   �̈́��J��Ջy����]��ϳR�面e�wA;���n��t�3G��7/_�[赭`0*5<0��:$>ˬ��v{�����wY   @�!���455)�\.����)z �y��=_j=��R�BFss�BE(   1�l��f�O���z��!�ovx*��닠<V��N�������O���O�4�f�;_�
R�j�8E�    �h�g*������) �G(��TWWk��X  ��#�>˻�����խ��e�=^�M���V��B`ƆĈ8�=ն��Y��O%E�Ɣ��`���ק3    !�@C?�p8*���4 �L(��jҤI   |e�����������2/�V�>Aעl�r��������{�v     ��Dޏ�����`�ƍ5}�t�?��+�bÆ:��S        ���@C?RVV�Pb6��nY�V��ͪ��W����S]]�   �c�i���M��,     �4���b.�������`3�E%��m�5t���Ǟ^C� A(���mۦ�3gv{��B�
   {���T����vͮV]ir���O���   �<��t��q��pc	�qz:��x{��@h����׊�����&[�v�nS(�k�B�:���+{^�o� ��[�ТM���?��L�B�5�E}�O6�v{�.w�   �����\�@�%�s   00UVV�Zp:�����}ۨ�m���������mCKKK������}L�0*z��/�O�!\��<ײX���
)��/�S ��\���5�^c�Vj   ����X58���$�ߒ#�U���    �GO�
\.�l�='��*�?��m��]���P�     0 \�}�~?�*�[�\�-ջ%���l'�9VǕe�֤��.�wg ʝ�.�yC���%z�x�>)�JmL'P#��֧���i��(   J4     �ay�&}V����KG�5�5�_�B�.\��������1EYAy�����h0�ϔ�Q�~�ٚ?�<��Ԛa����hA�*5����#��֧V���ܨ   @H!�      �55�uޒ�c�����:3�(�=d�.v�\��Un�k�����w�����RJJJp,ª�탒��b���A3t�7��Q��a���V띢ef����Z�_LLL���E    B�  �a�x��ˢ&O��+������H�L!���d��  �@�1�l,ׯzD��&��cꀇ�]o.�v鵂Oͳ��*�&22R���Ay,���:T�6���X�mv�>Yg����do��'f�73�/�����P���	V���D   j4  ��ؖ�Y������w����ߣ�  ��cTfX\��\~��%�s��s��;'^j.����������RQS���4�Z��t���t�_��̹C����~��)ט��mf���-����, �EZ#t|�a]���nS��B���>��f����	�>G��n�TyK����4��Զ5�����x���x�b��-��    �  |��q+--M�������R54�n�q���f���k-  x�PVkB������duݚ���g�7�ZU�g(��gL���]�QPJ��[��lW�P��E�1-���f��;H�>\g9J?{�>)��@��w`�gk���,�?}g���T�  ��IDAT�k�eza�G�u�>,I�qZp�}=�1^���ݿ����ݶ�0�D�;�j������w����~��n���D�ǳ��uy����  @�!�  �7Z#=���~f��5���������O\\���.Y�)W�в���˗�  �g�ڒt]��]����/�1�|���˧+��_���%z>}���G6�)uc��篳���2�'��놲#�l����Z�
V�"�Q�����\�쉻���e�����7�%;6C-u�MaS�J����F�#��jOА�4�v�:%s��}�+�Z�ެ�O�A7�9Ǽm�~�������~�)Z���<��6x�N��4��'U���i��do�   @�"�  @7233�#G���n  �~����gV��V��'����o�g�u����\G���qS��q���殉��3|V��˗߯�%��SI�:�b�>�bMJ�����_x��\�W
2*Bܷ�  �"�  @7bbb�			  @�9o�s��_����,��8����'������{%��Ɣg|v�rO^����|ĩ����[&|߼��z����-jt6�c��;�?gVw�����P�Q����   �  ����ԫ��   z2��53e���}X�R@W��f��O�E�F�cT�YZ�A��Ҹ�a��E���C�gNO��xtՊ�3���/��aǚ�_׍>S�l|Qխ=O+  p�zs�����j�L�  �QUUի�v��!��ô   !���V/�}��v~�]�R��]mzb��7��ѯ|����`.�J��|����6I�q:w�s�Ge��S���~���#[��sG�Bq���`�q�[�  �K�������k���f���
}f#�  ��JOoxG6����ب�s<��S�[�#��[�my  ����]T�Z�kG���=O�ǜg�Ml�7�d��~��y������]�.3K�=��s��,�\N�K�@2&~�yi����F��촉fu�{%+|�׻{M�rL�d  ��{�Z�d�_۬Y�FG}��g^!�  �7<V�ׇR�w�i�,���#��D>�   �9�_+��\�c3���'��g�ə?����@o-5�KW	�EM[����_s��8R�����G��3��Rqs�^��DO�x__��
��f���Qi��˫6���4��O���fm�v��W�R�¦
�Iׄ��ݶ;m��J��y����*r  Гٳgk���ڴi�����������H!�<ϖ��?h      N��\�mzEl~M�d�ԕ#���Ǜ���v�mo�/��#�ǘ;�n��:��F��U�S�k�?t�9�r�<�8�\�{�>�X��7�b�f����>e��"�jW�=޼n��4"v�YAᎉ�����Ӗ7v�O��	�2%��*Z��@C�����	Sͥ'e-5  �W��_����[UTT��6�����{t�m�)"��� ���Y�3�8��O�c�8�\����+O4��   ���q����b�r�Ǟ����6��^0�JJLL�cE��?k�f��>fTy9�cs1*�<2��;t��h�G������֧�.��}�%��O��{6���>ݽ�n��t�ۿiX�<_Wy��u���U��V~�J
  �UZZ�x�=��sZ�h���ڼn�e��t�M���5j�(3����x<���y��y�y�Wc�#� �����     4�G��a��Q��g{<Ҋ�-��J=u��{sP��ӠP������l��)I���nӚ�m��r=�A�S��o�_3B<MZ\�NO��G�*7v�ߘ��Cbd�_�N��3/�Z�m�f�b��  @�����n�e�]f����U__���F544��q۸4��kkku�w������d�zRR����v���ƨa�3�s89f�Ţ����iii1fE4�����p�\f���3f��뮻.g޼y���G� ��F����+���c�*zXr�m���*   �f��յ���E�OTBD�9���^5�v4��ۤ=�Y���(��if�:g���Y��v��P<��}���
�[���}*Tݺ��~�?}n_�T�����a��e�Ԉ�L�z��B   ������3g�����;�~�X:�����fUWW����������7�l��>  %�4b�ۼ>v�!��?���]:��^   �Ș���'�Q�kL����w��鯹��G���r�?�'d늑�t��S48:�<�ٝ���>��z���nIņ�׍*8�ص���L�{��%��  �)�RRR��_{�!��CUUU�A���D�2%F�#�  ��ݢ�|s*"�9R   @������#o��b�����M/���OT�L�O<�O�DwO�\.�[��w~�w��������6k}�NMJi��t�_��l��U#O�}���e  ���C>���
���{��*a\�0�     0 $Gƛa���:E����!g��7����m{K��R�	�eIs�Y����/2on_���+Y.`�xh��۬�*)2N��|�~����z�.1׼�Q�j}U�+   �/::�\�������)2Ve���r����g���@@[�U     �W��6E�zmgi�hk]���=%�J��JrgU��<������*1aO�G��6u=�B|e�\����r9�����n�+Wbt�XZ��?>F���\�fO4_}X�R@O��L��WiQ	�z��#O5���?�\�r��O[��e��I#����e�X�p��Տ	   �w Sd���v
>xCt\�m��r�ʅ~����h|q�� � �{�=��ڶm�F�-���Ӆ��Z��#�	   >�z3_��/
zb|�_[���>S�O�
��t�n�����ç}v������(�g�O�ṝ굂O�ޮ�e8|��<��7<��v��f�1-�E�~�E'�Qc������̬��������)(��s�mVΉ�F����U+�ƺ��}��Õ�=$d��	   8�ݮ��Ts�h0�{/˗/O}��lϔ �N���[����7����+))I�C���fz�n�M:^�ʠ*��
뾾a�(���'?��>2�����&  0�y��+++�k�!\a�����w�ZZ	' p��QH�4��E?�3��Lgd��M3���l,��|PKWy��	S�ś?n~��W  �`�?Sd�=MFnnn|w�	4  �d$䊊�̥�;|{�J�t�����jRM�K���zԷ��î���Q�u���Nn�x�����}n��r��X|���''<�)I��m��o�6��q��͡���;����eYK���*U�\���j5W��3<�|Y1����y5��
7��~q����1�]���z��{&_e�E�Ee�u�һ5y<�'��a�����G�j�=�����6�����No슫S�ͩp2>![W�:M���{%��2Zb�֧��W�m��kv�������z?���3ߦ�2�����ˬ���~����5f��w�������|��8\ͻ��������1   B�  �Vy��Uc�a��ս�Mrr�9U�!**J[78PF��{�|e���h�ݯ����h���~Ӂ��q����@lm(h_
����K�,�ڝf0"%��Lbh��s����ZQ�Y�bT�`�1�:�����?�+�c�;��!C��g#�#��d3s��8h��}��:G����O�7��	�v<�?�m֎�Z�:�5�̬#�>ur�t����o&V��O=4e�
��L�SB��ˇ��O�s̥���=   �. �/m��t�5�o��7�QMM���9餓t�Y{�R}z������`"��a&�:�\���jњ��ZY�E+����k��(�@b�X�Č�:꣛�y���#�oX���5477�U�Q3LLa�9鈹�l��P�K/�}��v.|cT ��N(PV�B��i�tu{��n��f����oY�F�O����7F ,h}�os�    z�@  �4hP�Ç �
cP|v�Ds�`�}P�R�'�_�s��w�R�釣����V�;w���u� OBD���}�9��Qiv�7^g4_�k�	�1*��=j_�D�^�!3:E��8���Kt��P�y��ڼ�bcc�֧d!�    �  ����7�v� ��q�����q�ӓ�S�L�ص@��6��~?�*�Y�X��U
U���#��)c����~�y�Q�ea�*s>����6�� � _�N4��S�9Z��5�Z�Z��z����m.6�f     �h  `MMM�ڮ��A .�#�Ͳ�Ʋ��@m}C��x�_VmH��ӽS��+��Pu��K52.S ��1�����5.a�y{mM�����^�[����+t�<K��.~��o�uʊN5Á���}��������sů�_$�%��I    @8 �  �>***z�ݶm�4u�Tx���~~���YlJ��U��f�'F�)����$s�$;6C�Q)晟�d�=1c�y��my]�����c���Äח�<EO�x_�U�(�tT�����@׌�7�5���\�-�_��p �Ho��^S�]q�9�     p4  �/��t�K�u�G�xVe����V�s� �D�``XW��,+FY�᱃4>a�907!q��J�`^���Cb��S�ǜ�V=��J�+�5:��Q�j�3���!��gܤ~$�ǥP�q\vB*��֘����3 �c����d��c���EK�ܮ�A�Js�	�_��ju;5-�}~�Cz5�=�s��T�    ��h �`q�� 7sƥ�"����n��}h��L��������~
T�5{��O �������Rsy�d���Fe��iuj�L�=�h�����7X�{�^��X7�zL��u
e?^��Niޱ���MI��c�Ӄ[^W��x�I:!�{uc��U�h�	@�[�\������:R׎>C��>N��>^��Uz-�=��C�xtۿ�B�B}g������~e,y�2�3�c�5��    �� �����%������:����N/-���.  �V��0�06���>i����Su��S��ҫ}^�}�O9T�.�ӬB�v9J��/��S�����I�������w�Rrd�8�>���-�iS}� �&W�YU�X�'d��Q�ҥ#暁'civ��ӻ�JVYK� o�[�����6��S��>^��=���������"%DĪ��    �w  g��][l^>|�bcc�mk��� �nc]�~���X��.v��x�9o����%'=��/�W�)^�Pe�_6�sp�'�`҃S�����N��&_�Sؤ#� ����Ͽ���zy�i���9Z�����>.[��w-���ͩ* o�Un4��V?����2��ə�ͩ���~M�V�;��EK��v
    �3F�   �~̘�ॼE��W���?L�F����a� �u��:k�m���K���)>:��^�������2+e��;�L��Sj8\-�w\���2���T�u�Q�kn�s�)[��<#�WF���J F����Oҕ#��̬�������>    �g   ���q�o����_�Y?շ���vk�j���/�E�&��Eek���1h��c�o�a^�w���j���e�X��}�h��*Z" �cTO{x�zd�ul�ds� ��PzoK}��Z����YG�}��v    �� �e����&9�NED����ڪ��� �^QS����6�9�Rs
�G���c~�)� d畿y�:=�%G����8[�g�~G�l|I�v��tx�^�5�Z��5O���i��iy���w�g��{`+ �%�.4Bj���>    �h@�8vU���$�ׇ����&u����/��V���K?.��f^?򸣕��u��({�.�yTng> �Y�|�x�bm۶M�G�VFF�ٿ���UVV���\��ޟ� �^3�3E�3��;������fܤ�.��BQIs��lnO��k�[&|_/�}����
�����W���[�6@`�{�.qJ�k�sf՚��4ZO~�>*]�_�<%��n�+555(����?M���Mҕ+����ݶ;g�Ѻ}�%fŤ's�#�&666h}��"8   ��yyyrl�5�O�t��0�۶k6�I���?g�j�D�#4i�8effv��f�ɺRr���?�J�6m2��� @ ܿ���Ɯ��v�v�.h_^/�T���mo銑�jz���ڢ�ȴu��+X�8�Z��㽶�\��6�& �eT����+��jK�a�W��ZU�U??��zjǻ��P$xW����,(���i��61q�~<����=o�f0�]�T7z�~?�*�c�����4�O��H   @�!�    `Ɣ3R�hv�D���{��z��3�=��ſ�������'>,���r�g9�\�)Z���u\�]:b�Omo\��Z�mXgd���Xݷ���߿�U];�]�}�~��E��U�<���/��>���c{_�ƨ�d�{{�ou��Yz��s��<�u� �S��(�^��s�n)#U����Q�o����?߲1��>��  .4    �1���_�I���Y�V�?LH����B�Jòʍzf���fԷ��}l�MZT�F�N?ˆ�!�bӣ�o�i����?���Ux��j���W�֧������D�R�	����}ck}���U0�01�F_$Ѐ����Rl�L=������ƹR�ؾ	5؛���r*�ڸ�w�\�J�j   �� ��1}G�Z��k�m���_x�9#9%>I[N�Py:g�_�jw�/���Mc��k���� d�_}���r�ң�zlgL�����u�c1~V�%��ڮ�͡��>) }#ݞ���z�*��4WiPT����ۓ��H�����>�>���3L{�#�,�2a�ۼ�P�f���0Ch0����.S�j   ��@��Ŷ���|���2r�!JKKStt����TTT�����ӱ�R����f2??_O=��&M��aÆ)55UN�S���ڱc��������ǈ���ԩS5|�p%&&�n����U���*))���}�M
G���*/st�	�l ������9[6��_"�6��zVj�U����9O�o�~�����^صP���~ٱ�}��>��s�s*j�����jV|D�9��S�$EƩ��B@W�>��s{�bO\Dt�V��a�}j�0C�ݡ�M��5   ��>iܠ􈄠=^�3���sZ�f��t������v���T]�d���kO�g��ɺ�+�m��x��+�W�59BW]u���������:t�fϞ�����p���T0���1}�yC���o*T�N\5�4�N��c;�5B�L�A�~������n0P���6W�m{K ����bE�욕r��Wy�^M��'�_	�1-�e#NQ�=^խ^�a@#԰��P@0�r��C C�f�`�>��R�  �n�@��U�
 �`�I�׼c�����-[����#�8B����ϟ>�� �?x�h�_�÷ҁ���W=�s7�zrJ�L}7�x���I����#�Ї7�|��q:=��$���J�끩��Ή���o�Z���	��k�퀮�[�\W���nm�+?�2e�Q���g�;#DK8�:"�a��   �;� ��.�Sۦj��5ߪ�j1������;O�1h�`匮��.�m�ƪ����̩;�����qu>���Z5���*�J��R��ն6�^�c�<Xk����𐔔����� �GƠ���%@�� YS�]�o{[?{�׶N�N��P���
>���E���7����;>����om������;Î�s��R��<��Y�F��'\��������_�ʿ�>7+��<�5�Zt�Ɨ��jݯ]�=���pj�L���H��C8�:t��j`�c��(��5   �@���%��ZS���V۔�AhH��Ԅ�Xٷ��i3�{hQ��m�S��#�	4�[Vk`����LU��g�w%��Q����\%�U���6��)������;�?kV_���܆Ƥ��I�z=����F�eymW�Z�_�<% �q��?iB�p]2�d��ʇ�_*�v��f٭����y�g)͞���j}w��Vr��n��ڢ��XmrY�:���q�������tۄ�u��3�>��>�<"��ÒF���>k�2��Q���vE�O�E��U���p3t0�~3��c�!�5   t�@��A���r��=��k�s>x�,a��:񉉚r�Dٜ5E:�QΒn����n466�7***�*���1�3�[������F��l�BY]�C7���^:��m�J����t�q	������s�VEK� GM[��^�c��t�yf�aߩa�A��>Տ�<���J�w�֤��S��X��Y;b���ֆB�X�#��9C������_�w�Y-�W9O���$��Ȳ�A�SMY%�ͩ� ���	5�s���  ��h ������3��.//O999}��C�jڴi��mk:�r��v�fΜ�3f�^W__�O?�T��y��uZW�l��{_�X��=�Xy�:�H����{MLL4go��p�1�M��V=;8wϊ���<V���e����r��{�O�+���������E��c{c�N�4��8�9�3�cs��M�]�Ŧ�gܤ�?���gi>6�FEY#����j���� �1�̏V=lVo9q�4�*CBD��嶿.*[�|G��?��&�=H՗B�}xaS����.�Z։��jT\�Y���kFX����z)�}���a����C���  ��h �3$QwA�u_}������8�������W_to��>[�=:����g�aO ˧�3F\��g�y�V�z���r'E���:sqq�6o�`��Y��;��ׯ�Z���w�7��u?޳���i��{?��~�����5���
?��a����װ���St鈹�Ǯ~?ƅ�'�̙^�g��_�8�쁃���V��"NLL����O��F��]�R=��C!p�֧d���f��S��?�:j   �@p��j
�6v�XC\\�RRRTUU�}���<ج�t���   _��E�Ĉ�	4e��o��e�E^��q�z�x��[|޿q��������oiy�&  B3t�*���5   �A�8@ƙ�����`���h�!##C}�b��A��������c  ��<n���Z�
'�l|ќ�|d\f��E%�w�����y�wO�\Cc���+i����  @ ��0C��C��,�6�ЁP  ��4 (2�����2�%����ghz�L�$* �U����+
'�2g��#4$D��w�7�TLW�~��q�5�n�m8�L=��}}Y��k۩ɣu�s|:�����j���  Bפ�w��C� }��_�:��w�Ku�65%j   �� 55�_�ٛ��z%''+}�Ʊ�5�������8����m
�@CbD����81��.Z�w���!G���f���5{�|�=�X-�yƏa�y}�����Ky�  (�0,n�����F���Z  0`h P_����-������о0��/��0���5n�8  id�`���n���`���1��9]�����:^?u����O�m�y�f�M����n�9��G�Kx      ��4 ���$��ܰaCP؍Juuuݧq짟~�����6B�d�9s  ���#��fC�.�������Ɨ���Wzm{�F�g*o���T{�y�/��z���      �`#� �� �Nl[�i�W�[�7����ضE1�<N������k�c/o����d��)h�]Նڨ����W]�c���i�>���5_  4i�D�M�k���:5U*\�q�t�\���c�{��;��j���w����$����(��6�(       �!� ����}Y�\������~Y�\��.��Jˁ�9¥�=vC�������Bqd���2���17�� s����*;;[			���Rss�9��Q���Z���nM�1u���]��]���vG輪�?�q%��uH嬚�7�2�(��ӧ	;���kd�SZ�N���A ��5o������ȩݡpfLq��Ǵ�����b�zz�{��b��uG�M�U�N��~��	5:��      �"�  ���g�N:I�_~y�M?پR�k�
�C';�5�1�Ӻe��f�!�c��R{��@�d� �9cw���hْ�i[���@ ��3���{�K�T�[X�J/���O챝�x|�|�Zx���",6=1c�O!�w������      �w  x�'�`��zlk=�r  t!#*I����vo.V����E�|��"�zl75y�ns����n{�yۛ&W�nZ�� o<�Z[[�v�e�X���!  }!))N�3���f��e		����}56����B       t�!g)�f�?���Ԧ�|�%�U�k�?��i?���7�.��u헗���{7����b=1B�c�ecڱ��s
2 \�5---(���wc ���Z������=$K�M�RzZ�����TΆҐ4L��)��������}5:\Z���@  @ h    ���T�<���{t�[�O����9�kՅ��X}z⃊�yH��P��7�"�����Na�Q���p�U""������GmW�����Z����7��FJ�u��3��P���-����Clj�U��zj0�6��E0   ��FA���`�ꍲ�Ɨr��Gmmmٷ�jUrr�y����RSS�� \dƧi��A�x����v�k��Z  �CӮ�:�¾
�*���ԟ8=.]��->�O�x��%�`�qգjq�=/�/�3���������y��2��ʫ���p0�>԰;��j�,�
�^�v�\�a�|  �߈�Ox�{Β�;w��8�3�Щ�ǣ��
�m�ڪ���}[Y,JOO�5�\�	&�A��s�VVV��ſ�Kn�l���e�7�v��+ @0�0�l}7�x���w�?��@����zf���zԷx_�|�K��;��� �����S�!��j�f   @�h@���	4��3,�222�Q�"5��a�������v�]Æ���8  `�|�Y��_�U�����Q����u��9J�'�z�N�~��/|aT��1�  �ס������Yާ�((*�0C��C�	��0{Daaa  �>D�   ��=��x�a�o���٬�V< ���&F+ZjuK�3zr�Oz��߬^M�|a�)%��v��am  .���r:��t��
�7Ե?�&�-]n�   �w4    H�5B�O�X��/V��3����u������H��S;�Օ#�騴	~o�S�Co}S�?���U__/���HLL�v      ��V}bP|��G�����gW�ͦ��ޗ����*�>C��R����N묎�E6+��VaE��Zj���<1e�%jvE�6�Vqu_�W_W���=g�X]�k�<��+1B��)�`9,i��>�f�J������}���(\����@q��G�b��Y|�5���têG��p��cTb0>ߴ������`Tf�6     @�(�Ď#�j���K���u��ݶ��j���v��RT�[NO�l�_���م���X���.��|%�8�,W\�|�����O���m������vw_N�}9��g0�%fl����?E �����]�.�E�'�]��`��t��Ԏ�4���٦�ܩ��4��1����"G@o1�     ��"�OT$��K_��( ~p{TRR����ė��1dff�Q�w�u 8،��I�����g輡sa�3A��z�C�~q��*Z��蝢e      pph �0jW��Sw��{U
nt4jʬi~Os�hm�Վg4�\�f��gڑ��&�d�i�D�桎���Ά7���@��k&(��������&'j�a��ڏ17�c���{�����Qii�����(,6�M���fYeh ��J���)�3u���:=���lz��jsu�{��.O  �bRM�~�<�ˣ7kWl�пW:L� ��G'����&    �#(���S՟g�Xn�[G|t��PW���ϖvZ7c��>FC��k_U�5�V8���RѮ=g�fdd�б�4k�4��c~'��@r*d�^�F��{�kRR�N>�d���1?r溕R���1�l�����b�?����9 ����x�O�֤đ:2u�f�M�����Rb_W������/��C��0���}--}WѮ/�#y/��X=E���G��@�>E�   =A	4$F�jf�X�<n���R}���:c ��ohP�s��K�V�'��y�<W;���m�+������H�٢���@ard�Ym�cI�'*;6CC��44&]�㳔��@s��z9��s�s�m,��3������p(����S���+F�e���Ay,K�6��3NV��u�    ���    �/1�p��nӳ;?���^%� �!#̐����@�1��        ����z~����H�-�A���f�w�A�	 ���<6��/Sk[�׶�qq���n�U��jn�   �h    �6�SK*7胒�z�p�6��@�IRr}�,�9�)��]]��4X[�fq�䊖������i��|�qG*���G�[�<��ok�[�+��vk�Z,�N��ڗ���. @�f��m�S}]�O�j58s�b�.�##̰~S�j�}��7sP�b���  �/h    ��fW�V�lӊ����|���V]�C �������{�1-i����.�{zЗ�]���m�'(��_���%z>}����j�蔺1]����v�$Ҝ����.��+u��������0���񨤴(,C����--+&�   �G4    a��qigc��5jK}�6��iy�&���iVe    �՛0C��C�Q
�	3t�;�-   PPV�E+�>q��y`�kz9�c}�b���D;v�PJJ�bbb����v+77W�+�8�޾s744���\JO��,mYY�v�ܩ*k�I�B־ϵ��ٜSxϼ��UVVj۶m*��31 ���lV��Ѿ4�Uj�T�\�Җj5U���J��K��L;K.    `�[�ڸ�H��&�l���OyE���)�57;�aK��z��JN�   '��c�Й)���� l������,˶���8�rIHF ���Q
4���E���Ҿ�����G[ZF)�eHH 	Yd:N��{�!K�%ݿ�qd[�<#��Oz+�ޣ+]��q���N�9�'��)�>mII	:;;����#;;���@BB���d'��d����N�Bqq1�f3�3"��r��k��сm۶a߾}HLLĜ9s0c�����h4�6������j��R�ףv����:{[�~��{�����2 3{�ldee!--m`[��"����Vn��h�Z�]� bAD4��ʷ��~�ۋ3����|-{}��-+��G����3k����n5�k��q���0�VY���������"3�~z�)����q�7�{ADDD���
ﭬ�"G���+ADDDD���!'N���y}&MQyATM��F�s�N����6|��r""�qf���Y��KN�����>��yV�� �b��T�i���:��ڝ """""""""""""""��+4���
(I�H3��hG9�������ȿ��z����������)���( $�cpo���J����艐4��PX��D�!.7mĶea�ء;5���(̮��⼮M�Dlf�m���W[�@�[�X(��u�G\VʈmO�5�}]�������;E�N��M��W�

rZ��g�� """""?����ǱC�/�`�j��ڔ�H�G��Ҋ����e�X�3�;soŗn@�.��_Ko'B��nX��W\qnYuˈM�8�;�G4����.yu�ƍ�vյ#6}���k�@�Z����&y}����ت����?'v�}DDDDDD��Z�{�O��Z�
~/;�!��|�Xݰ�������K��5aX��w�ö�C�㩗A�����ş�A;X"��ڍ��[bC�
�q闐�*�/����� ��Vtt����9xzl��
,�u3�������|ς>4�D�ҍ^�S�Б� �54N ��(r{#;�h��
����B�O�c���vu�_2���ܫp[���������R����K�c6�����yQiȈH�3|_?�0���[���v㿏=2A""""""""��8y�M����j�D���N~Ud�P���N�>����B�O;[�!��;��>)<�Ⱦ�ʻ
�bg�-3�{Qkn���a�G�6�~�>�M�~��.|w�����o��f�m���������������F�((�\���P�3\�����5�2XC2�p���4�rBtf_��w���f\�m��2��bWK�؂������c$:QyC��z�O�RgQ���H�ŧ��:���f��\yy9:���DFF�������Ǳ��0�4�u����رc��χ�0�nkkCQQ�[��x������Ø5kְ�M�t;_�D� 5�f�W�AEƱ �^�����L{�aNt�ʽw䬕���ϧ_��=�zK+(x��QmnNᆒ�jhx���4e�Zqq1����(9�Ny��"�U��5�0t]��_$��(;����a�Z����4�VШ�����v�����@oo��W�La�������F�΄�{\V��v��Fl	���?���c�h�I��q�ve��V��:�c������D�<�\d�A�b�P�DDDD�%�����Ykd�aUR�۲��v��r��Ґ�$��`�!���>ē[/z}�ay�3�Lr���n9����9����EW���^c͸�U�w�i,�m܏MDD~.�B��\�(��0�p>4�a>3�ܖ}9�������zK�~<^�/��g�K]*DDDDDDDDDD4Aj��c�\� ��0�g>	4̏��K�~�Y�������U[�j����x����06a���2��7�j�GADDDDDD��b�����9���ީ`H�kiK�����,F�Ǝ���f�~�a� 50�@DDD42��	a�s3��"��]U����f�q�H�v�1�@�e���B�Ղ�����h�"�t����c٧e$U�h��g��V�@�y��Pä�.j`�����ht>�嗨��,c&
�3Q�]�D�g��}Ѻ�I�W��;D��d2���O���t����F��DEFF"##���KA�/&&�g�4"(P���.j`�����hl>	4�6����qY�y0h���{1U���d��x��-uV�B�?+������b36�M�!������KDDDDD�}"�S��lzƧ�T0�P�W�.j`�����h||h(3�c��BfDnϹ��ۀ|cfD$�;so��4��(�V�{�ADDSO�3/X<��;�"e	4ϭ�
�<�ADDDDDD4%�8���0��5h�����2�@DDD4>>r��܌�?�_�x�&/�]�W�3.�g�Ώ��������Z�$�ǂ�ף˿���lk<��m'���T"&��8;���jADDDDDDDAHQp�������?%a?q0�@DDD41>4�8T�4��?�­Y�ᮼ+�2a.�4:\�q�@ۏ�X�S�ux��(Ϧ"���+��{/v6��-���y{�aXp �	�� ��
��!o�R�b'U��j�Pe��Ӯ'A�5j
��QT,U�Ph��|�'NAo����h��%�0TG�	�w�?r���M�W:��H5���פ��S��	�W��窷�No
l�=�W\��k�#7*kS��I趙�����ް�������ADާ8�����*���qI�CKDRf-�k�Ð�?��ލ&]ϸ�e4�Sk�����I���6�����EDDDDS#�X��z?�Z�P�b��v�Z���hWq���M�	���}͹��f{�����ʹ�*��w��?8�wlH[�O�]��+�S����/� ����5�|�5P�z�j���tC.NZ �R?r���/&�d�`WK�j<������bQA�E"� �DD�"����������M�����/�W���ZWtY/�w�0�||�_���C��	�N��a��/��'a��
5�0�Kv��I��%���"""���I�ኔ%xk�/`W����1ۋ��jw�)A-���|��X7S.�І��G��UV���fH�%Id�a�sZ?˭���=�_��7��&��?��l�ߋG��סGDH�T��LHOO?�u��}�uu��?DDDD�_�5����P���\j """����I����~UN$��]�W�a*(x՟p����L;
X
��\h�ZY����{ڞ�F���`�����'|��DDDDDDD��=���P���\j """�����r\N�r"Sqi�b\��k�!/*m`Yiw�s�M�3����@C__ߴ>���:�\0M!����T翉8�Y"����/.++�_��W���!&&F����˱%��1�u��CNN�F#:;;q��)��)�@Dg\�=Y-�(\��Z�L��ኚ`S�^�/�C��p�G�GJR�۲�m��z�3 "��(a�s5J����"""��T���SFD"V%�!%�0�cr��6����7ûM�Q�� "�8E�f����nG}}="�R������DDDA�L��j���ѣr�{��;S�f3<(��z2'�1K���`-���W"'#�m��f�������wS~����H�KF�Y�o�mzADDANt�/~�0a�Ɇ-���P����g�B�ǳ/��i+d����3����Oᡒ籽�0v4Eso��ܙ>�����ϱ$����n�L:�*}��z|���e�bʰ�X%��q�m��e��V<�������X`<Т�ï�v����ad�������Q��<���a�P���}�Oi����:й`a���5���P�g��G��>%��(��ϋ����#x��(:����sDh����[��<5N�>�v{b���tq����0Z���F,3D��/�Y�������4}ˈ���r(0���
���HOO���mmmr�rn���E���'O�����x�l69�ׇ�ǁXy���`0��D�����0��S�=x�޹�2�PC�l/CDDDDðg�����l ����֦C��@D~E�hpe��0�"�lջ """�3�f@ii��.��p82�`��1�f�z{{��K/��W_X��X�\� �"��k�'�U�VP�{�Q��|�O�aC0��}��BA��5��i�At
�7m9��|���ے@�k�ߒ�M\��X^~f�5rc��(ǻM��ۛ����""o(�A\��J�Ύ��M��qg�:dF$�w�/2�@DDDS�8�u�4�;q
D�R�V�Sl��.#��v{j """�
4-N������7�팈D�J,��ԥ�8i�8�:9�ھ�|LI�f�>��������ªU��(+��gZ�L&Y.�]�	|�c�Z�̙3�r�Jdff"22r`]]]]����]w�Q��5d[srrp�Eaƌ�u�O-�|�ĶnE1;'
�;�Q��*7�X�O�]�UI�PΜy�����������_k��١���^�����$�������q��g�Rp�5����r�#S�+8$/�j��9k�$�ɇO��Nr�Taa!���*��.\���t�h�.�~�ڵ�-^�m�5x�����ۺ`��_��c�E��v"
�61��DhA��ʻR�D�Ah�v��7��wp��DDDDDDD�*�;�]\��Si���^�����|hp�*n�� ��R�ӈ'*����C�4e>�}�J[.�Eh�ADt��0b8	d(0f�yf{/^�ݍ�d\���{��C�
>��߈�S�8?g�ȿ�'��ߒ�?������a�?,���q�m���YZ���>h-F�c�wX�	s����?�~[�{l�Q<����k���o�3�L����q�7K�%�M�ǳ/�w�~�b��f��s���#���/ȏ�������w��5���JE�i
����B�� �2�2���7f�-ﶙQgn�d�5:\�v>��Y�2WA���ް��Dvn?Y��Dn��_��u~�lY�cOk1^��@��7D�6��۲k�W"'2u��W�4��G���}ʓ˒ϓC�VG߈����sd���g���\T�:m^�y����>7p;9<�Ͽ$���[�*�=DDDDD`T�����W�8䶚���Hb���UFD"V%bm�R�13?&�m��f���"��rL�}���0������� >>��Ɉ��Bdd$���a�Z����ٌ��n455��4�x�RSSa4��'&��!_/����ڊ�������111��v��#Ե��L&���ɉ�ދ����iS��#�SݵmD�.�x���4Z���"ɹ߈�",!����⸙�V���֧�/C4u��ǫ�W�m�A\t����N�Kn�x޿_�E,�/�U~p�� �����Y�LԘ�q��r�v�$-D�6L~�߷]��@�>ڭ�X�`i���c����{�twݨ�Y�0�aQ����2�.�})+2y�u�D�D�W_�ξQ`b����83���U��P��.��tۚa_�I�T�}x�R^^���Z,Y�DvL�G{{;�W��5�_&��rSQhH�� J����ޗGl{��(��Ξ������T�m�u}�)�J�[u�'ǣ���f�\u�UHJJ�:DH���'Z�@+j1)�(�J��\l��u;����m���_�6�0�x�m����-�vni	hj�J����{?��@��X�k�P�O����~��^9l��f{��cOWm�x��%2 q~���v��Ӗ��փs���\}q�uw�w�\�����юr�Z��Κ_�J?=�,v+�(�ܚu~�����Wq���Fl�̅�G�!�o܍�Ί��?_x�{Roi�K�;��O�J4�|c�M�+�Jy]T��a�<���e�����)���6������
n��EO�G��x�0��yW���JJX����c��������(00�@�⺌�d���ދ����������edd 77w�a!..s��0��颬.9����3��4���zV)<Q�!%%e�aA��c֬YH�ƹ[��Ӡ�jgo��8!��3b[gΜ���D���@C���$�����3-۰e�ჯ��'nLӴ����U����6����|��}X7c����E��^VhC��@4Y�=��a��j �/�/�U��:|��n�4���ٝm�R�:�R�yQi^{~7�X#/Eu���6ā��!�6e)�S�y("
�*��;ytX��'͐�{fn�'s��=?ǿ�����+R�ȡ�<}��(q�@��[�͸����h�e��qCe�OkGZ��+#���>ۧ^�q
V?��JDDDDD�h�i���3B�����
D4�Mg�^c��e}�}�e������P�J�'��gկO[�;r���U����崿�OTl���s!�_8�;\�a9fD$˳�=�W���l\��\��<ԕi�CQ�^������Q�|������o4쓁�K�0�@�>��Wx��݁�b�k�W��n��k�\�}���-�����?�\��m\�?��yKUO�n��9������{D�{1�z�k���cLjd�!$�#|�O����4��z�dic����ϧ_�t�u����r�2��]'�c/�/���L���hY����P���i<����py�yb_��tPv�%�Ǣ��c`������=^4���ˣ�e��dÇZ9�^&/��B�N��ըD�!Q��b�����r���	��UyHTg20��hnnF��b���'���㩗�o��΋�ǟ�}s6������h<җˡn>h-��Bo�š�S|g� ��!�����}�`�RP������>�xa\J"""""�*�ę�7�z DCŅ��;�AL1�x�͌�-����'��DDS��܄�JN"������e���+�����bH��>�
D�%�R��ű�#�����S���yZE#+4�,��ogXϕS�-���R@!���ޖ���/���+�_�����ѿ���{������8e�	
L-�N|⃟�ງ�o�p�w�/�g��o̼D���u��n�D�P�$�b(o�d�91�/(Zv>����0��S�.5 >ވ��@�h�y]�f��Y����ςVw����e����{{������9!Ά�T�U�5�R3e�Qiw����ӯ�L� �	�gw�D�.B��^��׼�}li�""_CNܳ�!|��#�%k�ʻ%⎜�rg~��)C����dx��9u�NtU�ˬȑ�&su�a'\���	s������ހ7�*Bg_��坶��I�X����BQ#�X7θ�c�ATm��ov~���@1��Ui�CA��:ɸ DDD�b�k�bFf44��'=���p����-��q{;�m(>���KDDDH|h�ɂ��2a.��M���_yl�ǫ�����6_��si�bܙ�Wn�.���A�Mt�0�(���c��@[	�c��.u����bᛟ��u�z���4':ϾLIa��A�ET��Ti��_�	�l�2S�>�@�FQ�P�7�N�sqf��3y\�yf��>F�Et.��i5^8�N��b]
�5�����@Ò�Y#�Ah�oC������+��D(�����Y����:%�C����n����hL��5�t�A�NV���a���V9�w����0Ce�l/Q��I�Aؼg�5��@Q�{$�{h��l�eM3#���	s���2�خI_)/o��S������7����ucAl������&Jt4��R�̈L�c��}��_nT�9�����+  :�:��X?{[O��?�y��(�)Lѹ=���8�w	b�
-jj¯�@�j��v�|��2}�s纲��!�um�u2�Y�FSLT���G\�9�z�G:������l��'��4�j|kS��@{Ɉ�߄���K/�7�p�����466�?u?������2�6m��ŋe�H������]� ρ��hT�5��}b|�Ɇ���DDDD��'G���"� h=V���6����37����g��OWm��J���Ċ�`UR�<S���=&����53*m�n�0�`S�x��}h��
4d�p�M+��nljBqE)��'��L��9���}d�5��F����BcG���z�az��M�g._�$}��mq����u��*07Xyp����rS(�<X�4~u�sGN�.�7�tN�C)	]}�Q�m��+�ӯ�T/�/�����l�:��e���q��fa����(��u	�rN�j��b[��Rhz|2w����+��3Ȑ��a�-����T\m.NZ �ֈ �;�g@ll�@�A�j���̄�^q6:���1�����9d�'��IDD�1�P�[�! M4��f """"��I�A��uT����c�Od_10������?*�X&�1_��Qz�c����˱�)p��U�ANO����]A��dv~���3eEݣ�4���y��݉�( ^�_���y��=�J	����Ep��k;9�J5���M����^����}�K�C��2�G4���L�
�˻M�a�Ypu�rT�de����z���*0��R��������h4ݶ��V�.RV��D��}o^V%b[�!�>'l���8"""�b��"g7v�}[�9�;�E����yE{;��-`�����h81Www��ĉ�g_�L&y)�����(�I�!�//u����)K�8s��S�����/Լ�M��G��;�h:ܞsY�Ձa ��η��9�:�Z�Y!�eNt~�䋲ʐz�h"
cr�eIw���D儭Mqu�
t��$���>W�0f�@�+�0R����������q��K~&?�&K���U�œ����{�n�h�+d�aOk1�_��d���45�#;ݖ�u:��s�;k�l��t�[y';�?�N���!M��n���=f;5H���������� ""������Bp�\�+�p����vjUUG<��'�����@CK��3wę����8�l)�LƓ]�`2"A�Ot&.�/6?+2Y^�2fx\^mn昻D4)b(����u9������"Cr�Zt�1(�͑���ߕ�L��oι�����ώ^��+�Η��Oa,�������>u�v�OɐKg�Mq}Ξ-;2E^��px�@��ێ�m%#.�s~ƝW J|V�
3#��r��.\��8�����XA��|3�A�ٚ����~y�Dϗ��#�^����������(pM6���:�}#>	4�1S�8����y�9�6�z|����'A��J�Ot,�[���?t��=��ڡ�����Dݒu�3�p���VV�ɍJ��Eߞ{^�ى���@��MGd�����,����7@4�$-Ģؙ��K�;1q�����a{���E��V���|i\���(��DDBAt��CōVuM�4���Ykpw�9o��㈈������B��n������a����Ob�afT��嗦,���e�@�+��Z����I91�X�DD#�_���x*75ȳE�8�:��/�W��XR�x�����;[�Ɋc)3��G��.OV�5%ϫ�������1�X�����X�U4�&}��.��������r�!]^��+�ߘs��7����������(��b�`�@á�����B3Q�]����K����#����17�ۚm_��eF$���Uf�r��3Y�3��O�yQZV��Ņq]�Ex�p�֡�a��n����(��{�o���w��n���V�s�+�jY��Tw-v6��h$z�7�X#���tx������a�6{[O���DܴZ-"""|�X:ǭaaa>ۧ�?""""���H0A� &q[܏��'��7����f�g�����;�G��S.۔����'�om<(ۍD"��)W��������3D��u����4��k�����{j�}��B�h��C��.���?��p�}쳗}�ӯ�+7by�����G�;�=_�u�\���OM����o͹E��D@�o�پ�҆MG�06o\C�Q���t�����c�:�K����>ۧ4v��#"""�A%%%8r����<� .ϖ����K�"&&F�������4c�9O�7DFF��wtxgd�F#{":;;��*���'��[ܯ���m�+�1Y˗/_�tf����ov{a}h���W'�Ï
�Ě�E����<�/J2���'�=�:r"S�"a��.�DDDD�i^L��y&��׼�=���Z��6k7���s���Ǹ$i��\�^�����<	ׄ��so���ߕ��:K����lD��Bm�s��>y�z����5x�G��E��E�����������p���q�g�������2f["����7���&L��`�A��X,�Z�𦖖�g�v�x.�W^y�y��ܷq��
��'�������\�4c5"��㮺<T�<�l����3������w��dh����ˊ���Q���>�D�����vaO�Q�OXVܳ�!y����yTV�rZz;Qki���9��h~q��U$�;��@�?���F���m��J^5;��R���{-��9�[p�<c���ܟ�~OWncu"��˸yQi�ri�1�R�!%<N�{��~p���'����Y��N���_�u-n4_,��n=�|�|D4��т��= ��j���)�����B^ee%����M�r������o~SVI�s�(���6UU�|�嗯���k��,� �߲�'x!�Rܙ��1�ջ�:+�ײ��lջ#�W �I_�Ӧ:9޳(oJDD4b��}k��qٟ�~�Ę�c��.����<y��sz��kwM�����{��z���wU�~""On˾���a�{}x����#�C���4C�� q6���叧^f���������Fd�����N(̐������3x_�sz�^��@� ���g�V9M�8X�t��@DDt.�̭27�|"""Voi��b*{Gmw��4j�[��J�k�,M(�]-�N4��˪"HUknq����������ɢ}��}|EQ�F������q��T�4����&��Т�D鰱�=1㑔`�&�+������k{��b����KDDD��mۆ���	����t:�v��EQҝ��W��Qȸcσ ""
V/SNc�j�w=����ߞ���_���ۇ��q��N<'��8�Y����<�����D��p��qu���m���P�3����Lr�꤄0�@DD�v�Xu]a��������4�03����D�.����?�@DDD����v��	MEQf1�@DDDDDDDDDDn�3��BɉQ�3��BɉFQ`����Di�ZД�`������������tu[p��	��~���T�����u�z���@s�DDDD�=4�W$�F`Es�O�x\�tVPp���}�@bl�46w�)T45�ˉ�����DDDDDDDD�i�H�����c5E�0��;b}�O�o�M�@�?a�����������B��#..�7�Ӏ���`��>��������DDDDDDDD�"���R�4�h��>��"""""�@4m/n鿮j �~�NIU��Oǲ�DDDDDDD���"""""""
h��JF���$lڴi��Vᦖ߂��������DDDDDDD4e.NZ���V�06F]��>T��n�a�P�z���ձꓨ��~�W��,+ODDDDDDh """""""�ˋJ��+�-�|6#�,������r�.���j�Xn�ֆ�gJTP�T�yo���&(h�b����BDDDDDDD�U����CH5��dW5��چ��貙��0;:פ���ԥxq��ش�x�b��hr�3ިŢW�О{������G��F������{�} """?��7�/#���^}��@��O��fB�V�ן���#.c�������������C~x�1���`Wn�_�~S�.K9�����Ӳ/�ƃ�67���&�#C��k�7� :�^�f:�τ8��KDDD����}��xOD{q?o���>��Z,�	�!D{j�&��G�@M��C���_5p{��Q�����	�x�:3�5&""��Ǔa���k����٭nm.>��K���(+v�nqk��8	���6}xn�[��N&!�4ئ��潳ڬ,I@bw���n���vb����h��}JһP��=p[ߧ�ڣ�nmJ��O:۹��5Xwؽ��T�3:n��
�NskS�b���N�y>Lw�]�d±,�64hY|V'/�O�������ƃ�u�O����d b2�����}�ԩSؾ};�̙����鶴��8v�vv2@Dt�5�0R�~��f """�@MZZg8lM�K��$�=P�h ""�v�[� ̮xl�`L��m�K�v�#�k0�`��&�]��N����h��6���m�m:"�{���7�Ž�rC�Ž�:�MS�{�C��ڴ�j���a7���t���d
�I^,/E���Ұ�;+qi��~�&���`����/����:�			2����6pI�D��-�0V�~��f """r�@MZBv�=�
y]����Nj=.ĢE��u�͆+ρ����S�!N1Q�]3���Ă�\�?�ݲ��DD�&XB����P�DDDD�1�@DD�����5���c�tvN���U��t�Ry]���"����U��ZE�H��6���{/(�i4�����~F�O���l�R��R`��&ڹ������<c�����&..nR����TѠE}�Xd��/:X�3��'jfZ�}��~��vD�����9ۄi��w�hJsk��C�{�ȳۤD�78�D����&����HD�ªmRn��dgG��'22�L���:��lctk��9C�h=�1�P0��F�&�hE�ɽc=;;��vLTrM9��a�ث�B�*꬐��W�٪w�l�7����x��}P�ϱ��>y�pG&��H�`0�l��؃+� j�a����j`�����hd4ѴgqѠ{.��D^^V�^-?+w�څ��≯,n��l��m��n;�63�n3�M��m�=�G���h3gmf��M��m&���Ahx�a?:�L�ŢO���c�17��V�a��ү R�窷�_��W-��c��� B��Zm��>�;�Q��εs?�B3���""����Iݯ��	��� 򵌶d�D��;��K���̴6rZ"Gm��n@n�{�#ٝ���n�t�#�����#Y�	\OR����g
�щn��z��D#�<Xr�7́�9�n��S����6���s��̮�F�i�M�VŁ�6�6uF$���m�g���������؛�
":w�l�+��b �'������?a�{�9��ػ���ѿ��ʭnCJh'-��wau�B��x/����j-t�"oٮ��>��j�V�~��f """DD4iv��^k��ik_��:�����R̙;��z�PE����I~H�����|<��!C��tos"��-� :��nS�ڍ��, �<��T�hH�ަ<��-А�`Df�`�;�6,� BYCB�1�4�l�Bv�`��>,А�dDn�`�^�cX�!�9R�#\��D�1o޼aU��ϟ�@C�Z�`V�\�;v`[�)�ߖ��4C<�3�V������_���j�Y�e5�Y�LĄ���j)�M�~<�aU��h|�=����}j��%"""
V4Ѥ=�{}gp���[�kx�}sp�DDD��>D||<(0-Z�Z�.*B�L���<�7����so��)KP���hG9�t�<r�U���,�ND�oD���F�瑟U.���}q0�@DDD4~4�����qͣ�����.CŻM��d��1˘�}4�mT��b��^{����s��B3MDDDPj.��xe]3�#���6o�=����D3���\d���;8Dz��6�z�i�fp�1kc�&E7��J5]��G��bb��Ќ��^�α�11��γ��6���6�`�>��6�$b��M�:۸},�2:��a�Cm&>���c���ADD��b�ʊDD�D�a�&����S��`J�PC(m/M��hDss���p8�(,;=UTUme������Q��֞%�l�E]���T�>}���D?|���,[��U�X�pm��=l桍zV��3��zr�g$�����9+fb�8���d�ψ=3�sv�	�Ul4��]�C��{�m/MܬY�P^^>���L&��)s��"""
Hk֬�_0������I����ȫ.J,���wN�~�����;�/M�+��o��ք�}�vlذ45E�;�Ȩ���ݪDDD4~������w��h�"<xP����b0䏅�����{ "���b���ԥ�_yO(�ma�3��j#�ѫ���[���}�"�S�F�'Zh�!��#"""����B\z�ضm۸���Ob��լ�0TUݺ��'h�"-d*�pN�0 M1 E	G,�㜢�C��s���A�lPх>t�b���y�Q����Ɍj��Z���J�VDD���K������vP`�3g233�t����(�mi؏��&^����
|��1�x��<�?g�@Yd(�-jI��>�������#��pd+�HU����E/���(:D;/�G8�*t��N��Kku^oR�1VT�S%z`Q�""""w_����Յ�����>���7�_�B��G^�^������w0�0I�%G�B����)�y]|�֏�%z,:�Z�k�w~1i87+�P�8�v�څcj'*U#DDR���O�-**j�z�0�����f�i[(4�t:DFF���4
(�����n��.5m�py�u�s��(����a�B�\&֡D��8��+���:|�vt�T��YO:/��W"""
]�����~�͛7��_D}}�������=�܃�o��V�����O�JUUh4YmX\���V/v=ǉ>����bv��G9��w9�O���q��7n|�y)���	�P8_I�2M<(�ί־��Т@1��J��ybȊ�j��mΩ��DDDDDD�X,455���ͫ?���tDՕ�~�{�؆��Z477O������8���ȃ4�UI��<e	�^��z�@�EL���}�XJ��D��W�&|EŻT���Z���"����v&"����%���Dݓj'����h�V�%""
=�X������(���n9��&�	����]˞�y9M���+���=-c�a�#V+�X�M�_p���p����(oW�=x_m�vGN�&Ph�B�
Դ��b��ئ-ʊf�������5��֒Q�،NT%�\���<�Q3���w�7�6rZ��u�Q��0�6�FZ��`�m����ks��t��R�ى�$��%""��%:�����g����M�����bݺuSj���[o���SM�!|�`�ܹ>	j���8������;�N�x��-<W�f{/��(t%*z\�$�M�+1��aIQAw�+��59rȊ=�Vy����&DDDZ�	b�q�eh��xSkk��Ξ/6�?�R�p�פ�r%UVe43�Hܢd�M�7lu4b�ڀ���Y�M[z{G��Zo}H�� Y�Fv�����O�D��m���x�ISc�m�}��Fߦ0����1��*�a"""
nG���ݻ}�x���8}�4����1N�:�0� F�رC\X�p!hd;�����æ��X��TN���<Y�6-ی#�����3(Z�V��NI�M,-�0�դ�IT�}Om�fG=��N�D�/��-!&1�Ӳ����h8C|�^�I�5J�RB��8�F�������G^s�b���,1Q?v������%�2���� _��̙3e	t��ډ���Ӳ�|f�5�-�r|��F9�o+�[�d�۲-�\%
5�L�2-��NQ%�*%Wi�P���o:`Ϥ$"""��F���k�С2�#�]p|�<a�`�&7k���D"X����9թf��u~�C/�'%""""�sS__�����5��~OD����Z��&����<���X�;r���%2���»�J�n<r�U���!TF^����3�BI����I6>���&m�5��Q�FV�%""�i2� �0٪b�_	�@�(wv�&Sf F	C(IW"�Y��[�����
��kl """"
b���>���h̞={Jc�ܹ8z���Q�K���,:�z�x�9͋��]�W�p�M3V˩���;�(��zDDXDp�%AV����V��p�&�h��O9*��`�s	C��	BtttL����4���fȊq� ����߭���jf�i{^u���3b��(ĉD��K��)�"�&NJJ��}A|9ljj��3�###��!���|`DD��xb��w���1������z<xP�6�]&Q�a���)!�4���ķ��y7g���ދY��K]�@Q�C�~R���J4B�\�I��Tlv�៎J��V3q�{2�3������	O>����!h�-ܣɗ
hP<��D�H��~;Tߟ�EDD4�D��{ｇӧOCU�6��������ˎĩ$Ʈ߲e˔��,R�K�,��ŋl 
0���X�v-YTTV�Z5%��eee �g�^�� �ʽ
��Q:��_gn�������3LD�N|������,&Q��T"��L�TA�t�ϸ���Ӥ�9G��W�
��EDDD��<!*++GLF�D�![��4��XY�b��t�q@m�쥨Q� ""
"������T�/444`��ݸ�˦�1D���o��2좪Ş={d%�u�ց��ȓ��D9���ydE��Ҋ�����8�#�����0�e˰i�&YA��łwK�ag��3?��hdb��M�9Ă�J@��;_��59X��������nh����(�u�A|��Q��;�_��{ܖ*���n�uT�i{%�� "��'��
3�TVVN���٧��&q�S����"""!\��i�pG�:ܐ�
:E��⭆x���x�v'�^�cHu�������`@JL"��%"�	Y�I����(S;�T0Iu�V?��M~g+E3zADDDD���|ňoj�"W�M��L��"%	���:�gw�ڃ���S4X�X^N�z��ű3������ U��d��jFM{��׹��'0���y�Y
j#�o߾���On�q�(~R=9f��N$`�����U3�1�s��3F��Ԩ��L��֓�>�6)8���,I�����t��k�ʦ���Pb�����dD�������Z�皧,�,�Æ7{{\Vl�ƣu[@D����f����ɿ����GRZZ�@�0&WVc�����+���?���Ѳͨ�i/_Aun��(P����lZ��~{�&49bh�°X����8&w<����(T]�A���N�����*��T��[�<��?�AU�ᶴ5���"�oU:�&u_�͆*�]W,=�m��ǌ����|��nL:�ƈ�J�J6�T�=�s	�w�1�@�Agg�2��,X0��g�fee���
����""
m�/�+? ��l<V�&�Z��5�oPpGbb�O+¡w���}Jk�ĳ�Sb�-�\�� :7F��u�\�I�ol%p��-������/��)q �ѝ�� ~���V�~��
Jhoo��}�v;ȷ���%$$$���^�!ѨQ�@��j���L��6Q�z���Sh֮]+�Ө����g������$"�Р�h���OTlqNo����!�hz���j}76�<>
:T���)�Ewjrq�6��P�l���ٺh<h/�1�DDDD4��	4�V��}�|��6��)���n)�G��	"�����~�iS��ӧ�KQ�"L��&�O�6�͎�o���f���0$%'M�ci�/�N;�Ƕ�aGήO����nC�����s��K��m"$��o����l���5���1g�CNn����׃w���i���*{�r|��4���U�0~�}ʧb����b���J8~�[���x��۪zDDDD�&(5��6߹1�O�D��_:�l��^�͎z2��)3?&Ze�R�a���$�u���q�a,�'	�c���!������]��9ί/�O��F�M�,ň��#�CLL9-|J��\%
�N��!DDDDt�Aq���6[�@�����<���r��0�E#;!'CU�s�#""���
N�j ��jeY{"""""""��X����4�	��}�r%���v�ꗈ��h��4�C�ok��"M"hz\��D<����D�%��������	|ս/���h�ly���Ȟ �@�%��@Ji�\(m�B](-em��q������B���R��,J	KX�	��8���63OG��K�d�tF�}�;�4#Y���9��?^�7�ۊ��� dt�'����=(;�@ó�>;�떖���N���a۷S"""""""|L��W�I�h�!ӔB��1w�ob�9��,DDDD�#0h��1�+%��:]����46��ԑd��@�O������5;QUDDDDDDDvԨ��.}@�U����|/��= """��lh�F��9fa�R��l�?P��6�{r�,�In���� """""""����	�L�ɡ|�1�~o�� """"�D��0Q) �e�R����V���0�����"""""""�봉�%eI.�wCw�7b#CDDDD�	4�+���f�Ab�"����Y�-��@��X��2)//DDDDDD��Ly���}U������a�i;��Z�,��ym�K.���g�7`��"""�\f�@C����Fp�
 �m�R��t��w�Dv~d��2��"""""����2���i�׃S���|�^�v9T��c��kѯe�$�A�����X���?���-��e�����(WIhP��Vmf*� {�y��똆��o� ��R)�mmmp:��l;??�(
����H�(**�{]�� �������]�\eF��ϫ@�SUղv��P��4-��T�[����8�=��Z�-}Z� ����r��k��8U)�ˇ"��5���؁l�
�I�h𥥥�������4Q�x�ͯQ�D����.-�RܛAٯ��0m���ɜ����d���+�h��o�߀�_A����胤4\��s-7�_3�x�8�lb�2%/˖�������d�!f��7""""""�d�W
�=m:4V6��q������w���q���(�Hh8N-��	 {�V���f�4�cMKVg�L˶@��PCl�a""""""�dy��f����0D��ϙ���N�)[����ab8+��P<�_�ס��A�L<��㓾�hnK���[,�
�hj8�DDDDDD4Z�w�mj��.�����*�DDDD�B�@�*���@1���P�������l_-�E��iI�~4��������˅`0�l#B������E�A������\�6�d����7:�`{؇�DDDD�@�@�UZ�)���2S)����}7�KN�D��l4>�n�;z�e{����޷7�q/����DD�h�R�k��"��]��o��#DDDD�N�@�L��Tǂ��Uj���d���h �@CO�}_GDDD$QiӦM)ݦ�DVYY���r�K[[[�������Б��~��oA�PX⊈�T���VmZ�.e�Ɋ7V�O�"""�l'M�A4�o�4�Uv&d--���䘊���"D�h """J������
ӧOǼy�`%`X�r%�y���m�����Q<��%&�bt`��I/DDD�ݤ	4\��G��A�l7�hz�O�N�+4�h ""�D�}���CCCƍg�>v�ڕ�0����'�H�V�q�Z�nbb�7�)�zx�`�%e/)S�"|\����z�2Z����nh 0�@DDD������~8`i�����Ȅ��j��	�k���N���Qk��ne��D��H#�KM������1�fx���4�h ""�D�x,ؽ;�������n��I)�	&���DDD2�R����_��x�W-8h����(e<�p�Z��J(�����j<m��0�@2`������q���駟FsssZ�'�S�L�tӦM�ƍ10�����̛7D���BYYYZ��1ݠ�'�q�:�4S��U*n\���Q��K����6�����QF����h���HC�E����`��d�@Q����CӴ�nS���.⽫���p8����遝U��p�7�@k����P�?,�k��ƔN%�b[�7JХ���_���YyNb�Ɵ�Y���������}�cزe���=ǥ�� fΝ;��

b�]t֮]������}8TTT���.�PV$�G�FT5M��:?���S�>�_�N��ePr>�V�D�k�Ne����^�4�.Pn*U\�T���`4�� �����Hd�G}Ԓ튲�g�}6�N'���ى��z
��ݠ#�S�E�U;'�ۈ�Ң��Q��,r�Pb��<]33���=p�?!��6�ԩS��lQ\\���:d_NS�D���ֽ�2��N����#�>%�C��l�Z���������W�M˾L9�A�U|_ -���15M)��j(w}Q����5�������M��p�cZ(�]�����~t#"1!v�UZ9���B����݇"ְ�Wp�i�Y�z�D������	�\�B8p� JKKA9��A"�8Lǆ�pjpf�k����p�{��)A�w����]��h����R�|�?�����*�Qn�:�S+��hQ6�X��
�����t �3?t��˻��7�"�Bŉ��X!��K�z���v��$�DvRPP5���#�v��ii�AT�DeQ��|K?t�P�X���M��'���68#8	��SPl$_��t�#�	��>�O位��}�$��4K)�	J�o�2���:���۹��~V��|�[!�O�������DDD�E2�3(����Z�lw��[f�o�ٷ����d��n�=�P'��>\��������R��
�kec��㦘E�T)�9�?v�V\P��;y��"�����c�_�����hʝ�ю;�8����iݧ������X���c��-(�ul�������i[7��,ul�W���2#�Ց��b|��T��w������ Q.��6��g����
�4��i6o�6�^�l����B��_�׮	��/�ZA��_\h�'Osy?<y'�!��[=Y-��C���3�J�0Z@DDD�-2h�H����)���ë�������z{�\�}�6�˾���������c�W
��'k�E�4��)>���o����r�A*꺞�m��,7��ۋp8��}�\��,o�ˬY�������.ӦM�t�bM���Z<x� ��9��SQ^^[H0�(���DD��|Ӊ��N��1��A/�-�g㉼M���m�N%��0Y��x�٨!�6ں����
��)\xg=��y������P/��5�����鼲z=�+e����z�Z��Yn�L�g������J�n�YW�At��d��Wmz�l���nd��m���?4�o8S���t��s�*�y�����6�Dj)���$�\4��~��lK�Gh��H�#��=�\lٲ�����
YS9��vG�<�&�/��ݻw�,�A�5TUU�rQ]]�H�UTT""J\�^���>�r#=�|10u��	W�^�K�W�HD4����6����ly~�����=��7>ձ�[��4�ᝅ�/�3�n��U� {�8��n�e��"""�l���ڹj��k���^0����[�j������[����{���\�)7�����9JͷN�*�,H�D��s�J��h��� �,���%�L��dq��?>���2ar�_�}��+�����M�g��U�R@D��*��<��b��3���l�������\��m~!.O>��K�qV�t�V3ޓ%��K�z�3�@DDD�!�-���:�>��l2�-}���g�٧�Һ������{��N��L���J��ƫ�O5|L#u��H&4�N؈_�B����_T����P��\z�J��fE�t��Ug��(i��e��w�f������v��q�
�(��? "ʄ�8�`Y�>��~��F�'zۖ���r����ך?�P����Z���*�UJQ�xp�d������/�=Ӕ"LR��kp>j���s���=�9�w�q���X��7�.��'P��"�n���}�96ĺ[M�(>��%���#;o���`�E׍z�K�)��{Ftݚ�r\x�7@Dr��?D)��iii�ә��쮻�;zI���~�3�'�u:�#;�ё�t/��7/�a������|�O��!�Ȼ�a6��]�ޞ��}-��
zA��Ԗ��S�N� �f�s��\����֛����w_�f��?g��46�e}��7`�����}���U�EE���jܧ��ݥ�wa�ͫ3t!���w-}���F\�F��8�}��+Θ�����V�_]����g��9F��[!#Vh �0��oU�y�����=�@WuE	�����RWU�P0��-q��0��E|��d���m���eee5d!f	h ��r�*��*
y>��j�8��Yϡ+(��ө�f:ϥ�i;��4Q�$���vux�������9m�3��A���>�k��W}�t�Zb��ܯ��i���-����yj9�j��3����̚Ƈ���z>�/�s�_��u�}��[~�?C��o�a	�4�LGt�-�&[�A
�L��~+� ��'��H��K&���~+� �c*0���d4|g�X‡��3f "k\:p,ƆK �y��x�yk��e���444�e_�{;(�����혂�vq�Z���?�;~���Y&eI���.���M{�Z�{�l�ʖ��ep�x�k�N�Y�'��� ��&����Ch���X��{���=r������ۮ�ݫ8p�R�W�Q|n����p�������(/�y��Ң�W�+535�𼝉�PQQ8�u���ѯyy��1C��F:������0����83pduE��]��YG�4�Ņ(�xL�'+e��^�E��W�.���!����v�������2�^�7�8NW+�Fg������-m	�yJ%��M�;�Ў�;�X�6��e�W������U���f�E�I�Wu���@��N�|>�:�}߹\����cM;ވd��kS�:;;1~��h���I<���zL?�h�>�?gT��E�t	���Cii�{aԁ����c�޽ы8/'�������X�yDDv�!�y���A�ҷ~����v�����l��\�6v*l��j~��j�ɽw� -�T|Ȇ��m�O�Cp��;��O�aЎO������̯�&�0Q���Ω�e]����@�F��(9��t]��<Ȟ����M�`%$����¤pr�Ep�N��3�K�}PQQ��������úu�iӦ�>��8O�mF���7��iJ��o�����[�}�y��s��s�yj��H!8N-��U���Ⱦ�h���.5|�����?�Ε�^�M�yŒ��-�⒯a��*%�6S�"��t�o�r�f��d�@�(��i��y�)Iݮ��
��χ���H��NäI���3�D��ID����c�M "�#
NPKa'�G�>c׃O^v��`W��~���"ݹ���6r�R�5`������+-������3�� ���~���6�ʥ=Z��g~�u�1�8lT�\3o�4��@�(اYDD$�Ã���o7f�,X�`Ȫé����?�q<��c	/�vjpDd[Ӕ"xӷ�pJ��8�mɥ�]��di��E��כ���J�
����+ CDDD�A4�Ɓ��]��ۑ%�]��[�=r����1'�&Dr�O�	�0�@�a���(y
DD)sRp,�ϫ%%%8��
3*,,��矏�K�"��v�z!��حq�*��\�Ugx��4��y�Ȋ����6����ӷ�y��2�vP��F�C���Yh(U\��5���	,��9Y���8{�Rxh�Z�L�4���D�Yה�����
�4��w���d��tw�!��HMg�&�i�(..@}}�������'M�d��m��(e������(8묳�t:G�ﲲ2�t�Ix�����(�@��qJ1�" ��~��S�B�W��?���u��H�;6q�R�f�DDDDvdy�a�b�%�t�Xn�N��e=�2��w?��Uߙ�O6H�Y��#��+f;�hh4�(b-�<���~�ɫv������g�G��%�����}S��AD��iDD4z����pEB�9�cPYY�T�9s&6n܈����fJ���� "{qB�1J!��)���<�,��r��9(�5�l`�R�'�@ٓ偆6
4<g��|����Y������c}��sԚ�����rX��d�v��r�~|z
�PV��Z
**
��՗�}z�����nĽ^q�'ZA��$d򽝈(�/�fb]"��J��%��z���f�^""����.��7��'������]�d߲���͗���ӤC"""��<�0�&�aQm���9d����ϟ�V=�����0&=HB��V����^q��O��5ZV��s�1�/�u+�LD��
DD�Q�'��������*��c���	
7
L�y�9$"�t�>�^4Zo�|�>d�Ef�7�=_��I���ŃB8Ћ�U�$"""JK��x�����m_u�+��V4���]��L�r$7A)�.=a�a�Xh 4�""""ʌ23?��[f�����x0000�۔��׺A��t:Q\\��}�U'(����uL���^'ڤ����+͞�"�5>��~���(��}���~��""""��4�P�x���ˈ�0�ڿ���v�<T<�A�i���Y���j2}WX���%:v���	KD�0���D��MZ7�X�	4�M��+�HT���t����9@Ӵ�S�.w_���c�����nEx����*�:I�J���DDDdG�&��췌�g/{�1��X/Xtc�l�D�:u�#m�b��r�� Z�0�����|�'"�f߅����r���{b1}}}�ڇ8�o�}�}��(I�eA����`(��A�D��2�.��s7n�N˾��s�`���җ�e_>d�*T4(�U�Ʉ lR;nE�X�,���㞝�z@rv	�}�����m���1{�"�lQ|��F�U����1�:2}7h i���V���i�g�ʛQI�����;�m�@��ў�>�`�H"�1���)���B����C!X%�m'z�idĀ���(U:��c*�Zq����ͮ��/yx=r�[���B�-����WroReKՊ��@�Z� Ǭ3|�q�f\�
�UC��ZHVb�	""""�L	(��F�J�����WDD�T{|��i��������pэ]ǩ%%�X�b�ch44C���ADDD��t:c6V,4ȟ��f���}����1�_�������3K-.�Ī!�1�@Ɋ�"��(Ϟ2M��u+�� N[?�������^�����U���mGo������y(�JQ%���?���v1\U�T�殮�h��DIQQ��K躎����W�����$��.�@ :�.���"o��P��~KK�%������~�:��-�CD�N�6��ab���+��F���Ԓ�!�r�ᄊF�<��%�.$"""�	�B1;l�4@�R��1�9� ��f��HL��0$+���#o�A4�x��ǰuG��Ecj�0��y�2��I����K�}��±;�����4i"�������Ǳ}�N��ļ�ө��u8�¯�FoժUشi�?�4i�:�,��;;;�lٲ#fɋ0�y睇1cRXioo�O<���_�g�}�%���W^y6l8�BCC,X E��,�Z��Ī"�|�h����*��c׮]	]�W�_	Ip#"z�*Th�i�<ك�����P�ԁ�W��p�>�LDDD$K%�ɉV� G2�c�:�P�X7�+4��h "J�샍�����
5�0Ä���wɷQ<y.̚ր���j(�z0s�X���CQ�YS#�xgϐ�f�=u��J1C��aa�����̙3-��ʕ+�*�
����[0X�~�aA���g��UW]ei�c���x�7����={p����*dѢ���N�͑w/lܸ1<I�0��[o%t�����c��d"KY<�П�aa]A�C�������4J���@DDDd'�4((P4�̌��9��(r�>M�G�op��3R
#���&�����r��i��%J⦅�nC�P��逯?p���.�ʋ��$_�>�톦��=}<ڻ��y�1�e��G��8�}za�z"����:��}Eia4X�gq��t����VD 8�Rb�	+�A졈P��Q^^���g,�`��PLl��03\3�ۈ���ٳQYY��� ��g��DDvRl�@C�Z��m�/͋n�+�BH�PG""""�e����h����O?�9�����u���e�;}��&(����k:AG�Hf�J�X+���!o;���#���9�	;����L�"���G�E�1�˝�2rnwB=PUe�}�����,-�3���c���v&��~�6s��5����oi�!�����"�lrJ(� ��+V��/�.K2x������f�I�o/�����a��7�v8�����>ȲL�"��$6�#2�2ŝ�Ծ4��bs���($"x��l$�bpX,��Ab��J\������d�#��Ӫ ��^s��%�BM����Յ��z
,�Ñ\��Xfeٲe	Wi�z�[�Yc����a�7����DK���7ʼ9Ui;��>~3�� ��}���a=зE�L�ļ68�����>Ȳԁ�N�� �n� �p�ԁ�X|�y��ܣ�9KD��h�l%ӻ����c� �@�U����O*��{��&�h�RWi��J���~<���?~�����g�I*��ڕ���"?�@}OAZ�UPÁ�\Pp���Ly[�����cŕَ�Ð�ƥ�{��bY��	�a9�����/�9�B�,�mD�F�����FKS��(�___��O?�����[�o���{�`"�4w�\�ִ�W�iӦ��rE'�x"�N�
���ԕ+W�СC�5�� _MM�>�l��3z8�ǣl+�����F,��@C��Zh��}�~���	橼w4---x�G0gΜ�{�pm[Q�l�ڵؼysR���Jϻ���#^����iٗ��s�
�vL��Ht@��&@7��B0�/��A�=�Yh���-�LS��i���ArX��:Rb �Hf4���ի����޿����ݻ��s��.�t�;w�<j}o1���K/a���)�onn�o�q��|>_4dPRR���jXi���G��ŀ��I+��͛)�$����BA���x��S�~�|IdM�����SCY��3����3)H~���m#�J�؇n�4L��WM�x���*T�kKN�z����2a����.O��"|'�x"�'�ǌ���R���E?���w[[��݋}����3ڳ��WB 먑����J�����h�D/}����x�4�M�CrN���Ȇ,��������0DE8�e����$�l4��_wd�X%��������1q������Xmb�v�4� fξ?��~ɔ��"s[�<�\X���ҡ��|~�w�D��|SNӔ�{���%Pգ��P--]P���b`���N���WF䱶�t���ԉw>����2�䄕��
�Q2��x�������s"��;Ǌ`Ö-[�+t�~<��DDv�H��j*��@�fB��s��6FDDD��F�t�a]�b}}iɹE�)D!���!���)� J���P%�gZ��Gb�>��dj�]�A>�f�֬���M�C"��T}��g��o^��h:�N�"�*� �"���*��?�x��j1���+**����)}߯mdj�x��BN�3z*\`e��x����;أub�{�	L��D�B,9ADdGa���\�r~�ܩ�e�\L��X6
f�Ah�D���4�٣��6�8��;����oϪ��ٮ²�i��s���g��������c�?OGP��|-J
���tx0DG===��n�r&�y�b����V�7`*S�A��Os�1v�y�^�[!�`����/�n_}��t#Y��G(<|@��&{�y��\fe�!ֹET��E���Jww�Q?�2���jv�س��h��j׭to�Z�>ٕ��y\D*4�AS�> """�DXh���-�J�.p�.�B�ڧn)��C�ZG��pd۳"�0��x�ZZZ�u�V\~�� ktuu%�.���A��'�*#4�t���G����-�V�C������"п�iq������p�+��Ǿ!����fu��x}2�-/w8PA����8݅y�39���P�d�BC�m[u�$C2U�A��\�����ƭ=g�kZfI�NG�<o����B�L�&�Gq(���e�s��K�:M���Bِe��~3��vӥDq�5e$JU���>d_IPѩ+:;��ٓ��c��K�#:�=��0b@p��Ř={��nk�M��}�	�Z`�ah�ԐZ�䋷}�f��z2�~���`��>�*0eZ�󊕯�t��۾����e�R�.��LjQ}�e������̶U�}�U�)��Q����c"k�u���ȗ��
U�HN�㈈��h(��,�@��*%���Ԥ566�dKN<v�΃����4X5�!�E'k28c=��D@���5���j2F:i�a�ቿ��efR"S�0�Z8<�{��_b�C0���x�긲K)vU�וt-..�6����D�e��PGPIX��F�VQY�8i�����o�r>�p�w�4�ei�Lۥu����U߇�o��y�Z~�]�^u��o��d�k���� �qr9�`:����@ξ-"""�x,�ԑ�h��#��|ձ\$�_Fzݹ�Cg�2��/�����6��PWW��i�CS�}ϕA�A/+��|Yhhkk;���}M��Z��63�%{{��*�������D�܊UA���a���hC<C��yݎ�:Z����5�i(7�{n��l��/�_���H�ؠ��G��"��)�rH��W	���������=Jy�{p�����@��㓒?=�13��f��dg�@+3���I~R�0�ʰV��ĆU��X�q|Z��d(`��^���B�2d�w�K��UR��aw��n�W�S�l�I�c���x³	��{;�=Q��6�Y_��O@����[꫔<�+�
�&�~DDDd?�������dVb:�C�*U\�?�X���H0�@��k��(�Če1�.�U��x��ъ�m+K�W����Ē�����2-��0�@YL�[��ۏ��U�x���XN(�y��IbU~�}	ǆjqe�	(��Z�n���NG���M�"���csuy�n�_��ڥ�RA��ٍ��`�"���w�Q<���L�T���I��!����0�@42b0]6�����L��.�`�X���a��;e�X���m�T���2��Ub�C��İ68��'q�"�LE���	{��hU�u�}�� ��$]����B�@T�I�1�J�zm���l8�C]��Z��1�b8Br>3�>.9ADDD6dm��7�����E7\tץ?9��<�͋Ou�;!�f��%f���	�D��D�!S}�-9aq��xe蓷��h�b���@0L��/���0X�e�v�U�r��U a<��+��pl���aF���C�S�X�܏ծ���h��(�4���Ǔ�}9��qç>�%}�uL)����C64��v=r,аbŝ��N}6$�{CDDDDdi��i��@*���/9h�W�[aa�c�(�D'��4���'�(�~�С�~nլe!�@��KN�۶U�|�@ f�J�R��vU��p�0�:��b� �8o�A��εV���9�KN�FX1�ֵ/za�	�2L�+P�{Qex�o��60~�ѧpH���0�stq[R�����"-��kv�M=�6v�oi:�$��.��DxK������3��N����2�#Vtt\�a�R��1h """�J������`��;�����t����.��K�'����?�v"l@�c����h �X�M�\oŬe!ր��i&.V�D��x�-��B���D���/����S��X�9qNm����P�+�����E��A�	A�gk�B�׌<������s���X�����ZI�g�T*S�.�ض�#��	9���v���'"""��$�����>5�2��Ä&�'L���^u�?����k���Z߳8J!ؗ�rz3�]�AQ13���n�ϊ@C�f�$�>��4Z���MD�6\��T�H��>��Ԋ�j��e���O�@�P���9h�a��S���`;�����(�RX#�d ���hP�/�9ޯ555���ب#��5��w�������_f��1�@v�p�U��e0)7eb�X�_V.71H�����s��fC�K���Q����[Q� ��3]���c�c�w���DDd����)(��&)���w�7���{�#�)��T��.Vh """�JrL��[�^[*��u���E��Y������j�؀8v�hdd4,iy�������C^gW�!���X�'%*]Ř��:��tg�
V��Z��4���#��(�ūВ�
���h\BUS7���)�y�����;6�+m�"���ȷS��~���	��G`=f�`��S�#`�#���f�v0I�~g�қ��O���to���U�M����f�a����o��Z������3�Um� �e���H��`�1s9�e؇ۮt3��3��a��g�ߎ��k�t�2]�!��E<�⾥����Dާ=[�Ɖ���D?�]*"NU�����>u�e?y �ʡ-u)��OF�F�;z�Qj�ٳ�Z�`0f�2����^�-�vQ��\���G�]�,ԫ�>2N)v�&6Jp�4�M�h��3����N��5��b���c�/�la�3�� }*Ś�=8[\&Jo�⾗��G��m`_yyy())AWWrA����X�!�UF�7���X�U_��ADD41�^,�[��c��z�}�O�|�7d]i���x�d��X����|?+Q6Y�x1�	S����5��3�0µ���}��REp���E���Ϲ��=�,�%�,�n̇Mt ���5����D##����PU�4�[�"��Cʥz�1Ӄ����GB�_��ʤdPr�z��wvv"��z���\/����,Ý�R)��O��e'1�.��
���{���Jd�'��qAK_��*6Z�n����*Ⱥ�MM(A�Q��̀D�tPL�{
Zr#`��:�
U�jk�N��T�PQ�y]���1_|WVL�jj��,d��h�}�k9:�h �`��h����P�+����t~�ۇ[��>�j�oo�N�3Z�A�Q��'fҗ��f}�!��.Ձ�xۋW9!��;ץ� Dê�b��	i�׫����rP�nroiڎ�gkv#�Ƚ����5���J�?^���|��<�,�N_�3S�45tR�g��������n�����uX��F���1�:,?�_������bx�e�Ӹ���%��rW!�8�&,�=9��{�.�-~���k�J����W����?�g[���?O�>έ>�����U���W�g��j���9�߂M�Z��+��/Q����}��O<�!����y��(�85�}�H���0������^�������{���;"��W�����2?��}���ژ%��3��"F2R��8S�G�A(W��ۍޕ�'��xi;�oߺj��Ղ����d4��`j 3Ճ^B���L�p�z�隥�J���������8�\�a�*:�Ј'��?]�t���s)H��џ{S�xcmώ�9"���q�ʴ�kKq9��W��cjU�^�4���י]�6�	�&�D��j�}�[t�_��G�`s?Yt�S�`#k��H�6w�8�܆'"�>]
�Е?�PSTx��P=���ϝ-�n\��������pf�qGlC�U�e����R�[XP;�y%����=���^M^�>�XX��`/�p;6���*E����z�%g��2'D~4�T�>*�0�@ 0���<}}}Z�2Ҿ�n��V�|U|�<�~��_�m[,����\Y̶75v*�5I-���ŷ���'ac�X|�#S�����^kd��9�Tc��h�b:�s�_4P3��Kl�ڦW��KA3����64��G�(�ܥ��}���jt]OYX'ֹSt\�j�"oww�Q?O��.V��k�I�D��������̱��DH/mǔ*s��&���b�E	\�U_����Ig5��M�l�/�l���e�Y������a�;�[3��v���-�}8�x"*�ɷKz����>6�r�@C��Ϝ�#L)�GWȇ�Vފ�]�!�2͋��hx�]���E��]�~~��������W���>����4��:�F."�7"���a�����}���%�C��T��ޢ��F�3l����������Cߺ��߀����<U-�6���F/+4�]0�@4r�f-[Q�!�@���O�2b�O�g���T�ҡfG��W�3�'��?�(�x��ܔ�*1�Ν��tIW����'>��kE�u.UxҶ��M���v�����ZO�vG��'����o�f���SǙ�9E)73d_5h "���7ᣵB��ǗL�;�^��G�.Y%��}b��d�.���b-���~/����f�CO�篼k:�"��'&��q�����*.�ZሷaF���?���+*/���"�#�rǻ�i����+⢪�EQ��K_:���+_�
��hF��D.'���+�6̰YC[��x���[��yُn���|�-?���Ze�B4�]0�@4r�:C�`|*g-���+�O5�gE�X�2�)L+P�����T�:��m��]�Ϋ�4�!:��]>DD�F��V\�	�k��+�v��ij��I��ߖj��x~���3���t>�[�n�مn�@DD����+p�̫�������/��!��Dᦩ�G���w���<��'�MC������8K}r�hȏ����6&u�O(�ݎ������G���U��O�a4��`���+��.j��U�,�dW���35�v�a�/����WD��X6"8M�tsӖ�uDh�u�0�8��׮���A��+4��Zm��u,>LӼ��r�������/?9��_.��OST�հ!��ċFd�@�D#7�2��0�W�k��TW���=�b'J�xZRh�H� ���2� ����sDD�N-f���p�qJ�����>z��.�K�N��Y�K� ��y�lfVJ4q������w ���(�~��qa�)�׼��ߛ�k�_D��T������WGosˆ�A7�#�#B
�z��������l�z�ٽݡ>;0��W6��&.?��=[Ǽ_bI���O��.�����q�,�s�zxL��!��?O�~�ڄ��/af���%�?�zA#�
�U�b�;�0�Y�z��c��ଂKIl�E���Z���.��v�����|�z�&���׾����inHd]��مc���d���n3�[�`���� �Mwz�]t��S��S`S�.t15L��l4�@Y�^�	z�u/��B�xL't�@P�ѣЬ���ыm��ȿS;�<�*�L�+P�F��n��sP���j}8�vc���oGҋ7k8Ձ�X��霹,����~�ϭ��K>+4�����v��|m�z�(���u^M��n�9��5"�pY�T�J� �	"�>D�}���D�A-Z/F�~��׭ڻ�GD4Z�����+�)���P`����k.��:H��-���f��-31(y}є>3BDD)t��F��j8;�����������Dp@޷�m�M=�u�wL�⃸��+�����}cާό���"�7��[ܿ���~'B��j8'z�硽+b.V��#�(t������Z�*���8����p�_d�"��E߁���i����fEQފ|}3��߸����bE�A]%�����f�g�A�|���k��>z۹_���A"�>�������+���ef3d�
d�h���
��١Zn��hP�z�ֵ�]�Ѫ�`c�%��;'4eFb�!mZ�;��e�.�ӺA#3\�!�d(�k_�~�����jt�"J?���T�!����u��Fk[��J�h�M����x�C���{�6�sn�R{AD�k�5Z�Em"�H�>�*TwIHu���E����K��$�t�O�S
>Up}f�T��ȾFW�r7��{9��t!�U̎���a����g�bl��5�6����u5.�9�ל�E�KP���c~=��=��؁���폣%�5����ET�80Ў�����/�'4����Z6���F��Æ�w��Ō�IH�+�+������@�ۉ �n��^����r�����x���<�	J~,��z�S���6|a¾o劻8����ߍ����7�AO<�s�΁����q�4-<HTfxY��&h ��{�A��p���¤�!euz1���с�x�y��l������P-.�O��DL���0_����)��h�y���y�\�O�~t7]���^rb(�z�b�QQ�k�0@������
-r/9!���PN�?������&��
N
�v��h�-Y��C�@F�}o9��� Q���(W��F�Q�`WN�j�����߶��(�����؝��t�#7�o�~3NIc
�"�M#"��Y��Z�"�kn�;���Fb�� ~�mi�2��]���~"aG�箼�uыw �D���_�E�y�	���?��K�B�ڋV͇V�-���²�|)�LG�xk��?�(iɏ�]�x?�拒`'��&���r�.V���Dc{�꽮����=|���|��M�����w?��o��$���e/�g���(&O��a��Tt�gʔp%>�Bty�T9��^68����,�P�G�pEJ�;)\��}�a����~Vl�I�{<�|G7�S9�'�D#x(2Th�U�ץ*l�o'k�?WaF`Z��7;�g�c����Di�xe�6_
-�@{*��2�?\��T��b����ĈM����쟃1zjK���D/����H��M�\D��0�:�0�Aɟ�W��\t�g���|���J���ŋ��e�S=s��c ���j�2Zm{������ B� ��~��`��8bj�G�:t+~t��e���tF�U�����;W�"hTF;�W<#4�0���j�,X��\q�;�����aS��՗��gEQ,��?n�ģ���V��N����@D�����ej��>�`�~D�ajO��K�]��w��\���h1P�ݞ�x<�m�˳	�fM|hH� _�
2D=i���Lz�
2Zշ	'�v#(�M+��G���ܷvk�=U�-�_\ٷU��D@k�P�8?�>8)�2Bv儆����遉G���J��7��{�c�{����[f7�1{0UI��L�STu�R�����5�_t��륷��x��#'���)m��ߺ��Y�z��a��%���ҜDDDtؗ�,Cs�{��i�����\����Mt��yj%�E�⮁��}`��~�ŷ�?A������Hi��ӏ�ٰ5俹Dq^Uf�J�5���V�h13�z�QX���Dt��*�/�*Ë��>�Ҫ�M��?):����5��Լ�t�Zߩ�j� ����&��}�j�$%�c���dXrB�7WD��}�f�^�
o�;g�;Р�jtI���E�Zb��������������^�b��u_����c"�d-1��6����Ap����z��/�z�-OW�=w76��B*���?.������%AuZ��]�G��!<mp�	"""iڳ�Q]�!/oŻ�:y��lQ���M��A劻��o�0���%���7��j���^�4�Mjj���r�ٯ�~� �sú:v���e���L6�M~6FPH�����1l�ჯ�L�z)��=EfBo)���x����2�Jzʈ����w:j�B�یP5n�=�(\�.%5�9�"V)�Tz	���k5U!���W�]j���ݖ� ��I�X�q���rX��Zh����Ӌ��H�+�N
6D��k�KwQV[e��j UJ�>c�C��pN�w!�X���;��|��C�a����Ht{O,�s�>=�I����=F�د��=n@ �9���(p�S�.*��.z�M�<(��f���.��g�F���5����/F��E��4X��>#�7c��(������J��~�fV�)��r�ʴ|Ek(P��T�Ij�$�cy���vӇTyfVK�O��?Qvnى����9�-�[��[��#�te�>LW�z�i�ǻ!��{%�7���r#sb��o���y�E�*W%�L�5���@C���t��u�\1+���"�,����-޹N�wE��ѐ-�$�7mmmG�<U�:VhHL�Qm��JU�"�s��;?+|%J��SҲ/%k�#�}D 8]ǔbÒ�b�&c/���lU�8�K��h�ۏ����]|��W	��V�4v:�u8��a(�ը�Fi��S�)��6�HqV���lP�?��o�X�e}���䡘���h���P��/�@�p���;�G.Р�ep������??h1-Z}�
����K���4*b-���ݐ+4��db&d"Ġ�7|�3:&\�/����x_��J��t���2fT�{q�o~Z�`g���@�,}b�R쳷���ߥ��r��(sb���@0u��X�Lb�7UKlpi���N��d�a�x���}�,X5�J}4zb�9^��Trp���'ޯ�uL��=;�͸L�G���J��&B'E��[�ȷS��K�޻R�Zb�G�S�����F":�N���@C��f�<!	��7�=x���IJ(w�d�c��1�@v#:e�A�5}��ؐ�s�P�g��yo[��O���� �qz)>�7(X���D*f-nk(�����@C ���K�e� �U�E���
4�k�郬^bC� ���;��}'G�ݒ�X��"�L,�lYo�م'�7Ӳ�VI�(��1��vLE?v�a�Ac��M�._�HX��e}���h�L���y	X�я~5>ߌ��+#ߝ��M���ĉ�R����a�Ö��!+�nd4|b`&��!�f`���;�S��y��89� ٜ�7���kr]��'q�OŬeA�@C��ku�x�&"�W���dtK �%\rb(�o�B�!�!�c���31-\ٜw���i�����4_ Q��1w����!\�֣A��R�z���ɪ�DDD�PЄ��2@����/�ȳ�p�a��-��P��G��c����h ��5� ����@ݧ�O�-��Դ+��<\�,d�Ɂ9x�y>%�\/T J��"� �@_�ʰ������e;q�*А�@S�sH��`�r9�X�U��.�`�ab����� #1��S}'�?��B:�����ַ�y?��u���~ DDD$�H��k�A��.�ڢb���je�rđ5z��d7���?!��D�TUE}}=���3I���X�[,���c�޽hkkKz�uz1�L�3�HQ�"�L~ W�����Ř1cPVV��=������۷���Io��pE+S<���L�^�`�X*�RU� ��W&J���'˰e�X�T�b�C2h��\痬�����9�v�h�v_iii��'�A�o����&��*��.��"�l����j���\�7��V߁8���H�F4>�*(%R3����z�4�)���iw���}����4�E�Af4���h����pER��gϞ��A��L�8'�tR4���k�E;��q��T�t��l�r� ��%u[d�:u*�̙����!�3~�x�p�	����ڵk�e˖��uZ`�y6�K��U;�PCRU��o�
���,�6�ID�f�3�Η���XE�^��&K�e�d5^/��PMR�A�Y�f��c���<N�0s�΍֬Y�]�v%��s�S�"o`In"�N��1G-�{�^^1ۣ"""���߃R&u�_��;�f�1� �P�0S)e�7�n<ep�R�T�1а�?5�ۉy��Ϗ~���
\p�غu+V�Z�p8��ӃS��ʵ�����o�>��9�{�8{o��@B!�P�IJ-����_��A[hY?(�R(@����VC�� $$dg�egy�{k����;���N�I���R,���dK_}u��}�P\�<,�j�袋��������^�aÆ�O>1������x'yb�L���N�܊ ����ξ��ne��+�|��-���͍��nsy��/A2Lh8��77�
\_|1rss��\��K/�����|�r�\.S���%�ܖA�Ģ�\DDv#���=�:��_��ų�} """[i����2�E�f.Z�9����M1{SY��g����fG5)}�W�n�on����@��n	Yj2F�J�G�FrBBB���J�?33|�����)�!N���6_�A���⊠�HI櫮�
���G}}��۞������r�u�~�V�|����`;%4�����������؉l+\	��d�%q T2���Ԝt�$^�#����1�$p�����IR���Ӎ�fI�.��-X��t2�����@D������w�����s��Z�͚V�DDDd/c��J�e,�~�O�������� nb�pT{Q-4�֑�	i��p��?0W�Y���]vYP���w�iӦIf^ǃ<9�S�P�0���tw/����[��&�����d���I+R;��&a��;���nŜp�a�	؄�<y�dl��hH����_ )��6Y#\c��ĭ���Kh��+4tl�����i��GHk0��Z�5Hr���7��7���(rր�(y��	�.�5n�E��Z�Q�����lDVt���RG�r����Ր`n=G=��J6�td���z�
�z� 0��"��F�{���?�N�j���T.�̛6m
�������Kh0�xŹ�k$$�JJ5�}��F�3F{z�tB�� �-'춒W�($����够Y����W.u�pU��k�?\)��^�n���%���ѳgO�7����n's7&4Q4+��Z�;��O=<��Q����lf�[�d)k�_��z1�? ����L���³�	H��s�Z�md�k�f���d��o7S�2d��n�*�ǏǮ]�L�Gx�cYbp�'���L]_*IH���9۶mCee������2A(�y3�κ�b�ܷ��y���-��-'���_��h�X���&���K*r��8�{�oQ��رc�c�S��#<yX�݈U����C��ۃKP�жJ؁��M��e{7mBUYY��yq�!h�
�l�)G�C&9r@��o��([Mَ�>�\�_�/Uw�gFs�h�ޝ��y:��P)Y�5Q�B3�Ͼ+�BE";%4��f A3WV̘1��C||��߸qc����	�B�<֞j��ۜ~�鰒�d�˗/�6�=p�//�M����BC�}WTT�t���_ �-'����
-�����]��5��1Q�.���H�̵ݲz�'��Q�Faݺuߦ�'�����@�j�s/ʒ[@$�V$4����
�v�������WC${�6˴�_oDDDd��0듵 �Y��*oN{��J��X�V�� �s�E�{���a;0���.$�o=���#/�\��@<�TBC���x8�����PӍ��r8��D�4�h;hR�$3tW�P�E,
g�;���x���r���(I6��E'"�����3���Vhu��5��&�ĺ^sI��^ثW/��C�}f��d$iqhQ�����"M��	�a�v<w��y��l;�Z<���$��d�j�@a����y�Wަ���&$>����U�n�Z�7�C������C��;�c���o�Q
���R<����~,���ơC�ЧO�����]a���`���&��Gn����v�)���&��Qo�~r���ݺuKE���D�j��D���	ҷ�Wvy���jYرb�� ���}%Ѵ��'��'�_�2V���o�kBC(c��q�n�q�I5C�n�CVV������Z����� "�-;�:�û?wZ���:_\xȻ��%""�E{��^�|
OBÃ��;�������@�e�W��	e,)]{P��S�5�&��d���DYY>�}������7V�������(??�=�����K�ގ����^WW�!C�A�p�SˉD�ܾddd�e?$� ����}7�w�{<^���i��&��y�t6y~H0���᤟��>��;Vh`v���׿[�tt���7�{�5w�8wL��6c�ɶ�<��4�T8#"
�j1�))���(��Ń����懈�Ȇ��Q~
��E1f.�s.�����&5/~�݊�če��S��p�w�A$
WBCII	�9b�6׮]���?�0rrr@�X�z5}�Qc��U�@��;0lذ�$�ة�D����,�lvۉA�5&�<ο��m'"v��Ñ��/p֕�g�Y�]tuP��z%����SP��[�������c1,�>�؆�5�~�wm�󐛐�=�G�������pA�m.�j*J�+���r}U�f\�PL�3V݆m�� {�7���k2��u����r�;&A37��Ӽ�윕�(�I��<%�*�@�Cf5�zw�&���Ȏ�G�%E��	o�����K%�Z�u��g�;�1t�����nAyg�#����EE�Ϥ�����k�e5:���� O<���d�{����#�r�V�����BUUt5���>x<�K~2�m7����&{/���v��+������vLh�B����:6,���p��t��p����������MhH�Kƫ��F�#;jb��?����u;ݸ__��.<�k��o��\��&��o4���6��	6��v��\H��߿&&4��'��A%��AD{�h�=;�1�d�"�3޽�\� ��.4x�
��f\�q1�\t7��#������;�V<�O���v��{��Pk }E��k+����'��}���^�!�d���~:� _G���o�>�v�ip:�Ӥ���BWk������J���v�b� {�������[E�p���1D^��\�z*�k�*4��{����8#�A����R{������T�뱯��8��������L�����G����U�:�o(ns;��o`j�|���7�v��&_�T	�C�(�����nwP��q�cͰ�<HZ���� "�Mr��^�6<w�)|/������r�'�=i*�܌���/�D��<����{�u��P6�C��C��x0n4��67�N!����6�����i5!P�mݺu�裏p�嗃��l�2�ڵ+����҂Çc���n�.	5���ﲲ���GM��`����q��{T+��G�5�gd��$Y���ܪ�*Gh��H�
2���%�֕	g�bY�*�W�	5��-'���^g_w�2ZJ��O���m��m�5�?���y��F��i=&��3��m��NvB*�z�8?��������r��k�+�МH������s0	�D�1�s�p������6R�r���HD��E��<[�xܙ���̮�T��!�m=�Y�W��.�	
4��N�PZO��Z~�݊��Y��f�e%�w;6kՈV&4H�R�����W_�\��Az���;��@{���-m=!	vP�4�:��������Ȱt?�2�Վ��V�}��4}��������V)2ҕ9·J2�#���+y%�B�گ^��$B[=�_��.��h���$�����{˿��9`z�ɧLhh���7~�8�O�q)8'w�惢��ya�	M���K�QB�/2^Ӟ���)�㜡�i�����d�c�~��~��B��b��DD��n�ڻ�w��`��iv3�{/� "���p��p*|Z�	����:�^�s7�StN�뺅���۠h����Mj5~�m�C�ӑ�0�����}�m���AV���O������q��W�̑�{�����ę��R8вm�%���YU���?@�m�6L�2Ų}�d��۷���gp�X��2V�e��'�lݺ����Q�d��hcu�O�y%���!	�&40�׵�����y��b��1Z>L�~&R��h����VQS���~L� I�0�!j���l�I_)6I��zl��x9�S��'��"�Ģ���w�y��̫M��������Js�W�Mx�y:F*�.0����{ �Q�-� "�$�g���/	���U�1�������?7�t�"&4����'��bֲ�^-؉:/�5{�0�����nJZ�ƻ:G#[�^�T�|��n�~-��%[Y�AV u�ŋ3�!�ׯ������B�~�� ���Тxp�Y�A��W��ر�G���J�l���ow\��TvǕc���ח���b���V�&G�1u�]��|�$��&X]�]�!�%�W�ړ}���j�vlF;�� ��íz��l#���\\��L|P�������%99ǎ&�*���7Fvu%�VV��ƹ��)��W����FZ��3YYY����ݻ�y��S�yp�w�s��XŚq���B��޽X���(�I��_����_*\�&�!+>�Ӟ1�_��Q��0��L�m����;7=�w��u@�=����o�N�|5�Z�h(�vku��w#��y:{�u�B���x�4s��"��춊�>�V�@iII	z��	
��l�\���Us�� vĕ�Jh�J&�~�)���
8���kך�O�/E��fĲe�p�5��2����/7���3��;�B��=�P8|��G}0}�ɼ�{M2�~T���댄��{�TBCߔ<�ki��� ٟ��y�J"����7F�Di�_���n�R��̃�$4�x�ҥ�1cFȿGI`]�j��ۅ2�#"�6����l�ϜC1�aM�=�#�|Uw`�Z	"�X2�hJ�;��',H����ޯ�� �2�R{��D�)u@�1k�<'�,й��Y����ׯ�û
rC�\�֌_z7�^�(��`qg�W��{u��'�XY�A����5	;w�dB�I�½+���GeB�	�0��4S��D	�_p���+�$0��G�����};�p�| oc�����?(/�.\��.�,违<Ni3#�#3�76�!ֵ��?_�U��}�H��u[��Ҏv�	i��;
�Z��:���q�Ć����7�����a*�& �;�u_IUTv�\HLL4���k9�+��\[_��UM��������I]tQ�ɬ�\�y�<�ͨp4bFDD'�B�߼{Q���z� Sc:�F~��{�a�ƪ�D{�5+�nQ�حO�����$R@:?�u�ǅ�{�P��?x��/e���n���@�t��d;�4��\�a��eШcҧ��jf�-=O0]��*V&��)���Y�qU��6u;��!�/��Bӕ�=j$���	�E�����"Lr�3u���"̟?ӦM3��_V�.Z��x�f�O8�}Ii���T�������[N�l�I�<��2���=&!Nqbq�zx�c�R�;��������%�g$D�$G������j̥��o�.?����o��Ϊ���(m9�k\�8��Qg��U`������߿�x�������Jc�L��5��϶DDԖ�����G�ǯ�#����C�ڪ���T�\r/��>���Ph,3ZxJn�+)�)�vգ�9�D��Y�M�@Ys��Pş��t���SV�hO�-�I΅Sq�pS9<�/h"�U��
�ZX�t]3+��ɇ�s�O�s��bsX�?� �P�;�Ñ���x��w7>W��1	��� 	]�}Ia:�PVd�BZ-X�n%�%��͞ɦoWXX���z�'O����OT��M�6a���A��Z�'�G�%�2�� ��ʌ�;q�D�9򔥗�1n߾����W$
�%�#A��	�^̪e�-'�,�.��Xc�Ta��&Z����0��d�	��Vyջ']��� nX�((��{����l��f�����[�K��	��d��+q����d4��\B�8t��Νk���z�y��=d�'s�`��nŋ�	{ADD���*q�g���l��<�����1��(0�� �e����L�M޶�\x�='�όOţcn��.FZ\�q�\���E���v��ߞ�\��<tK����e�Ǿ�����=�8�ç߄��O���~ͣ�u蕸cص_V�|�h5f����]�G��������4��ʜ��ϯ7��h�ё������9�Fa�G�by�<������6�f�m�zωH:޾��3��G���:�-�{�cz�[��:�Z��%�.�v����%à�WVmr�Z�]Z�r��h%d�]Z-��D��\V&4t%+��"����9g�^��	�pe�(�𦛾�TYX�d	�����v�޽��Krr�Q����8x� 


�
��4q/���8����b��6�sT*u�\�6l��!Cзo_����WH�\V"Jk�}������!�0���W3F+8�����+`&�}�pV�a��~�:�"ಞ���K���L�v������ަ|���M��Pc9(�X����ڷ�8�J��}�o0���r�;�f}t�Y���L�%i?�n�:cԧOdgg#))ɘ+��[�}R�!�yߊ��:��s-Q���	�y���A���ͪ������j�폈��ʈO5Z��%�'O��=K*���o����z#�or����30,����U����1������c� ��*��S{�Jw#�@��L_q�II�308�4��nǏ�������}��$��\��݈���/��+�؏�I���,^y��q��ޑ�'�\��q��'C�0�����
�������cqA��I�Sx���~��Ȏ���}�3	��49���F�I�� �-u���6k�o0�Y�c�6Y�5�מ͸��3���d;$�!��z�{2[8]Y�?3����X'�C�#,+�'vj9!����p{��AoC��_��8�C�Ҍ����V0'eF��@��$O�oٲ�8��GQ�^
�ҝ�_ir+�������� ��e�E
K��T���|R��%fbs�~��$�^V'��m���8u����K�6�������07�s����4ֳ��-�*9���'43�s���y#e���^�7۸q�q
�Ņ�I�ADD�q�����z����,ث*d$Z�U�	�nT��QP.^vr2p����￹�~|Rv������M���{��t��T �L=ㇸu�\�c��s�I���К��E�.ܒ�6T��&	3�^�&��Hzx�̟?�eR�L�>��~��5�6W�����]��L0�7��2ܹ�yi:V1}l��s���O��)�}n<��3�;F2�\����O��	B�J��$YB*2�cȯ�c��{k3�6^3�hSq��������+�^�P���ȗ���S�^)���X�Y�>�~�[���Q��9C{�r�4��<�ݍ�Zl�.�z���r��!//dN�=��_�-!!V�[B��_��	�1��v4'e#�$�:�v�7�;� i������*4�W��.+y�=I�+�"ȉ�M������cs���H����s�vB�(.:���n��T�C��=���ڗދ�\����Fi��}�7V�\�(�X�r���h� �����*s}3��DcΞ�r�I<��[���Nތz�DDd��7{���p��'�5���� �%>W��*	��{:�\��uO~�D�G<.]~;��~y�, �c�F[�)=�v폡<r��d��u�q�_�Y4"�o��8��ٿ�]�Gv����'ݿTAx~�ܶ��//�����Em���⒵���?�y��X��X��֔��}��.k*��~�+)��]����^4��DG[j���(!`~{�wq���NA����%u���|=����&܈�l��}��M���q�g#f:��:g$ �K��Ьy����-�2X�r�W���0b��9��`���_�e�q;&4�WR�a�'����_$�O�`����c��;{ra'���(�m�ڳ�����[�l�x�'4�������r<��/y�޾ʂ��=��r�gzϳ|&4���/��>_�O��%���M0-��>�	_�P����)��8���Z�z��}��'I�]�X ""
N���_�{�R;��;����
̧Z���G�ƪDD�I�SI��3�?�V�Ifh%H�/Z��7�*����g��0�߱��O�~�gL1��2�e�葔m$G<�o�Iב䄇��о>����o�=��.4Nq�zbB��NC�#�hy�]s}nW0����FB�e='�oQ� �G0{	W�؄="_��1g淡U��r����j�2a�Z����p�#�Y�~� �B��?=�Q���)juBCFFF�'4deea� {�������c޼y�L�B0=ݺ��vMhhT�x!m5~Yw⵮/�/���+������B�j�]w	��D�A�҄��V�Fm�J���>b����Kee�^�ҋ\UU8�?Y�=x�Q�8�ޏ5����|,1Jz;����YÌ��A�)Qx۰�qy�I��7�U`����W�9?<�l�?P��W���X�/q�_�DW�(Y�LB���/�s��(�3e5�D�s�bG-���DD�|�
7�_�
Go|�9 ɰ�q;8�5�9u��;#""����2v���:;N��@l����z�&'��q�)������|����1����FBC���V�-58�TҾJ2CIs%�&��CO$I
bU�v��U���m��94���$2<�YKن}f���zq��7c��&(����E���Gj1~��ኽV�t��Z^�_c��	999(**�|��:u��g�y&233QS�y�9��-'ZIu��SW��¡umbY��O�Lg� \*��x*m9�Z��mV<�{�
T;��c���T0	�P����mP���z����@ߩU��
R	�¼3�ߢ�O����^FAi������E/}��o�o����>f�>���xF� l���~���C#���.Ž[_2��6CMh𗸕-'�$(dgg�_�����U�9W�g�V����!N���%���7}Ԥp��U<��z�iGq�c .vt��ȾT���z�8���%��:��l#V���9��?���{�s_���B�~)_���qY`�>�|'�h(E ��g��������o���JB\�c<������	$�@�r;f-�;�V������0�����I�Ic���-Zn�l�8G���m�b��D��@k�k��:���	VKń����Ɩ�����A���nƌx�W:�>{��a���� 6��_)kpS�Y�P��>�l�_Җ��������{�
���\�h�%����p�pH��M�^�o?�[�Аb���Ⱦ[������S�$�;�]��O���5����Q�_?-�d$@���k��uQi�Uf��Riaz��'4|\��͕Fe������ׂ������I�Ih�m;�������Nmg\�OY�5��xtM��JG#���* ""�Uh-x»��0���9z�tbC���[�a��-�^�}�`�w,�]*0����mN��y��֣���j����*n
,���m�! nĬ�o�lǞ��Y���7/)��/�߅e���
��՘��ŵ���d �l֪��0�Ъ*AK�QI�w�ި���*�_~9z��	
�W\��T�=�ՄT����ĺ�ChP\�q�ٝ�/����i+Q�t^[��qG��O���j����(w��%��m{iZ+
44�vX�W^ة��-6�KIau�@�e�;�e�709g$�\�G<��-�탔(�y����B�z�;�U�#�z�7�/.[����Lh�u������I��r`~5b6~0�2&4D_��ذf͚��!�	�vW�?G�5N��E�ٔP��8��R�Ν�:�X�
UDD�W�5��=�����~��莸Jl(�Z�zj%h֘�@D-�\ǎ�J+ϩ�މ:O#�Z�:��?.]���#�$M+��\�o/Y�%�F�f/������b�@���G��iJ�q��%��V��*V�xG�`����LR�V�����z?�8q�7��'�o��V<���a�	0���FBB��_��2+�{r;�>?K܏7�7��t~��#�<��1��8�]};�>%��R�Z4��r@|%4�]�+"�׺�-6|=^�5��?Z�g�|֯�^���O�Ȏױ���ąsrG!+>EM�Vs���R����?;�4��aG%O�R�B#����S�-1G[ؒ,Z�z��XW__U���_�VJ��ZN����v�M�w.���8Ι�'�(J_��&c��[����x5%.�A%"��T�5^R0��Ǩؐ��m�N;�Z��-�
�^.#"�4*�����1�n[�W�]��ʩ*ev�����=�X4��w��H�jܵ���B�m�;�5s��s�$����WХἫ�����HS�p��gL�*�:(������Z)>���l�J��(�������ֆe�������m|��L�<�^{-�~��l_&�̐��h��%Q�ሌ�,)�x�RLuŌ��H��s���Y�7R6`[\	���m~.u&��ŷ�!CO��G3�Iڌ5�Y��	N�����/9�#�� ����4��!n�@�9�\�=�Gp�i�aj�Xdħ������xj�;F[�I����˱�b�)_��Z�u����R{�ʵ����V��{���Ԟw�ۍ��e囿��K��������/-��͕��ڗ9�̵�?.��3�'��T�s�U��?�/��Z�ڦ3��y�T��y������ź
ͅ�x�[�)J..q��$%'*�Q4��ej9�Eا��QW�q7�'q�J_U��U{p��q|��C�i넆�E���0"�.�1��ײ�jL크�X�̫����߂�V�����;�A\����9F������#���Ne���Z1>P�1@I�y�n�H��JxO�R��`�v�գخ�2�eB�$�=x�`�ٳ���P�������>Y�{����&dɒ%�o������F��+mG��aI��'�כF�k��HЬ��
G#>Jځ��A�We�G��2\�<�C�Em7�,Iڃ��{�̪��
N�*^��k�5�kկ�^*�؅U�L���̔��H�L�\�͕�瓜	FB�?o��8��m�Tm���۵j�4c֪�@������3��ʓTۺuk����㍤����}B�̛�:묀���k��tǹ��;�T̒*R�6���-���YsH��ф�wbER��YNDd}��L;��<G������s�a����Vs��-�j,��b�ViT�%"��#�(%�`PjO|��馎����T�r����+{��{G]�����3�&�k��sU�vT�:�B�;GV`[m!Fgċ��¥�c|�KnB�QqbAq�����ʌ�� ��=�"�i���.�Z�<("�?�A<�����7.���*eXg����x1LI�DG&)��O��Q,eͤ��:�
���^}ߙ�-��%�5|�p�r+����{��СCA֑*��~;�����;�X�M��8��f8EJۉU+Mx3e#>Hށ�Z�c�{ �y���$qa[B�QfxS|�>6�� C������X��\}1�5�(�l��EF�]qeX�x�H�h��U���)�Ґ���v��Z�S�6I���H�5Nd6������ ��t��@��*:�Ղ��~ٯ���6�Ib�����V�BS�4��M�0Q�����l� ��ގ��ŗ`M�AlL8b�V"":�Q��{�㔧$&*���B�QA֩�Ʊ�MZ5\|�!"
�&����+j,�՟?��K���!3pǰk0){��A�zl�������ʳ���yg`V�𿣿������K�����I��5W���)=0��$�A�e檇�b�S蝜��i���i�&7U -.C�z�
�z�Ǣ��'%4|P�����}�C�%�-7��-�������4J���Ŭ�{A�~�Ŏ|{��w�X47ݧw'�t�2dIح�a����і�t%���юSґ��-�.����zl�j�M�տ�%���$P>d�����ȑ#AoG�cS�N��Cddd��'��o�cƌ��+BږD��f�=Y%�Z��)KK�wyr�ӛ�<5)Z�Q�أ��͊u�f�:�Q������w4���RIaeb�qJU0������K�7�Z���j����x[�R�ŎZ싯��24��%��de�	v"c��'���os�U	))\�LdW��:3m"����3���'~��8g��K���L5	#<��y_z���}��(I�3*z5�m�K�u��}��o����ș��Wʵ�crQ�8�Õt�R2�㭧92���=�!�jǎ�j�ت-�Z@DD�'-N%�G��ny�H ���vm�Zݵ�y�$>��5�`g�!�9b&&f7N�l��oT��*�B��%�/N��HL�q�Ʃ�Fo6��;��?�~ۨ�p]���=�8�����!��I�s>%�O�5���"Ld%4���o0wڻд���t�.H[
)/����\'�Q�1PI� ����$��~YV��*ͅR��D��M(�'�hD�֤�5+0XM��f�fd�\}�ո馛@�7nܸ�$�dذN),c�������NN�@�w���à��/'�gR^=P�z��q%�<��	�Bb���o�_�/���lK*�Hrm����.��~�v}��J<`B�=�8��V�󭍑y}E*�l�j��[r�����$b����HC?��q���$f�K  �IDAT�a�դo�TkF�ւ"��hk�*�-��@D�i�T�4���W�jw=�X�;�B���蕔���k��NHf��?׿���w��|a�O�����T?���xz�qe�)��3����m6�����6�7�|��?���(k�b�\G���ug�c�H�K�V?�$�������䜑���$�*�Tg8�Rc���T�K�I�I���>���3����r��8F�vn�O�%�A)�Z�\�K/����=(y]�+���>	��r���Y�>Tf*�HG��ܐ�O����m��oФ`��zŋZͅZ}:_�y�J�y|�����X�O���)�lf�%�NI_�;_�򁯄;�|��{iii��𗨑ʄ"�j��Ҿʂ�
-555']��bߖ�I�p�}WA�8GV(Mn���D:�3r>CG��i-����,h��(tZ�q�GU����@�������Z�Q37U�k��^�4͊�:͍Z��㬬nKDd���1�p9�P�\e��y��g�����"�t*����S����S�d_	�I�D �T�4N��pբ�2�� �����f-�7(�EnB���Lf��cΥo��д[�(���Jvo�>/�	�N`�"
���`B�9���f�$�(Rz��z���ѭ[������2�Dr��X ���	����ӧO@���8��d�M���2O�1�T|=VI*�D��I�
�Dd�w^U�(RI5�*����m���;���DDD1J��?���nZ�u}@�2�q$f��J�������S�ӎ�:��Q�DK�	����o��L�yٽ{�I�۱儯�$(�x'/i��v��^|�N����f9����&�8�	c�<޼�S���r���m���p'=��.�`E��Hhhu�B)r;�L{
��(� ��@)`Lh�h�U�D�� U�R�򾐕����UF�c��_����L�$} <�Ϲ]��D�_��ॗ^
z�)6���,X�69�9	��5DDDDDDD��ie��G<��5KX
/
Eg�k֢���0�� �-Д[�` �N�	X�(8�j�� m�/�������<�@ǐ�ړ{�p�2��cL�k�_�CH�*_-r��q��{�q"""""""�R6CQ�A��e���nљ���X+�?��������д+؎���+4�W��}����\.���1��_@.Ԅ;>V"j�ꀼTuINN�ɾ�㭫��l�爈�������&%�Կ��ٟ�ń؈z=������qz��,���?�g��_�������
d%"��+�׾bCGZZZN��uu����IRF��I_��\&�?��IIIp8�+&4E:���>e��C쉍��]��Z��%�4�L@�8.ӿ�SPL�̄9�:v�ؠo?n�8P球�?��O��|h?z��BQp|�L7��PYYy�ev��8!��0������y�����������ש�_�2����Z��&nu�]д�p|�z�r&1Ķ؎z�Z,Q������/_�sm��u�~i��@�ܡ��ur~���_��\<��+H%}��Ș�+`f�@�<��I	���0`�)o��D�6���d\�y�U�����3_�jv�i�Д��׵а�J�ZV��b;���o-ٯ�/��/� �C�zN׿(����I�M����P�PUD���.D�����w�J-Ҋ�Wŕ��f#顩�餟�9�A������e���Ñ#G�Ĩ����8 mll4�/�ٟTh8p 


,�����ag��7o�$�#;;999��Zl�ޏX���������,ҤĪ����9(Q U��b�bkRP�bBCG�.����<~��s�ѐ�����(b���Ǆ,�K~��;��Q��k91)c�28��(�}�ip?�˧Vo�_0������*AG��О��6N��d+*4�iJ�>V�Q�;�y�����±���?III(**
:�W��F��!C������0m�4lذ!�q\HR[�=0e��Z�Mp�}�uG���y%���� C�Мրt�3�7�(Lh�7?�;~�
1��y'���Lh�h��D�#��x%��6���a�%oev�j�V�W��,��P9V9��
��i�u�y�!VHE
9�I��X˱���������Ԙ�@De�r�(8��˾ZG��+Y�la��""""""""""�LLh :��(Z�k9AD�&m'�LhH�����s�Q��5?圕��������b	�^D���0E&4O�����nϮ��7I!"k��ןtY]]���������b�^DDQ�ID��ׯ
-�V�nݐ������5�*466Z���}����u��A>��e�Q�`ċ�8Vh�h���9���ؾ};�^o�ۑd��S���E���^��K����&��8�N�; Y����Hj�߿��}YYv��""""""""�X���qLh�h��H�ʔ)�<y2�nwP�p8���G$�޽;fϞ�����<Vy�Dd=y].\��6��������L��r�$��F���cBE&4�F􉉉�			 "{RU{��E>��1b�8p DDDDDDDDF���cBE&4P��MDD���>3Z�������������È�q�Q4aBE���F��744���Ȏ��FYY��������(p�x�+�a�ΝLt �IKKC�~�:�(���V�#�s����8E�/�ӳ���(�r�)1�E�Y̄��@���@Ѯ���6m	��e�^�v-�l"���r����0F���c��	(���-&�w���B<x��{+�Q+F���c ��	(VHk 9Qdk�)�v�QQQ������������Lh �(�0���"������'����.��o�DDDDDDDDDDd`ċb����g��]�HZZ��&�d&4Q�ٻw/�����������NĈŜy���onn����*40�����p��:��� �V�xݬ�>E%EQ@DDDDDDDDDD&4PR���#���T��)r���t:A�n��b�˹ """"""""""��Ƅ�)��Ͽ^Ӵ+=O����@?�455�ӿG]]ݡ��w:���/
�lDUզ���b_?S�1++���կ���g�E���ܧ���*�~E&4P̘7o^7UU�T#?�:;;� �RK�,9����V���PRR2zƌW�������������(�0��bɟEɓ3999 �b��������՟��x����}�W�""""""""""""����	��ϿLӴ��|bb�游�	 �b�.##cxccc��m�~��|�d���� """"""""""""� Lh��7o޼UU�>�j�����@��W�����������|7�����FE &4P,���(��LZZ�J��q�~�DQL*4��u�Hr������z�ꯃ�ϛ7�3f,��1���ڼy�&)��s9�p8�����8��E1M��9.U�rssk���Z���9sN�5kV=�������������l�	��.]W__��~�)�gggoU�<M����z����ɓ����_�?��t:�����455M�_���Яr'�������������l�	�����ֿ���			;��9��-����ָq�A�&L��Q~~�$񼟑�ѯ���Q?��(�/�͛���3V�������������Ȧ��@Qi��ý^�=��H�}-++˥_����Oƍ�Q��0a�����)�s����`wUUՅ�����[�n���""""""""""""�%&4PԹ���^��EQ��������c�ĉ Q�0aB�ƍ/�_/����x<}���(..�� �1����ĉ��4��~گ(�;55��I�&�Q;vl�����'�|�k��}�\��>����_���ˋADDDDDDDDDDDDd3���0�9��    IEND�B`�PK
     �)K[��R�(  �(  /   images/d39a4f5b-af2c-4f90-bee3-bb82593c1b3b.png�PNG

   IHDR   d   @   ���t   	pHYs  \F  \F�CA  (�IDATx��}	�\gu���ګ��z��j�$˒,ٲ���e���16�C C�@�I&���dN֙!0�C8f���2f�A^�U�$������R�����m��U���-�	�N�^Wջｻ~������{7v�5$��r�{WH~��]����D	�eH:İ]�T���5z�cK����1}��+t���ε�tlб�K��@Ϥc�"�Ƕ��F�WJa��wX�����Oqӷ�b�hV���C�¶��c~I�8�m�@����W^�ྦྷś��sJ��=��eͻ��"���wɝ�K� b�9lzN\�.�m��V	��@�g���6��m���H�~�fC�H���.��O��{�H�.`�A���MU�$��z:�K-OO&�Ǻρ�&����5%�S�����xDZ�;�.�xf�]r7>c�K���ǰ�)3���}�r�Bv���v��}薚�sϨ�,tY���hq��[^K���Ct�狑�lQP���(��$��m��}�VjA�+:�������yX���~�uR���,�]ֆX<��k%lXߎ�IO�X���G�PȢ�W�1rp����~|=��� ���VF`X��E�����M����$z$��mE<�w�]N�N�����CD/�Ao���n��w+=(��=�?�_"6}��*���C���J)�ٖ�K�?��&Y�f��0)�q5��d���߲�T9�fB��B��G̙�	�q����EQV�)�b�Ԅ2�r	�� �ڥ�4�{d��jS��MC"M�=2��L8��p�x�a������/L�s�}�XFv��-c.Y�<i��Qpj6#����V��9��w�P�w��^l1=š�'��-ay�a�k���F
��j�������&��4�t�U���6�?��#��Vd�c]���'����������.ip��mE���KM2�\>���Ja3)"B�WZH�Z$w�ȺM��¥��%�Mn�ݰ`�t�VP"�3q�KE��c������&�c�\�"K�:VqN#=�J�L��KHg�s�pL� ��=+k�F�;�X���ێ ��KB[��-��y���=��`l�Yv~ �`�^q�����x�r�(������j�.�e+�+�f�X��)Y��^(�=�,�f7��e�?<9�E�@�q	�Vv5c�t��Ī�f&��eCt<B�&��������"a?~G�R���$M��K.�;I�
�H/H�z~���__��Co��ZBO�Pw3u����q��VwI]d�ߐ�n�e��<�o8FA���!�^��B�&a(� �3b�i�X�v�;�Q(���Τ13;#bE�R��oٲ6l��XS�~~`�F���6��o��2^����>�Qx�t�4H�S��Ir%<�W���J�@�I�ԩYd7�}�6ff�H]�@-똈%���D��w��Mgă$֫HR�0��}lV���=	�f	��1�'Q�03�<=ы	z��gz�e(Č��
b��'�>������w���s�q��)l=�$�K!ږ&�1d�L�����E���c��J���~<���hmm�W\QEYt!�0�?���kZ&j�1b��aa8҃��u�c�����fG;��\)��Q���?	u�f�k����U��)WuL�7�����/(��F��\�ӛ>?).�m�T�ޔ��No����+��@O"z6z�<P��.�8��1$���ˎc5���r	���a26B���TI�-J�Ix���r�֙���-��"�L�-�b��"J�R�B����bŊz\R�8JB��3�1��a|X�%[ǛYۗ���̂�VE$�Q��k��,F���3�Y�-� fK	:V�7'�{��f4�B�̗S���q���R{�A?�U��2�::�vw����:�µ����v�^y�p�⃏ �A�����"({In�t��14X��ķ�B�*>L1d�;�"����P���z�r���X8��Y�&q�Da�Qě��A��?��o��C؈�3�$��k�?=�&͇%Y��=��f-����_� c��F�0���涍t�8"$8�Ta^X�9bXQ3Q�P����t-1EH->T_�x�sdvAG�ۿ��>�GZ�������W��Ǿ	�,��Ʊa�֭B8�� Ԭ��6��[���C:�RUe�X O���W�''+���HT2H�Řd� ,%KB�u�Ϣ���|^d�9R٪����Lᤆ���}*�f/&\I��*�Z���Q���(Tӂ<S�̞ch)y��X�*M nr�����e�&�*�]�Zn\t�8ÆGW�*(,<��Y�Hn|!����r�Q�t?k���
E! ���Aoc��.�u�[eJ�f[��<ʫ�m��0���d��'Ռ��w<��v�L��Ǫ��d(����eQ��`vv����ep�\A]!0��p�����-���Z��<87|2%I	��0��ŻƧ�e� t�w����ڮX�-"�N���Z"Ɵ/wlG �W�+<��@�nT�処i�ET�)t-��X�	�Zz_���Ep��hT��$��L,4�ۍ�/����B0�F �rM6B	-�^��j��}5�I�z���C"��j�x�J,��	�H�Xϡ�׎�$Wg�+�
Ʒ�����ɪ��
Yנ���N�p��vCxb
��	/+�E�E�����ݍ���%�������<�����A!�K��������g1B�9�w�,QQ�!�"M��8��9��܄�:��\[b��=f|�~�8Ŀ�EeB�U/���G�]�R[���<��}�2��������x<.���ZL�d)�(��Vq���]�C8��ȑX]�*=S��d�\+�7�H��Ȯe3bLcLp�5|��+��!&.�5{i�'��ݻ���"f�kb��q�������G1D�s�K&1j��%q*G9G��͝[	jk�}I.E� i��N�XMs�KKo��]���@���AKX���^�����2-�R�~��^1W����k$�k�ڊ뮺�K���F����Y��j�t:�{irI�]���ۏ�ˇ�Kc(�s������
1�h�D����v��S97-a8[�l���hm~l���^��%c��
��t'�9K��ބ֒�ӟ"Hl8�Z��ǟ��^�w����s,�m'K���X <���y��Sƾ����WdDD��iѯ��B�9�n�%�{��8� >��*��)�Wl�ucܚ�xi��Θ9���1�?��z�>�/��Ԭ�~�Vk%b�~��v\�1�2��%��g��JIH��0	P�ߵ��2�nڈc��v�W"��w�=�uh��T���Z��y�ِ�Y�ov���"�W���>�}AC&~$`KG̃d���ZKH���d����w5̊)
��@H�i?�n$�:Fù:a��-��l-ˮ]�!!�^���B�D���(r��l��<�ʫ⁧ۋ
k#(yE��BT��X���y��/;~p�N"k��~.��&[�Z$��H���(x���5F�^��	��E''��N���$�=�zk���\���q��jv���E�
=|�_��34*����+��uK��i���28vTEȖ]��r5��n����T��r^wY&]դd-��I>�S^`N�mJ�Q\�6-l���~q�ݭع%����#�7���ȴ/؎�����w(u+(㾵}����(9�*.�]N��V�f{�#�g���I>5C"�,~��#̘hH{%D|�{�GB�-�G����CQ��Zrkk�u�p��7���0ƶ�#�0�#�r�PC\�����}�v��kDS,Q�S�������J'�WYH�H OϽNy���&[|���Ϝ���*h��Pa;EK������I��@��F�h�h�B�l�H�x��4��nVq� �R��s��T�v<<Q�8�Lcsd��$�z�X~�B�.t4{'�7sUr����Q���D*V��%�:zk��1����)�Z���S��:�z�9�I�9�K8	�/�::�����,G��V8MtKT�%m.�)�H�ֆ��}v�|m�`�6�h�E�2��\��OT'�i!�/�.%��%���^ �y�)\zeJ6���I��izϑle	�B;��U�m�E]������݁��Q�d!**�׵���Cw�P�$2F#�	�U�9�.�B�r>�}#�țO�� 7�����zv�-7��e������8fb�iSčf�a�!+[d'�xU�^H�
=F�b���R�snՋ�Qk��1WJ���a�߁�_�[���v������x#�d�w��(�t��qw�u�{���k�,����*���뵤=��u�����Ks���IX��}�e�`x-I]���.�!eY"�y�FS�՚�,��|�m�E����s�w�y��Sg-Е4�
=!�5�^|f��d��B�(�c�YL�'�K �o�8�뙃�T�GY6+���@�w��Kq�/��hî
�l�������u��bk�������&��y�wun���"�wz��+Y�.�t@�b�
L�)�ǲ	����<��M�X(�DͲϳ�O�9��B���h�C&��>\��;�O��$��)��f��9a�T�BG��@n��.�P��9
{�Y���,+��d%�ӹL�����Q̿�c�kޏo�E|z�
�?U�!o���X	o�����y��	�W <�va�Άޤ �i�f�x������`�N��:Al�"DW%���Z�N����$������wuve��Y�S�n��+nq��A�5ж���$�(ŏ�侾?��pQ�3�IO�������'�.3��gݘ	Z՚��9��\!�Ǜ*�3cX��77��D��6]F����.0�^��^��1O2�t
�����el���IQ�Ad�^Ry�~t_x����iUl[:�j����8f\Ӳs�ni�D���_̾������HIt�K��Ħo<tya�Y#C���$�G��RZ�r
�H(����B!��>�˽q�l�0���4�'s�T<� � �~��f4�^'k�m��d=�"d%S�9|���8���Gv�k�O�iT�-�\�B��	�FM����yr�BI<ԇ����(dm^k�)\����<n�C1ã:���ߵ]n\?���)����
)��(V��(�j�����?�:��ۅ������D���L�;	s�1��n���& ���@�6�y��� ��u��N�qlA<��#LD�:�ć{Q^t��v�pe���^M�U�w�*޹�A������*_��B��2�t���ږP�e�%�;���	��,��v%Bm�����zdB&^ȑE�#��7݁����4gc��W�����x��7��]�A��۝�g4˷J�����&;�I/XG1GJ�S�z�:���xT�Z��u�͖)�ٸѵ�s�y׿>��l�4m�*�e�����(�ݞr&�g)�g��b.w����V��7P�t_y%��={`�M��1�˄q+YU�tI�L.���[[��t�_J,�\���=H>�Cf!U��d5�qԘ��ʦ�g �|�<���h�P���d��O����6s �w�&(̫�TY�"��PP��Oe���Y��*	���������<4J��URQ����������`^M}�[��(�2�{�m��n��T􅉶��S����*x�x
�-e(Ѕ6w���Xn�������3x��ضmT�3��!3J����)X��1Q�T1_����;��;(1���Iea�0��H��E��B���.��Q��Q .��LyI��,\�K�tQ���ԃ�N�ń�X�#a<L��r!r����ȉN�T0��N%��WX�9��uOr3Fc}��w�w�釳�D(��6���H��?҂��Y��f�l�0�~?6�A�'��#薌 ǣ;��W:=��<���]ۏ=�)A������~��K;�9
�RRt%rMa���[se�L��>�}^�5�y�S�Ͱ�� x�a�(�l����T��'�(	��T�d�;�bn� ���!��rX�?j`*hb���B�
����Wz�r2���1�]p�M��:��N8�bӏ){�ze��w�)j+��3�ٵ��4Qr����;��K.��C���������ߨ�����8�ĉ��2*_�-:�-��j
��N��?g�1���0S��~�� �Y�z5�̬D�hm�{?��Q(�z]nQeW�?.��A�B\AŇ���~�)�\D���?�/����FX�<�y��'��])��k*�'O��T6J/Wz���o����XQ���,�$�Z���+��Ќ�l�[#�s���!�%Q1t̓0�Kcg48�6v����)X��͐��e���4+��eZ�©' ��(�F���(����� 㩈��7yעE�qs�kYΫ��SF
���4h�2Tglye�q9
���y�1�;�eܨ��޽8�%g�n�4��NN�Ɛ2�����ړ��B1_�Q1p~�^��-��R�������1�90+cS�	Qw	O����z�QF�G�k��H�l���kӘ@�@ˡM����ҳn����yY�]��0�mdK�*��%@)�e�U}X�l��c�ڇ�$^���D��j���/�&���#m����W�r7Cg�2J�Q�q>�LL��UF��q�53+�P!�4�~��"c���v�vIxFN�fk�����&E�m�ʉ��R�Փ�n5)H�]_�
�f)^�A�=��j)Ģ������r��n�R;�����;�p���X�eQ�d5N%���
#_���cQ�^U�U�����	1��yP�my������S�qݞ?~k!�v�rI'�8ױ��A�YX���'0�ʷ���n$����"@�b��?��|ߍ��F?��Lz��,��M
�j���1�e��ꫢ}4�N���B�Om?b�\]F�*��k�H�^T*.��=mK����.�z��ڎ��x�me"�l��@+�zbO�B�ii���'��*^���2�y�ν�kg��/���R�IBm��_� b����b�h�F��[Z���Yc����wR^���=���N��(�eX� �p,d�ڵK��mmm���2uj����z�^Ks&�Ȅ^�ʯ�Tt���Pɻ��o������ƛ�&�i�t
s�(��f���G���r�L&�n݀c��bw�;�����ٱE�pbZ/�`Kx��F~j�el�A��&��@o��2;��b���to��JC�,�׽�-�k7�0ķ���>I��&��Sݘ1RU"�� �7�ۍ{ｷl����Bv��C�w�'H$�7�h���Ꙡ���v�G�.���O��n��N��e�KE�κ`�1��l)�	Ç�6[4���y565�xn������iq�k��s+�`轢�p}h��鸷�&�d��,&�&��4��u�Xf���&!,^S��p͚>p�i��&{YF������9�u�NK��zb+P�\��\WW�[GUP9U-�\#�)�*bߠ�,���B�Z� <�
�2�� !��frv�j�J�%��R1r��ɶbU�3wIvn�͜����_;�<�bJ����N?�����}8�-�� 7m�?$�S��u��B�<k{��D6���9�D��[�Uäh[�(Qkrc�(�VD Ul�OdQhS.�@x:�qP\q�����;+�+�z}�"�RY�#�Q�ʗ�ؽ�.z�����=@5 ��������	i��岈���δ���|��v�a@���?�!�K)|��3hu7��������
k�1�͏��	�j��3��g����#��e�6�u���cyP¬^Db���J�S9Q��j�o�z�: n9xK��6�	�?Պ���N��;CY-3��*��z�(�8�V
���ͮ���o˓:�eb2?+���G�����q:�B�m������`9��\Ηt���`����7(7�g�"G��^Y�����6	MI�'h�T�ao�J���%���)aI���d(���^��*�̴�Pe��9s�W(�P�7���l�����_�MvC�3ao�p��g�B5[�dE��I��t����M�b�s��x�8���<J�)�ϭW冎�s��}�6TrY��(��X��2A�c��>��ś\����������;U7�TY��w������ω����:���\sNm���Ny;�Q���]��NO�x`�͙�|2���{��S-2AV������ژ�8��5P(G���ļ�8�#ig�\�u�u4�]��L��U��}\"��!�YEe����e�S��.�{�~�i�s�=�oL�Xܨ:�db��}r�$�����9��[%mm��oj���X^�Kx��&K�@U�˟����ˇ�Q�F�ŐLL�6�voo�w��\t��]H$�p�o��l;*�Q-2�y�����!tn;ކh*���^D��`D��&l/�&���y�����gE�҇B������_���g�9��f/�u�{�&���K� ��@u_��*��WKa|Z݈f�H[-c-��5je�n9�G7|
�e/2}��~!b�`�n��Q���g�P���P�-�x˟(��}��^�c��)	w�����#O����z�!�Y�]�d�s���+hy���B&^c��[Dy��J(�4���
�!h��7ލ��S�	�x$y3"h���k��?��~��+W
�հ�FR����~!�,�������$�?Կ{P�~D�b���Aط��S,�7SӸ|�OF�>Y�bn�*�En���ӱY���bW'J�Q�ނO��r�N_,�'������t��մ3�'v�ii�����]ö�j��&=�E���"��w�]X�Q��|�'5[�A��=rO�vk�V��답v�VǪ߅e�j^�O����/��_{$e���O��_����%ϊnJ���]���MCd�������Eq����H�H&�"�N�]��Y�}>��]mk"���Ɛ��gD|a����FV�EK��c,Ȋi�u��#P��7�-���eU��(�2�r�g�G��O���x��I)#���h� K�I��s�W������[�'�{�$��$�c��/��A��σv;�gWZ�Jih*���S���`f�6Vi���^�K����<f�,��	w��Vu����θa��EQ&��P�u��XS��v�N�R��JB�W"˼��JQl��ex���^��S'�*�����T�W\����'տSl���q�G�}׸��y���g����M���dq��*�$��2�t9,VޑH�hEE�R���`�z]+J{Lی_���P���5�ݤ4=P�\���n�+\��O3������J��ɦq0cL���YB"P�P<��߂?=�Ѣ���c�I�TG��(��˦�;f���k^�4�/e�nH7z��4�m�������O.���l���d���������������Z7q��><%�bV͢�����ё_a�5�I�1��x@n�����c���;�z��:Z9����N>?�����DQ-�����R�Z�Pa�:[������Z�C(��Z�>k��)	�Kw�=J��^�%Mx�n��$��uBKF�$6u�]4k;6OLL��4���UlW���8��EQё�ʘ��,wDT������j�D@ˇt$��
#�
�xn��Fm#NTgY�\�eIι���Wgy�8zJ��R��|���3�&��ɶ#�����?�~�i���G�i;��0F�e�oH���m��us��[;4ofpud�8�r��8)>��D��b�J���G�hJ<��|��P85o��$���sl�N+~œ�,Jv�ه��*.- �î���7ԑ3e�ƍ��O��^*�6���/�y��9�E��-�rw^a�����xW6��X������^ޯ�@z�م��U��m�lt����z;Y������H�ګD~	K?��ڭ&I0.͇�T Ϸ��&��V���9<�����/e��I������IғvͲο��p�����/����"K�]����t�b�BW�m���.��mQ%߾vɽ��9Wx�(�k���n��ó��x.�&��3�L���-������y�<=������ �1İV]��Z���gM;�j�*���ۥҍi�W��%?�iQ`TŖE�ة�G��?��Ϯot|sEGw��s-K�o�L<��W��2HeBP��m�B�bƇ�[��`�{��U|���
Ϙ��JI�*�A���.�����͛�q�IN/���k�X�x�|��	    IEND�B`�PK
     �)K["1^FHo Ho /   images/6b6fcb51-98f7-4a52-b90f-3140c0078893.png�PNG

   IHDR  �  �   �r��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ��IDATx���1mA  ���+w!`0�t ^z )�-(R^$E�}i��_]���s� ����\k�       ����|��5 ����cp{��朏��s p'         �%�          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��     ���<F��~��k�fq�\��PVeqU������T��T��aIl���6�4���%��5�j)mm<j�j����J�"" �s>�V��@X�3�x$��?;3���_�y}     � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	���7�o�=���������r�l��ʲ����1(5���z��7       �Z�vm�1�@����}����c�3?�7�۲7�S���?p��͹.x�%K�
���q�GF]]]6={��#�8"�u����o����///�~>�y�>/         ��k��o��F�ڵ+���Ν;���cǎؾ}{6���Jl۶-{=I�~s
^E UEEE444dӫW�l���ߺ���UUU         t���ټ�bڏbϞ=Y�e˖x�嗳s�l޼9���g�>�;�\.�썍�q��G�QG}����޽{g�         ţ�����z�󝝝�u��,tߴi�[�q���}���������������c�9歨�v         `��r�^�ze3x��w<�w��x���^Ȃ��lذ!����ަ��>�?��8�㲨=���#          TEEE{�ټݫ���ׯ�b��������6x(UwJVuuu������          ]�{����ܜ�~�v��>�~��l�}��رcG@��S2�8�,b�O���������          HEMMM455e3al���/�O>�d<��Sٹm۶�b%p�h����'?��2dH�766F.�         �B�o�d~�<���M�6e��ڵkc͚5��+��;E#�����YО�UG>j///         �bҧO�lƌ���y��,t_�jUv�ٳ'�P	�)huuu1t��lN<���          ����!��ڲ��������}��ձe˖�B"p�����/ZZZ���'>��z         ����ʷ��mذ!���X�n]tvv�L�NAhll��O?=N;��         �ֿ�l&M��ms��b�ʕ��3ψ�I���d����)���E�MMM         ���իW�;6��_~9�ꞏݟ~��T�IJ�޽���5���\.          8�����7o�U�V�_��X�~}��$p��ѣG�1"�          �NCC�[����?+V��Gy$��]M��a���>dȐhkk�SN9%���         �ë_�~�L�:5֮]˖-��<�����t�#�<2F�g�qF�m          ғ_f��ܜ���۳����}�ƍ����C����[[[���,          (=z�c�f�nݺ,t�Gb������C�gϞ1r��8��3���>          (l�|6ӧO��+WƟ���x���;�	'��ƍ�aÆe��         (.�����֖�ڵk��{�������q�9(�!�СC��sύ���          �42$�M�6e�z�سgO����TWWǈ#���}��          JS�>}b�̙1q��x���O�S������RWW���q�YgE���          ���)S����_��{^z)�����Y�����ڢ��2          �TWWg��?��X�zu�}�������;Jccc�{�1r����r          F�=mii��g����+�zꩀ�"p�}����ĉc̘1QVV          p�����_�B�Y�&�׭[�vw�S�޽cҤI�v          ����2dH�^�:~���Ɔ��C�^�b���q�gDE��          �F.�����:th��o�%K��K/��63����7n\�;6*++          �B>t?����SO�B����7�iӦ�4	�K\MMML�81۫��          �����a�b���t��رcGPZ�%*�`�ȑ1cƌ�ѣG          @
***���=F������{��A�^�\pA80           E���1}��3fL��W��U�V�O�^Bz��ӦM�6��7�         @����W_}u�Y�&n���ظqcP��%���2Ǝ�'O����          �B����_}<����t��عsgP|�E���%f͚���          ����<[�<r�����<�@�۷/(�"�����͋N8!          ��t��=fΜ�G������nݺ�8܋L�[)�sNL�:5**��          �����c���q�w�믿6t���^x��	          � ��E[[[477��ŋ�'�
���TUUŔ)SbܸqQVV          Pj��k���+W�/~�رcGPx�N��s�F}}}          @�;��bРA��_�:~�ᠰ�TmmmL�>=��          �_=z�/�8N?��X�xqlٲ%(�4|�������.          ��6t����W�w�yg,[�,:;;��	�HMMM̞=;F�          ��֭[̝;7Z[[cѢE�m۶ ]�1p��X�`Au�Q          |4'�xb|�+_�[o�5V�Z�I�������<yrL�4)�          L]]]\u�U�|�����c���AZ�	�������hjj
          ����r���'�pB��'?�6��'jԨQ1{�쨩�	          ��jll�뮻.�.]��sOtvv���=1ݺu�9s�Ĉ#          8t*++c�������-��[����=!������իW           ]#�_���ӟ�4�x����'���-f͚�          �juuuq�5��=��w�uWtvv]OM}��ok0gΜ�ԧ>          ����b	�����rK�ܹ3�Z�èw��q�W���          @ZZZb�q��7�ƍ��#p?LN>��������           �ҧO�����zk�X�"��.��m����cڴi�5          �������KcȐ!��_�2�x����w�����袋���5          �����G}t���?��۷��������/����V          @a4hP,\�0~��ĺu�CC��������/�nݺ          P�z��_��cѢE�bŊ���bcƌ��s�Fyyy           ����2.��hll��K������r1eʔl          �Ɀ����;�#����C���".���1bD           �i�رQ__?��c�����'p?Ⱥw�W^ye4(          ��6lذ���?7�tSl߾=�x�QCCC\s�5ѷo�           JÀ�뮋�}�{��/N�~�80��ꪨ��          ���e�K_��o�9�|���������������           JSmmm\{�hѢx��G��N��1><,Xeee          �����lyvuuu,_�<�h�C[[[̝;7r�\           ����y��EMMM�w�}��'p?@���1k�,q;          �.�������"����w��#p? &L��ӧ          ��9�󢪪*�����	�?��lʔ)          �a�lWWW�m�������&p����"���          �����=���c���"��!p����b޼y1f̘           8mmmQSS��rK�����	�?@>n����O?=           >��ÇGEEE��G?�������r��vq;          p�����%�\�E�����K��?���ٳgǘ1c          �`:��Sc�����,:;;��#p��M�g�yf           
�G��]�v�m�����{�:ujL�0!           ���:+^{�X�dI p���>;&O�           ]aҤI�{����	�ߦ��=fΜ           ]鳟�l�ݻ7���(e��o���1k֬           8f̘�v�e˖E������5�ϟ�\.           �|�<w��,r��G��|�����^zi���          �ᔏ�/���رcG�Y�&JMI�q�e�Eyyy           � �7_q��o|#�{�(%%�y���}.jkk           %555Y����=�l���$�����ꪫ���>           RԳgϬ{��7����z��������K.�          @ʎ;��⦛n�}��E�+��}�̙1lذ           ('�|r̞=;/^Ů������Yg�           ��3Έ_|1���(f%����Ĵi�          �������'{�(V%�80.��(++          �B���b���o}+���E1*���G�q��Geee           ���������o��[�F�)�����<��޳g�           (�%��N����v�ݻ7�IQ�3gΌA�          @1ijj�iӦ�w�Ťh��#GF{{{           �s�9'6l�?�p��܏=�ؘ7o^           �9s�����c�ƍQ�.p����+��2���          ��UWWg��׾��عsg��
�s�\tttDCCC           ��>}���_�������3
YQ���g��O          �R���'N�?��QȊ&p6lX�{�          P��N��ׯ�����Q��"p����V��r�           (E��z��q�7�֭[�|��.���֭[           ���ݻg}�w�����BS����ɓc���          @Dsss�}��q�}�E�)��}��1iҤ           ࿦M����?cÆQH
6p�������(//           ����"�o���سgO���gϞ}��	           ޭ��1f̘��v[���O=��=zt           𿵷��O<�V��BPp�{�^�b޼y          ����r1����b��푺�
��܋.�(�w�           |��������w�������
�'L�C�	           >��N:)������L�޷oߘ2eJ           ��M�>=V�^�7o�TD����b���QYY     ��ػ�(��;��)00�.��4�R#�A��c�&z�9ɉ���$'�����I�;!ш�b7�=XŀH�D�I�����DQʔ;3��9Ϲ�/1̝�e���     _ݺu��+��o�1�����Z�i~׮]          �#WRR���_=rQ��M�6���??           8z�]vY̙3'6o��&��+��"�ׯ           ��%�\����"��t��F����7           (?C����z+f͚�$g��+��K/           ���_|�A���F����=��5
           �_������Ϗ|0rEN�%%%��{           *�i��3f̈�F.ȹ����(������           *N궿�������سgOU�qr/p?묳�E�          @�;��c��SO��S�V�%��f͚�g�           T�s�=7�x�زeK��9r*p��⋣nݺ          @�)..�"��￿J�9�w��%           T�#F�K/�+W���?CN�yyyq�e�e�           T�������K㷿�m��r"p6lXt��1           �:%%%ѷo�x��w����<p�W�^�w�y          @ջ�Kb��ٱ{��J��*�ǌM�4	           �^�V���N�g�}���J�}��          �i�����cӦM�z�U������U>D          �O�W�^�w�yq��V��VY]ޥK��۷o           �{��?�|�^��������??           �M���1f̘7n\��g��%%%q�	'           �k������OǊ+*���$p?�s          �ܖ�����w�qG��_��{��nݺ           ��_�~ѩS�X�dI��W����}           ��ԁ�3&n��
��J����           T}��Ν;ǢE�*�~*-p7�          ��:��s㦛n������}���Ѿ}�           ��9���{��1o޼
��J	����Mo          ���?������+��WJ�>x��8�c          ��k׮q�	'�|P!_�R�Q�F           ���ѣ�o�޳g�h߾}           P����+k�W�XQ�_��w��          j��O?=&L�P�_�B�T嗔�           5�����G��?��\�n��G�����           ��(,,��#Gf�{�~ݨ M�6�           5ϩ��O=�T�����׬�����OϪ|           j����6lXL�:�ܾf����ՋSN9%           ���8�x�����\�^��#F�����           5W�-���1cƌr�z���ȑ#          ��o��ѹ����y��          @�שS��ܹs,Z�訿V�rJ           P{��<���-[�	'�           ����z(�m�vT_�\�#FD^^^           P{ԩS'/���Q}�r����c�С          @�3|���	����M�4	           j��;F�bٲeG�5�-p?�S          ��+Mq�ӟ�tğ_.�{��ͣ��$           ���&M����#��r	�������           ���_�~0 ^{�#����S�~��'           >���޽{GӦM           �t��ڵ�U�V��u�>lذ           �}N>��x����*p/..��={           �3p���4iR�ݻ��>��~��Ea�Q�          �i֬Yt��9.\xX�wTuz��          ���޼���FIII           �?K��C=eee��9G����?


           �Y�ƍ�k׮1o޼C��#�SM           3`����5jݻw           8��?��QVVvHD�{�����           ���7\}�ܹ���G�80           �������&M�D׮]           �H�������={�|��v�>`�����           �"6�����={�~�a����           8T�{�.���~��ѵk�           �C���'~��V�ޫW�(((           8T-[��֭[ǚ5k>��+pO�<           ��={�_�����Mp���m۶^߾}{�ݻ�S�N)**��z�YV�^�          *_�ѧM���sȁ{�Ν�A� Gc׮]�iӦ���c��ͱe˖غuk��p}�J����Ǝ;b��ݱs����={����N�:�J�{��������ׯ���o�{�q��ѨQ������u 
         �w��{�%<�C.�N<�� �ϓ��6dk�����/jO�zUK?���I��*E�M�4ɂ�f͚E��ͳ۴Z�h�ݦ8         �?u�֍nݺŜ9s�1w K��?����裏b͚5ܦi���)�W�>��4l�0Z�j�[�>���c��y         ��z��u�{
�:v� �7n��U�Vp{�S�k�-[�dk��şz_��޶m�l�k�n�m�         j��={~��)p/))���� �fJ1��e�b�ҥ��%KbӦMA�HS�Ӛ;w�oO�{�P֡C���{Zyyy       �^�v������ۣ��4{yϞ=��;w�ݻwǎ;����y��ԩ��}�ի�@�����������կ_?�ur= G�c���-[�ڵk?�������# �RX�����hѢ,hO7T���ͬY���O�F��S�Nq����_�       �����6d���͛��~��[�f�z��sɾ�=ui5l�0�6m��6n�8{9�k޼yR�@-�����⋟�>�;@VVV+V�����g1{Z�ׯ��t���{�e+I�����w��%�u�mڴ	        ���}͚5��裏�f#��7fa{��^]�&�ɻ����f͚e�{�-�պu�hժU�� ��Q��J�!@�KA����c���p�;wn����c�޽�z��l���k��҅`��޵k�())�:d!<       P�R�����=[+W��?�0��S�^ZZ�#�Ok�ҥ�z_�Ҕ��(��]�vѶm�l�	� �\�wK?R�Ͼ0p�޽{ ��V�Z��~̙3'�����I��f��V���J�{:���O�vA       G'M+_�lY6|0�i������5�[�.[i��'g�{��۷o��;��c���( ��4h�=Ƨb�L�P�lٲ%fϞ�E�i�c���6o�o��f��6m�d�{Z)|�[�n        �-E�i��%K��im۶-�<����O~~~�Aw�q�J'�w��Q�PMu��M�P]�ݾ��n���{1o޼سgO��Jǟ�5mڴ�S�Nv�K�޽����1_       P��ر#V�X���,�ŋg���=iZ��ի���odo����=MyO]D���� r[
�_x�O��s�F�E�֭�ʕ����}�̙YԞ�a��k׮���|����}�{��      ��n�ƍ1���+��ij;��'���ӧgo+..�B�N������[� ��!�n����b�����E�bƌ��[oŦM�*Zځ��SO=�Ms�ׯ_0 �t��9        5Bj0� �>� �׬Y�l۶m�Y�fe+)**�Z��D���C��#7n�Z������܏?�� ���޽;fϞ�E��	���������c�ԩ�jڴi�4H�      @��N7_�`A�ϝ;7�-[fB{-WZZs���֣�>��;w�b�����T��x|X�{� �W�`Z�pa���曱y��\��c{��լY��߿6�=�       �&�qi��{ｗ��i� L
������-[F�^��O�>ѽ{��S�N P9�@��ӧ��ѡC� �|�Z�*��׿fQ������u�d�c�=6C���w       �
eee�|���Q�ҥK��ڵk�Lq{ ػw�l`ӦM���Y���o�>�֭ ��۷�[o����ij;Tw+W��?�����#�dGt:4N:�$�       �p�v�9s��̙3��wߍm۶����l�t��z(�,�N�O}D��@�J�zQQQv��>�Ӄ2 �o�޽���^{-�y��I/�4������dS�O>���رc       @y�Ϙ1#�0v��PYR�hѢlM�4)ڶm�Mu8p`�2 G/???:t���������5�Óv�I�S�N͎-��"���wLWz�p�)�d�{�U       ����,>����>}z6���]�*�^�:��l�݇�Z�
 �\�N�-pO%< _l�ҥ���/gU��Sۥ~��4hP�92�=��       �ϓ&e/\�0����o��͛r�'c�4pȐ!Y+Ѹq� ��w�q����{aa��3 >G
�S�>mڴX�re JG¥�iu��=N;��۷ov�       �f͚��_���6TG�N�4)z��'�|r���'


�/�σ�?3po߾�V�ϰiӦx���^�-[����͛���-[ƈ#b���ѠA�       �vJ�g͚�M�;wn6�j�={�d��*..�ĩ������ �M�6Q�n�عsg��g�L�dɒ��_�o��v�D8|k׮�ɓ'ǓO>��TNS�[�j       ���H�g̘���5ٶm۲Miu��18dȐ(**
 ����{l,^�8{�3��P[-X� �y�lW%P>v��S�N�iӦE�޽c̘1ѩS�       ���7���矏��FK�.�֤I�bРA��|������{*�j�t��{�O<�D�s��{m߱\]�t���:+���       T�W�Φ�O�>=�o��?���Z��0 
��k߾���?�Q�m۶P��޽;^{�lb�ڵk�<i��m�ݖMr��W�}������       ��H���Ν��Ꝇ�ׁϖZ��z�8����N��M�@m��~�S�{z�,..��"��o��VL�2E�U,��0v��h׮]�y�1d��;      @�+--�7�x#���lr;p�6oޜ�L�?i �Q������&5c�~�;j������'�x"6l�@�X�jU�?>��K�����#???       ��q���˱m۶ �\j�f̘���ݻg�DϞ=j��F�F���?w��ٳgO���Yؾq�� r׾���瞋��;/۩      @�Z�v���}׮]��y��e��c��ѣG��c���>��m�6 j��{���o��<�H�Y�&��cŊq��gGp]p�QRR       T����4��7ވ��� *�ʕ+����=�X�~��q�)�Dݺu��J�g�mڴ	�����ߏI�&������/^���o�G�q�Fǎ      ���hѢxꩧ�����kݺu���f߇��zj�5*�ի 5�1���
܁-Ű?�p,X� ��#mZ�;wn0 �[�l       ��}a��Y��z�7o��<^x���,tj�V�Ze��EEEѨQ� ��6l�O<�D���+vC����z뭘9sf�;��sύ���       ��,\�0�L��rϖ-[����_�"������kݺuv[��o����ꪴ�4�}��x�gb׮]�|{�쉩S��믿g�yf�~��QXX       �U�Ve��3�}i���ɓ�^j���q�i�E�:u��jٲe������PݤI�/��r<��c�7��ٺukv��ꫯƥ�^�z�
       �غu�⩧��~�ZVV@��&��f�^���>;��� �Mz�j޼��'�T7K�.��'ƢE���?�[n�%����]vY��      �O۸qc<��Y؞N������ǽ��S�N�.� ��� �M���`@u��5�c��M��Mp��Y�fŜ9sbĈ�E[QQQ       �s�ά�x��'cǎ�,�V���o�=:w�_|qt��% ��Գ���� �.��.��L�۷o��ٽ{w�+��wމK/�4���       �U ���oǤI�bݺu�l�-�믿>N:餸袋A��Գ܁je����1:K�,	�C����;�O�>�}-Z�h       ��ܹs㡇�+VP{��-3f̈Y�f�g�g�uVԫW/ rէ�f͚@.JGc=�����s�e��D�XK�h3z��8�쳣��        j�6�#�<ӧO��ڵkW<��S��k�e�܇yyy�kRϾ?p/..�+�I��NL�81��8Z�6̼���o|#:u�       5��ݻ��_�G}4JKK ���c���1mڴ����u@�9`�{ӦM �l޼9~�a;��
�|����/Ç�K.�$���      �&H�[?���v�� �,K�,ɺ�4���/�F�@.HM���=�s�3f̈��?��*�޽{��_��s��UW]ݻw      ��j�ƍ1q�Ę9sf |��M��iS�E]�	�����TXX��{�&M��mڴ)��~�� �,}�Q�����i�      @�TVVӦM�G}4JKK�pl۶-���x�����_�z�m�6 ������@UKS���غuk T�}��?�����ꫣs��      ��-[���K�.��1����Og�qF�{�Q�N� �
��ƍ@UرcG<���YX
P�֬Y�_}�5*�?��(((      �\�&�����^x!�P����<�L���;q�UWE׮]��	܁*�dɒ��{�� W�����ڼy��k��֭[      @�HS����?�-�
���o~�>|x\r�%QTT �E�T��>��s�裏f�� r��ŋ��?�y\|��q�)�      @UڱcG�ZL�6��v�¥Ǚ�_~9�̙�Ms/))	�ʰ?poذa T�u�������� �.�ѽ����~|�߈���       �l�g��~w�~�� �L�������iH�i�@E��7h�  *ڌ3���m۶@u���D�k��&�u�       �a׮]1eʔx��gMm�Lz�y饗��6��ַ�K�.PQ�)M@����c���P]�I7�pC�92��կFaaa       T�իWǸq�bŊ��4����7q��gǘ1c"??? �[Ve�׭[7 *¢E��������K;��N��=�}�;߉-Z      @yJ��|�W����;w@.)++��<�̙�\sM�j�* �S�7k֬(/// ���/�'N�ݻw@M�dɒ�����ճg�       (�7o�	&�{� �,���~�_~y:4 �K�7mڴ^ ��]�v�������j �T[�n�[n�%F�^xa�0      �ٳg����شiS T;v����ǬY����F�����@9ٰaC�q��tc��.��3���ի�ꫯv�      �4Hp���1mڴ�w� �͌3b���q�5�D�n��hd�{qqq� (��͋��+;.�6I;�����;����h׮]       ��+W�=�ܓ�Tg�ׯ�n�!F�_��W���0 �D��QTT$p�J�=����#�<eeeP�Y�&~��_�UW]      �����/�ĉc���P��l�ԩ�lٲ��w�M�4	��%p�ڎ;b	���o@mWZZw�}w̝;7.���(((      �OڵkW����+P-X� ~�ӟƷ���8��p�ܝ�?�0Ǝ�W�j����hذa�۲iӦ�z��W�ݘP��I��߳�ȍ7      �dÆq�wĒ%K�&ۼys�x�q�ęg� �*��֭k�;p�f͚�ƍ˦S}իW/5j4H�X���!�ԩ��~�����y��׏���O}Ϳ��o�q�ƀ�n����_�"��_�5�;�       j�y���]wݕE� �AYYYL�<9V�XW^ye�|�;pD�d�?��O�rS~~�����mڴ��m�F˖-�U�VѢE�,lO�zyK�!p�H�������k�_�~      �>��g�}6y��P+����jժ��w���K �'��������<[��w��%N<���ڵk���ѡC��رc6q����}���C:�"18f̘8��s      �=v��&L���~; j�4��g?�Y\}�Ն�k_�� _`׮]����>�z� w����N�=zD�n�8�gԨQU�gJ�;p�}��D�+��"
      ��>���;vl�^�:�Q�F�Ջ�?�8��J�~Ґ�ѣGǅ^yy�U�Ӳ�����#�6o���v[,^�8�z��q�}���^�zEQQQ��;\:Yaݺuّ[���      �fJ�� �t�35Gf��֫Wo�˩�(((�n�`�t[\\4�VӦM�y����������?P��!��<�L���k��O ���yyy�pk֬�[n�%��j�m�v�ްa��Uw�|s�΍_���q�u�E�f�      �Y���x衇����!��-Z��V��4i���"���p=M`?�
�?�f͊_���o��oѦM� �'�����	��gZ�pa�~��e˖�j���={������:Hxig�����l�V��_����}/ڷo      @�WVV'N�_|1�=�e8��G�1��شiSt��)[�s�Q��"�yyy6?�������W���~��ѽ{� HLpꭷ�ʎ�ڵkWP�:v�'�tR�x��qV�M�q�|�� n�ƍq�7ĵ�^�"      ����Ҹ�����rG�WRR�E�)d/((�ޞB����4>�����[��M7�W^ye:4 ���IO=�T<��v�V�t�U��~��'W�cw�ph�m�7�|s|�[ߊ���      P�lذ!n���X�bEP�RD������7�t�?j�i����{��l�~�w��j�� �'S�L��<�<͚5�dۋ���&H�;ph�Iw�uW\u�U�/})      ��c�ʕq�-�d�;U'???�v��{��&���=W��b�(c}��'cݺuYC������~`��ᡇ��>��۷�aÆeV5mס�OYYYL�0!v��#G�       �͙3'�����|T�&M�dQ��A����M|��_=>�����w��������V�{��ꫯ+���|:4;��r1�/m4z���c�F�      @�z�W���˚*W��|�	'Ā���lѢE �o�ܹ��_�:���h֬Y ����?5x���A�IGa��ib{�֭��KO,

bϞ=��?��ñy��袋      �-�wz�'O�g�}6�\�5ʢ���GqqqTW�¡Y�jU\��Y�~�1�P{ܡ�KS�Ǎ3g�*F�%|�'�i��V�vঠ�y����Gp��y����/�v�      ��JC���?�k��T�v��Ő!C����G��7nEEEQZZ��[�n]��W�����N�:P;ܡ۹sg�;6�̙��4��W�^1bĈ��GK��w8r)r߾}{\q�"w      �bi���~���1cFP�Rw���/}�KѦM��iRK��S_l۶mq�7������ҥK 5��j�����o��s��+E��k�ȑѬY���Z�j��~ G^�����oֈI      P�����w�y'�Xi�y������I�&QS���w8ti@�M7��^{m���#��M��P��v�-�ĢE���չs�5jT�m�6�Z;���믿;v��|�;QX��      T�4�j�ر�U���СCc���Q�^���R���x|뭷Ʒ����ׯ_ 5�B
j�H��Z�.]������g��:u
�O����w�}7ƍ�E�&�     @�H�����A�ٴ�!C�D�:u��04�L:Q㮻�o}�[1`�� j&�;�";w��v����O�ƍ���O�>}�D^^^p�t1����ݻ7��7s�̘0aB|����      l۶mq�M7Œ%K��W[��}Lp�#�gϞlH`�:lذ j�;�i��w�����^��JX#F���u�����(5j�6m
�|L�>=


��+��     @I����c�ʕA�*..�SN9%���7_KC���eee�����?�1��ӀR�f����I;���Θ={vptRLڻw�8�3���|���X����W_�z��ť�^      @�Z�~}�����5k��'<xp><�}gm���&M�Ć82{��|0�o��sN 5��j��Sm���1k֬�褝�g�}vt��%8t)p_�hQ �����&�@     ��v�ڸ��ȝ�N�0`@�1"6l���T���M�2%��P@�!p�,�P�����7��\�:ubذa���|4֑Jc@�Hh�1��3�      ��lܸ1��.n/?�;w���:+Z�n|Zj*�ϟ��KEj��cP�)5�{���W^	�\III|�+_Ɏ���ܡb���Ύ�;��S      82�7o�o�1����K�@�խ[���Z�h@�IE���8� �7�;�P�'O����/��iРA�=:����;T�tZ���ߟ]���&      �óm۶���c����ѩ_�~�92������T@�KCaӠ��ÇP}	ܡz����g�	�LϞ=����"w�^�F����(JKK�)r���{���E      ��ٱcG�t�M�lٲ�����E�>}�a�z�C'p�����/k(@�$p��W^�)S���q��q�9�D��݃�.b��ʕ+�8eee���.6l%%%      |�]�v�m��K�,	�\�6mb̘1ѡC�����I�i�P~RC1~��,rO�o��G�5��ٳ��g�4�=]l�O��cϞ=q�wď~��h׮]       �m�������͛��u��ȑ#cȐ!�����T�X�"���;�3��_�%kÀ�E�5ĪU�����v�q��.�Q�Fŀ��ӢE� *���۳)?�񏳓)      ��;�o�[pd:v��w�����w��63]w�uѭ[� ��;� 7n��o�9�9t�;w�.�@ Z	�nc��]�6n�����~��      ��޽{c���1cƌ���$x�I'E^^^p�4P�v�ܙ5������9@� p�jnǎ��6�&�5bĈ8��S]lUcP��.]�ƍ�k���q�      ���w�}��o����$ƌ�5
ʏ�*^j�� ����Ѷm� r����td�=��˗/M�&M��/��;.�<�8�ئ��@�5kVL�<9{�     ����'���_~98<���ѣGǀ��'p�ʱe˖��[�'?�I4n�8��&p�j���EM�=��΋������� �5k�֭�r=��s�&��#G      �Vo��V<��c��I/���h޼yP1�[C�r�v��[o����� w	ܡ�z���^�X���:�4hPPuҎc�;T�|0�G��}�      �6��Ϗ����޽{�CSXX_��cذa���T�Ե4m�4֯_@�[�ti�7.����ls	���P͘1#y�����d.��lG1U+�|�A �/��Ogir�N�      j��>�(���ؽ{wphZ�j_|q�i�&����C�5kVL�4)�ʀ�$p�jf���v��;fOB6lT�t1T��;w�رc�?��?���      P�mݺ5n���ؼysphҩ�cƌ��u��'5�������/ɾ�F�@��C5�.�Ү�]�v���:�����Ow�L�C�۸qc�v�m��(�ԩ      PS��"�nl͚5�KA�9�}��	*���ƃ>͛7�6� �E��DYYY�u�]�aÆ��
��s���#�#̀��lٲ���{�ꫯ      �������b��kӦM\z�ѢE��jܡj�&oܸq���?�?�� r����I�&9��4j�(.��h߾}�{�ի6�-[�P��O��:ur�      5��ɓ�7��X�޽�A�i�;U���:;wc�Ə�cߋ�C�P̜93������9昸��ˣI�&A�J;���1[�ڵ�N8!      ��x饗��g�>_~~~�v�i1|���5h� ���c۶mT��?�8n����я~�����	�!ǭZ�*Ə���g�ѣG\t�EQ�N� ���}ɒ%T�t���w���_�͚5      ��.\'N>_�F��K.�:�#M��C�I��]w������M@@��C۱cG�C���4�lC��3�<3������-�7o�;�3~��Fa���      T_i�n��מ={��k۶m|�k_�&M��%\�|y UgΜ9��c��\@�R2A�J������ի�OKA�駟j�U�V�ŋ��ɓ��K/      ��RԞ�ȝ��ٳgm֩S'�=�Bnx�駣}��1p�� ���r�SO=3g�>-MN\�z�
�����=�?�|t��%      P�L�81,X|�4Dpذa� ��2�IS�a�`�֭[G��w�A��~L�2%��z���W\��C5��8K;�w��@n�0aB�k�.;�      ���^{-^z�೥��_t�EѣG� �	�!w����;������P��c6n�w�}w���JO����8�c��)�OGj��� ����Ƹq��'?��#	     �V�X���ي���k_��!��D�f͢�� ���@�[�vm��]w�u���@��CIǛ�?>�n�(M��ꪫ�8��-�8�CnJ� 8iҤ��       ���b�ر�s���Ӛ7o_���u�H��S䞢Z 7�������O��g�@��Cy��b�ܹ��R�&��ȝ�ϑZ�ۦM�%%%ѯ_�      �\��s�=B��h߾}\~��ѠA��zIM��א[{��ԩS�x�T�;��˗ǣ�>�M�6��v]5��r߄	�c
�T      �5���={��c�>��:�Ï_��Җ����e�K�jX�l��j�؊�=��˼�8�E�v��$��E�U�UHt$$!�*zG4�����h�([���g�_$v{�9�>�뺃ˍ3&����:����򣩀ғ��~��_����0`@ �C�%���1~��_GSSS�aÆeq{�޽��p��w����p����,*++      J����c�����&L��=�XTUU婶�6��s�ԩ�������Gt�;����~:���|j������XܞC)pO/z---��>� ���C=      P
N�8��F���r�3fd��UTT���@(][�n�^x!}�� :���؆��^>5bĈ,n�իW�?ݺu��������(m�`���}-F�      ЕR���_�:Μ9\쮻�o~�A��Ci�7o^|��_�q��б�Ѕ��%&�/6l�0q{���J_�i!����?�yTWW      t����\�[��V�y�A>�^���� ������W��_��ѯ_� :���H��Kq�ɓ'��?��O����>� ��w���x����'�      �
�w��>�TEEE���1{�� _RS!p�ҕz�������}�w1�1��E/^��np^mmm���w��A��R�˒%K���.Ə      ЙΝ;���MMM�y)�|��b֬YA���f׮]��6d��}��@��Cؿ̝;78o��Y�ާO���P^ҭ#����㗿��A$      :��O?��:�y)n��c�̙A>i*�<<��s1f̘���hw�d)���~���AD߾}�?�i�ScP~�?�<�L��'?	      �iC�e˂�R�������Ӄ��T@yH7����g���kTWWо���,X۶m"z��?�яb���A����d[�Ϟ=@�X�bEL�6-���      :ҩS��7��M�H����o�����6��o߾x������}	ܡ<x0^x� �����1lذ��ҁL����C��̆�      �#��=��'O�λ����;��/-��֭[�(}/��r�(�_�j �G��$�~���Fccc]eee<���/})(�t���ݻ(/G���s�fCJ      �/^��npޜ9s����!u5)r?|�p ��m(����e�Ў��I��k�֭A��?�ƍ�m�����W_}5�M�f�     �vw���l��͚5+��ޠX��@�;��#G�ĳ�>?�яhw�Ǐ�?���A�]wݕE�P[[@yJ�ǿ��������      �������o���A������'�@yY�lYL�:��Wh'w�O=�T444D�}�k_���/ q��6g������|'      �=���+�u�� bԨQ��c�EEEEP<�B�ICZ��������ߢG���;t���z+֯_E7bĈx���������[�n���@y�7o^L�>=�      p#�9�?�|p����~�}�N1Y���ѣ��?�9����pc�A����?��Qt���GQ]]Ц��2�
�<��?�����       �-m���o~Qt�{��Xt��=(.�;��ŋǔ)S��n��	ܡ����ǏG��W�*���	�T:�	ܡ�mٲ%֬Y�g�      �˖-˾w*�^�z��C�ѳg��ӧO�>}:�򒆶~����/~�7q��:Ⱦ}�bɒ%Qdi�>C��ǐ�<�LL�81z��      p-N�<s�΍���������G��gA�����1����w����CHSXO=�T���D�}��_�������`�p�ԩx���_�     ���ӟ�gϞ�"Ky�5jT@��T�ܹ3��4o޼�>}z6,�k'p��v���_�5v��,p��#p��H���q�q��7      \��7�믿E7gΜ�4iR��4Pޚ����C��g?���k#p�vV__�=�\Ymmm<���>��B�0�~Nҭ@yK����K������      |��������7n\�s�=�J�P�Ғ�5k���ٳ�6whg/��R�8q"��{����OF�=�H�y�۷o�<y2��u��X�n]v�      |��W>|8�lذa�lp�|x�gb	QSS���C;:x�`,^�8����!C�\����!G��l�ĉ�       \ɡC�b�Qd�{���^��2`���֭[455P�N�:�?�|��?��	ܡ=�쳅~��1cFL�4)�Z���m۶�Ǐ�~��      �J���?�������}�{1p���ϒ6����f7����k��]w���rK WG��d˖-�~��(�#F����p�\�����/g����      \(�6l�"�ַ��F�
�"���C�kii���z*����9^����Akkk<��3QT麬'�x"�	�U�6򥡡!�^��?�q      @�����}ERWW�g���
ȏm۶�ڵkc֬Y|15*�����k׮(��~�n���ȧ+V�׿�����[      �ġC���R���#�\-M�˳�>�&M��={���p�������dq�Ѕ�կ_�쥭��>��H��<��s���      'N�����GQu��=�|���ѣG���C�|��G�g�c�=����Z�dI;v,�hРA&�iiJ}�޽��{ｗ=�ƍ      ����s444DQ}�;߉!C�\��STTTdƀ|X�hQ�}��ٟo�	��|��ǅ�.����'�x�d1�"M�!��Νcǎ�~�     @1�ٳ'V�^E5y��8qb��J]N߾}��ɓ�Cccc6�����|6�;܀ę3g�����7��\���k׮x��cʔ)     @1=��3���E4hРx���W��,p�|Y�vm�{�1r�� �L���ԩS�x��(��Çǜ9sڋ��-mq�4iRv�      �����{�ETUUO<�D���Wj*v��@~���������������rw�N/��R���G�t��-{���E��v������;�#      (�����瞋���7�7�|s���T@>m߾=֯_�'O�rw�ǎ�e˖E}�߈�C���t%[�hnn �^|�Ř9sf6(     @1�%H���"���g��Qwȯ46q�Ĩ���b
#���͋���(��n�)n���������Ƒ#Gȧ�G�ƪU����      �/u/��RQϞ=�G�����U[[@><x0֬Y�Ƀ+��5:~�x�\�2�&ȏ>��i1:L�8�C���/�e��     ��k��V��z��߿@{H?K������@����1c�-\�F���/���9s�Đ!C:�+� ��;�]Cy�]w      ������͋";vlL�81���� ���?G��e˖�7�� >%p�k��GŊ+�h�*F�ùR�!mq�={��c     �{�W��ɓQ4}��Gy$�����wȯ�R�q�ѣG� �S�5H$E��2;|UUUt����i�x͚5q�w      �������~���ݻw@{K�;�_i(l�ҥq���p���R�)����ӧ�M7���Ơ8�ϟ��~{6D     @����gϞ����׾�ƍ�����ۂ�{������ҢE�
��=]�u��t��={f?s�O� �:o��f6D     @~�����ŋ�hz��=�P@G�4�/5S���j|���@�W%��-[E��<I�1t�t �C1̛7/�M�     @>���gΜ��y����n�Q����jkkk ����/�׿�u[�!�pU�dTѮ��җ��Ǐ�L)p߹sg ��gϞx���]�     �iy`
܋�+_�JL�4)�#u��=���}�Q ������k�o}+�������
w}VUUU|��ߵU�N�J-(�����     rbɒ%���ޭ[�x��:Cj*�,ȶ���(2�;|�U�Vŉ'�HfΜ)4�K���bI�ӭ#G�      �Wccc�&w�}w���t��Tl۶-�|;y�d�\�2�瞀"���hmm-��Y555�t�;ϢE������     ��|��,�+���y���0�cΜ9QYYPTw��6m����G��{�ѳgπ�п��z�s��P�֭�����_80      (?---�[�<��ѭ���ci Ǒ#G�7ވ�3g��,�E;�6,�L��U***����@��_x�����c�      ����_�ÇG�����m��Й�P,/��r̘1#멠���<�mp/���ߵ&t�t �C������=z      �e�Q$UUUq�}�t��}�fߩ644�{�쉍7�����H��!moomm����W��F�
�j&��xΞ=k֬�9s�      �#�w�w�"����cРA�-mq����}��Pi���������n���Q���{�(w(�ŋ��w��j-     �2��IMMM�u�]]E�Ųe˖صkW|�K_
(�;\��U�
u�ϤI�bذa�@�Ŵ������E      (}�M�6E��s�=ѳgπ�����Y�ti���?(�;\���ˣ(�u����7JE�6������� ���W_�     ��E�EkkkE
��N�Е�P<k׮��<���P$w���͛u��̙3����"]0 �;@����[q�ĉ��       J�ٳgc͚5Q$�������*�+	ܡx���������w�D��HE�B��o�=�Ԥ-�w(����X�jU<���     @�Z�lY444DQ�9�MĔ��STVVFKKK ő��x ����B�8y�d����Q3f̈�}������|@���kq���g��     �����H�+**���P
�2�~��e7c�q�ԩX�n]̞=;�(�p�+Vd�c���vJY�8�)�ްiӦ?~|      Pz6l�G����4iR�1"�T��_���
(-�S$w�?����r��(�iӦe�P��a(�4p&p     (ME�ޞ��{��$5[�n�X�m��w�[n�%���ҋߡC�����;�(Uw(�w�y'�^�o߾     @�h���(,�i*���-[?���@���H�ۧL�� FI����޽{�ٳg(����x���m�      (1i{{KKK�偔���� �i�����ODϞ=�N�����!�|��(���*0�B�8���(��˗�     JHZRdy t=ܡ�R�v�ژ3gN@�	�����Q__E�`(uw(��{���ݻ�[n	      �������ɓQ�R����mo.J�\,-�Sw�_�V��"p ���8��'�|2      �zE��>y�d�)i�����0�xv��{�쉛o�9 ������c�֭Q'N����;�����������      �Ή'bӦMQiy�]w�P�RS!p��J}SOy&p��֮]���Q�g�(w�ԩS�y��7n\      �uV�^---Q�R�w��R����G�n`��O7���"=zt:4�\����KXSSS ŕ>��      ]+�tE�n���r`i ۙ3g��wߍ)S����Bۿ�ٳ'�`֬Y�$�� M<x0��z��7�?�aTWW      �o۶mq���(����flʁ�X�r���\�Shk֬�"H��o��r�dw(����l�x�ԩ     @�[�zu��픓A�e?�---ӆ�ԩSѷo߀<�Sh���zA�ޞ^j�ܘ8��y-p     �|���ٍ�E0v�X�QS6�u�-�<v�X Ŕ\֭[��sO@	�)�]�vő#G"�w��*ʖ�߀$M744D�=     �γq��8}�t���PN�@���--��Ww
뭷ފ"�<yr���3����s��e�<��     �s�]�6�ছn�[n�%����b˖-׶m���ѣ���Kw
��{EEE̘1#�\��X�9nmm���՗w     �Γn�}�w��㎀r#hRS���?��y#p����������(Wݻw�~���G}@����������     @�{���=��ƍ(7ii �����SHil̚5+�ܥ��������{/&N�      t�7�x#�`�̙QYYPn�@�gϞؿ>< O�R�2λt�J�����QUUP�ҁl۶m��[o	�     :A���K�O�<9����D�^���?��RO!p'o����ǳ���kii�g�y&���ƦM�(7&��6��n���FEEE      �q�y�hll������޽{���T�޽;�b{��7㡇
��;��~��,�+�ӧO����cŊ1jԨ,t7n��(w�ͩS�bǎ1z��      ��M�E0cƌ�rV[[+p��>���;����Q���oߞ=}���I�&e�����2�;p��9.p     �8is��"�7�tS@9�T m�pڷ��퀼�S(�Ν�-[�Dѥ���S.�@FϞ=���> R��裏      c�ƍ���y�������M>E��m�|�M�;���By���ȝ�.��>hР�:ujL�2%jjjJI:��ٳ' ҵZG�ͮ�     ������Q)ܴiS�����ٳc�������@��;wƉ'b��y p�P��W��رc�hѢX�dI�;6�Ꞷ�WTTt5�;p��5dΜ9     @�J���w1E�n_�n]��F"������
(i�e�ymnn���g��⮻�
��;��6����o:��'Eœ'O�6����;���8.�6i�     �ߎ;��ɓQ4)
ܾ}{����7&M�ӧO�������s�n�H������8t�P9r$�z�?���}�ҥ1f̘lRy�����Up��6o�---QYY      ���ݩS�b���bŊO���7�wS����R�$ipcccTWW�;�;����r}���>��B�4�<eʔ�޽{@gH�1�6gϞ��;w�     hg��Npޅ[�S�N�Z�����R����$���!�l�uuu�N�Na��$n��Çc޼y�x��?~|̘1#�Б�]���� I�\�     ���Ǐ�޽{��;v,-ZK�.�1c�d[�}WE�����6�6�;y p�ZZZ��$�O��Z�n]��1";�M�8��&t�����ȑ#�����      �ǆ���|����ظqc���ٓ'O�z�^�zt����&��7P���Ν;��ٳA�طo_�,\�0���5kV2$�=���h��������={      7nӦM��K�_���˖-����ǌ3bذa�m����&}>����N�N!l޼9�x)4�p�{
��!.m߆��Pssslݺ5��     �ƴ��h+�SCC�E�D��>q�Ĩ�����޽{[�	|"�͙3'��	�)�>� �\i��ܹs���mWr80�z	܁K��w�;     ������̙3��I�DzR+QWW�-2dH@GKME�s����{wʞ���KS�۶m���ӧc���bŊ5jT��7.*++�����6     ���6��~���?��~뭷f��رc���*�#܁����Y7�ѣ�	�ɽ��t����ؾ}{����7&M�3f̈���\�����v�ܙ]�أG�      ���M�t�ԭ��O�>1y��>}z0 �=���@��g�fM��ѣʕ���۲eKPZN�:�mu_�re�9�Vw�J
X�pD��H���cǎٶ      �Ϲs�eut�ӧOg�Ċ+bԨQZ	�U��p���]�N9��{|�AP��5(m[�S�N�)S�DMMM������P���     \���}SSS�9Z[[��;�;p�����
(Wwr-
�m���cǎŢE�bɒ%Y��&���rEEE@�t Kۚ�lݺ5      �~v��e���ѭ[7�*�'� UsssTUU�#�;�v���8s�LP>҇�ƍ�'�̓'OΦ�{��`���Ν;�A\�     p}҆W�֕Z�����+�j��KS�Z)����!>���lp
ʑ��\KSH��#G�d��K�.�1c�d��ѣG�%p.U__��n�)      �6i۳[�K˅�D]]]̞=;��ERS!p.����+�;����@�6�<bĈ,t�0aBt��=(�;p%i�M�     p�RW������J�_�>{�Z��'Fuuu�������>�������ʑ��\��Ͼ}��g��1~���1cF6,(�~��e��Ν�6�����      ��֭[����J,\�0��>k֬2dH��,.�>�[[[���"���ɭ4a�w�� �bݺu�cR�8��V�8޿ �1�     p}�m������OZ�[o�5�ǎUUUw�R�q�Y��ʍ���ڽ{wv]�gR�XҁL�\(���~�׳g�      ���ܹ3(O~�a����'&O�ӧO��%p�$-�S���֮]��b�pR9}(��}���&�sƁ�T�NkϞ=�|%      �:��S�N����ӱ|��X�bE�5*�M��ƍ���ʠX�B�4�~& ڤ���;�(7wr+mp���F��s�f[�Ӥr:�80(w�J���     ��m߾=ȏ�*�w��~���ԩScƌQSSGmm�����{ʕ���J�0�I���Wb�     �ڤ����ɓ'c�ҥ�lٲ;vl�J�f���"ȷ�T�ڵ+ ڤE�����-PN��RSSS�߿?�ͅ��}���I�&e������K�6N
---��`     ��ٹsg�o��ͱq���I���ɓ�ؽW�^A>Y\*us�3?<A9��K)nO�;\ɩS����+W���#G��ٳ��n3�\&�u��cǎ@�����w      �/��{��	��ȑ#�hѢl�{]]]�J><��;p%�f�;�FD.�޽;����m[�S�N�)S�DMMMP�ҁL�\����[n�%      �|�{���Ơx��j�ׯϞ#Fd�'L�ݻw�_mmm \JOI9��K{���)�n�T3fLv�5j���%*�[�l	��۷O�     p>��À��Zz.\�mu�5kV2$(_�n�N� m|�S���R�4��^�7nܘ=)��<yr����+(�����?     �ձɕ���Ǻu�'muO����㣪�*(/i��A��СC�&�����=z�(wr)M�:r��e[�G�t=�;p%>�     ����ϒ�s�;wn��=-�>}z0 (���jmm�={�ė���r!p'wҤщ'�˅[�Ӥr
�'L�ݻw�����     �X���|�ӧO����cŊ1jԨ��7n\TVV�MS\I���SN��N�$M�1���+=,Ȯ�1cF6,�\�{�Ξ�g�@�ÇGcccTWW      W�n3������پ}{����/�N���555Ai����K��PN���t�tS��u벧m��ĉE��h����k׮ h�~�v�����[     �+KK��z�<y2�.]˖-��c�f�D��^QQ�܁+�URn��N
۠3�mu_�pa���ŬY�bȐ!A�J2�;p)�;     ���q����c�ƍٓ���<yr����+�z鿓4t���1�F���;�
�
�
�����zk���媪����R��Ç      �M�N{:r�H,Z�(��>f̘�={��T]�G�ѧO�8u�T �9{�l|��Gѿ��r p'w�m��?�0{���S�L�&��ܸt�َ;b�޽�?\�{      �������>��>bĈ���0aBt��=�|i����TzаQ.��J�ZG�F)I���^{-�/_��v[v�K������;v,�y�x�������y��     ��RW�{W:ھ}��g�QWW�f͊!C��'��J7�;6��ɕt�FCCC@�iii�͛7gπb�ԩٓ���r�*�?�U�VŮ]��j	�     >�ѣGut����X�n]����)t?~|TUU���6 .�ʉ��\���rp�ĉX�xq����D\��>j�([��|ؾiӦX�dI9r$ ��ɓ'�_����3      �����B�<w��l���ɓc���ق@:F��p)K)'wrE�N9inn��7fO��M�{:����;�(f_z�ػwo ܈4 s��7      �U��N�>˗/��+W�m�ݖ��_��W,l'�q��yǎp)���;�r�ر�r���[�`A�ٽ��.��o���(�������իWGKKK ܨ�w��     �r�6JE�6oޜ=�:�)S�DMMMpm�����~l۶-8���p%��lll����R'p'W{�_�>{��M*O�81z��y��,?����0@{9~�x      p�C�����ޢE�bɒ%1nܸ��9rd��Μ9o��F֗襀��`R�5|���R'p'Wm����㥗^��_~9ƌ�f���V�49���OG}}} �'��     �2�)e��ͱaÆ�<xp�O�4)z�����G�k�����i�"��J�wʁ��\��G�@�q���馛���������u��e�~�r��	�     .׶��A
0�͛���J�H�VbĈQT�t��x��ׅ��1�F���+w�n�޽�3��� 7s��:th����z+^|���' ��      �������ƀrr�ܹx��7�'/K��{���_�ԩSp���;�q��٨��(�4�����'M(O�6-&N�X���?����v�C��     p9ߡP���Z�����~����^,�\�ɍ4iE�o߾�I��)S�d���A��Լ����v�S�w��wMEEE      p����h[
����92��>v�ب����H���ٴ�;���;�!p���-+V���+WƨQ��нTp{��^xA�t������Ě��      �<[ɛ� �ر#{�����R�D9���������<ڛ�ʅ���8u�T �p۷oϞt��<yr6��U�3g�ğ���,8�,'O��     \@�F��>}:�-[˗/�d)�q㢲�2�I���z�8w�\ t��Y��c�w�P���F
ـ��\:����]q�K��s�=��'��ҁl���     �yǎȻ��E���H��ӂ�R�u��ls{SSS t�4�6t�ЀR&p'7lp���U�%K�Ķm����     �؉'�$�̿��+�t��;vl�J��Qj����ӟ��@��S�䆐�N�.���v[̚5�Cp��6�t�      �ST��ͱq��쩭��N�:5z���������SOŹs��3|��G�N�Nn��צ��%6oޜ=�}�K��͛����     �������ѣ�hѢl���1c���G��?��x����:���r p'7Μ9��i�����cǎ�U�      |��ٳ����yMMM�lu1bD�IL�0!�w�ީ�>R��k׮ �L'O�(uwr#ƀs�n�С1}���8qb�����5���c�Е�      |ʦV�l���˞�:L�4)k%���w7o��V�
��潀r p'7�lо</��R����QWW�gώ�Ç�?o͚56']��?      γ��XZ藚���muOK������VCCC������ ��{�@�Nnܡc����ׯϞ/��+]i�v�� �j�      >eS+\����K�,�ɓ'g������_�ҥ�\]��?��;������ �`��?~|̜93������7ް�(	w     �O�>}:�k���,_�<V�X�F��B�q��Eee�u�k>|��@�K	�)wrA��+]��nݺ�i��^WW�W��R��      �S���imm��۷gO߾}cҤI1cƌ�߿�5�k��/���� �*�
ʁ��\����k�mu�?�������      ����O�|����Z�*ƎӧO��#GFEE��s�n�;v�����������m����¹s��Z�v��455e[��H      ygS+����}�ƍ�S[[S�L��S�F�޽?�bŊ �j��H�o555�J�N.����X��޽{      ��б�=�-��K�Ƙ1cbڴi1z���w���g{;P2����R&p'� ������      �̙3t�t�t�V��Ç����c	���+W��R�vJ���\� ��~      p�������/��B,\�0���bӦMP*�P��䂀 �Tccc      ���@ר���u��@)�n@���w �R�      ��	 p!��:�;����  ��     �< p!��:�;����  jmm      Dl �żP��䂀 �Tsss      ��[ �bwJ���\�� ���     ����&ߛ  �S��䂃 p)�      6 �rnw��	�� p)�      �3 .���P���� p)�      �3 .���P���BEEE  \��     �� ���:�;�PYY  �~      `C+ p9p�:�;� ` .��      ��V �rwJ���\� ����
     ��� ��~@���w �R       ��Z[[J���\� ���     @S \���N�N.� �K9�     �� ����R'p'�u� \�{��     Pt6 �R�(u�`rA� \��     �� ���J���\� ����     ��� ��~@���w �R�      l �媪�J���\� ��~      ѭ�< ����R��\� J�H�      "��� �B�KJ���\�ѣG  ��ٳg      p~1P�����  ���R'p'z��  m�      |*Elw ����R'p'��4q���  w     �O����ٳ ��)uwr���"z��gΜ	  �;     ��Dl �����J����H!�� H��      �	��y7��	���Z�6�      >e9 p!]�N�Nn8� m�      |J� \HWA���}�� ��_�~     �y"6 �B��(uwrC� �1�     �) p!��:�;�!d �|     ��� hӭ[��޽{@)��B6 ���7     �O���+  ���;�!d �|     �TMMM  $nv���! ЦO�>     �y�
 �M���J�����. ��I����      ༾}� @⽀r p'7R�^YY--- נA�     �O�� ��^@9��)nO����� (.�;     ��Ҧ֊��hmm ��lp��ɕ�
����      ����޽{Ǚ3g (6�)wr%m۷o ����      K1�� ���r p'Wm ��     ��0 ��� @��*(wr�_� ��     ��� ����y��u�����0�0�30ð�"��b�7�D��W�TJ��m;��{�U7�][��ʹ�̫�l�i'��Ina*����2��,2���t��PYf�.��9�3�R�����|>���xO@>�SP (n���     �_�իW  ŭ[�nQSS���A ����l{M      ��i� @z?PRR����������  �O�{      ��� ���B�NAi�ںq��  ���\      vM� x?@��Sp���#p�"%p     �5[ ��w
N
����? P|�      �VYY555�y��  ����|!p��� (NMMM     ����B� �K_I��Sp��� @q�>      �ͥ���V�
 �8	��w
�� �SUUU���      ��w �8UTTDMMM@>�Spz�oݺ5 ��a�     �[3� �WZ�VRR����ܷo�xꩧ (���      ޜ� ���\�'w
R��*p��b�;     �[K������  ����|"p� ��
 �ǅ     �[�������ظqc  �EWA>�S���� (.��      o/�@�18�|"p� 4( ��&����      o-Mo}�� (�������/�����,tkii	 ��80      x{)p �KCCC�����;+Mq�@q�     ��; ������;+�n<�@  �O�     �{R�VRR��� �;�F�N��@�H;�      ��z����/ P����;k��� �����ݻw      �{R�&p��ap �F�N��իW���EKKK  �k�С�6�      ���w�} ���J��;w
Z
�V�X @�J�{      v�)� P<�y��@����&p��'p     �3w (�7w
�� 
[Za�|     �gjjj���.ZZZ (lw����6dȐ(--��;w Px���UUU     ��IM��~��  
����#�;�{��1`��X�fM  ��E     ��I�Y� P��������|#p���9R� *��     �sÆ ���m%%%�F�N�K��w� @�5jT      ������s��  
S
�!	�)x)pO+�Z[[ (������      칊���߿�]�6 ��d�����WSS}���u�� P8Lo     �7i��� 
S<dȐ�|$p�(�)�w (,��     ��1bD�� ��������H�NQH^�_ P8�      ��� (\���|%p�(�3&�n���5 ��WWW��4     `����;;^|��  
��l�3�;Ea�������X�fM  �o�ر     ��K�� 
���|&p�h�)�w (w     �����˗ P8���uuu�J�N�H!��� @~+))�ѣG      ��tW (<���;�;EcĈQ^^۷o  577GMMM      ���	�--- ����? �	�))nO��ʕ+ �_iW      �Ϙ1c�W��U  ����$F��������� ϥ�9      �G� �c��ѳgπ|&p��p�q�7 ��z��Ç      �O�A7M{mmm  ���k�������hjj��> ��������      ��&���v��  ���B p��L�81~� �&L�      ��4�]� ����<F������	� ����f�     h)p���� �_#F���ݻ�;�;E'�N����-[� �?����     @�5jT���#^}��  �S �@�N�i����_�: ��1q��      �c���Ř1c���  ?	�)w���,p�<���      t��	� ?���/���P��q��EEEElݺ5 ��7hРhhh      :N
�KJJ���5 ��bz;�D�NQ�޽{�[u ���v     ��WSSC��'�x" ��"p���)Z)��@~8蠃     ��7q�D�; 䙪��>|x@��S��Yyyyl߾= ��5`���۷o      �����[n�% ��q�DYYY@��S�***bܸq���. �ܕn�     �9����_�~�nݺ  򃶂B#p��r�!w �qS�L	      :O��~�� ��*++c̘1�D�NQK�r���#^}��  r�СC�O�>     @��@��0aB����;E-����}��� 䞴�
      ����9B�~��  r[Z��F�Nћ2e�� rPIIIL�4)      �|tP�v�m ��ݻǸq�
����7f̘����M�6 �;F�uuu     @�K;�
� �p�QQQPh�������?�i  �c�ԩ     @�8p`���?�}��  rӔ)S
����a�&p��V|��     @�I���� �{���b�ر�H��k��1hРx�� �z�'O��     @KSao���hmm  ����[70��o6���ӧ� G��U      �Z1t��x�' �-i�(Tw�?i����Ŏ; �:MMM1lذ      �륞B� ����>F�P������������ t���JIII      ����3m�4mM�o0c��; t�����"     �ܐN�81��  r���B'p�7=zt455���? @�;�����.      �i^�; 䆑#GF߾}
��� m�q���M7� @�{�;�      �q��E}}}lܸ1 ����A����8����[o��۷ �yc���      rKiiiL�2%n��  �NEEE|���N����:&M�˗/ ����i7      rOx��Gkkk  ]c���QYYP��)��@�)//��     @kjj�Q�F����  ��GP�Æ�!C���ի �xiK˴�
      �+Euw ����Y��@�o��|g|��_ ���.      ������hii	 �s͜93�X��ML�<9n��fe ��ƌ��2      ���������G?�Q  ����29䐀b!p�7�.���Z��zk  ��v     ���Z���Ǳs��  :ǴiӲ�����B�(�����ؾ}{  �O�>1a       ?���g�w���  :Gj����-���Ĕ)S⮻�
 �����%%%     @�H�x� �9ƌ(&wx�gώ��;Z[[ h?���1}��       ��=:���c�ڵ t�#�<2����m455Ł+V� �������       ��)��^{m  �O�>1~���b#p�����w hG)l�9sf      ���N���rKlڴ) ��������;�!C�ĨQ���G `�͘1#���     ��ԭ[�����  �_UUUz��H��)Mq���+++�V     ��Ҏ���~{l߾= ����UTT#�;즱c����c͚5 콴]e�^�     ��V[[�M���/~ @�I;�H1��n*))��s��W���  �Niii�+
      �a���q�w�Ν; hӧO��={+�;�<0���c�ڵ �iӦESSS      P����{�7 �}��}���L�{ Mq�7o�)� �Lo     (L�z׻ⷿ�m��� �o�±>}�3�;�!S�`�L�2��v     ��:�ѣG�ʕ+ �7�sL@���JS��ΝW\qE  �'Mo�3gN      P��=�X�; �������������A�5k� ���M�fz;     @>|x�5*}��  ����'w�i������K_�R  o�[�n��'      �4��s��\  {nܸqق1@�{-mb�1 ��#�8"     �:
- ����/���K.�$ �]����w��]     @qH;�
�`ό;6F����a��@&L�>�`  ��#�����      �8�=:F��=�X  �g޼y����Q����CEkkk  Q]]�sL      P\�?����K x{'N̆�!p�}����zh�}�� �EZ]ܣG�      ���Ho	��� ��JJJ���~w M���㎋�����u��  "�#�      �S����CEkkk  �v�!�����kwhuuuq��G�~��  "N<�����[M     �b5`���<yr��7�	 ��ű���SA;�={v�u�]�q�� �b6jԨ8��     ��6��X�bE�ر# ��v�a�E�>}�{wh'ݻw�VS]{� Ū��$.\      ����~x���? �/***b�ܹ���ѡ��]�=��� �(�      �̛7/��x��W ��c�9&����5�;�����X�hQ\r�%��� PL*++�m&     �MMMM��]o�9 ������>:�7'p�v6lذ�:uj,_�< �����={      �ёG���/�^ (vix`EEE oN�`��q����^��ѯ_��9sf      ���֭[w�qq�UW ��ƴi�xkw� ���1gΜ�馛 ��I'�eee      �2y����OO>�d @�:�����$��&p���׺��cݺu �,݌;vl      ��I1ߢE��3��L��� �I�&�������CISl/^����\�P�*++���      �vӧO���+ �����ǂ�=w�@#G�ta@A;��㣮�.      `w��K+V��-[� �9s�D�޽�=w�`i��<�7o ($C��#�8"      `w���ļy����n @1hhh���>:��'p�V]].����: �P���Ʃ���}     �=1k֬���c�ڵ ���O���� v��:�ԩS�W��U<��# �ਣ���      �4DiѢEq饗Fkkk @�?~|L�81�=#p�NPRR��vZ�˿�Klݺ5  ����Ҷ�      ��F��vX�y� ��{��ق.`�	ܡ����;�ϟ7�pC @�J���8㌨��      �'�pB����y�� �Bs�q�eC�='p�N4k֬����� �G3gΌ�#G      ����X�pa\}�� ����9���#p�N���.Y�$>��O���� �I�n$      �^�M�˗/��+W ��	.^�8����;w�dMMM��w�;n�� �|�v�UYY      О���d��m� �����aÆ�����:�x���� �3f̈q��      ��>}��q�7�xc @>�ݻw̟??�}#p�.PZZg�}v���klٲ%  �544Ă      :ʑG+V���<  ���Ē%K���"�}#p�.R__��̮�� �\ն(���2      ���(��N�O~�}�� �|3cƌ3fL �N�]�����S��=�� ���̙Æ      �hMMM1o޼����� �|RWW�| �C�]lѢE�jժذaC @.4hP�     @g9�cbŊ�z�� �|�v!Y�dITUU�>���z��g�uV\z饱s�� �\PQQK�.����      ��RZZ�=������k�� ��f̘�Ǐ���!><�����   �r�)��      ��c��o}+  �544Ăh_w�s�΍������O t�I�&����      �J����#�Ľ�� ��Ү#g�}vTVVо�#�Nv���'m�@�I+��,Y      ��/^�V���7 �9s�İa�hw�!)*<���k�	 �lm��z��      �ժ�����O�/|���� �+��@��C��>}z���=�� Й�?�x+�     �)cƌ���:*~� 䂊��l�`YYY C�9hɒ%�nݺx�� :�ĉ�裏      �5���φ�Y�& ����=�� :��rPyyy��}�O}�S��+� t�޽{�g�%%%      ��[�n٤�O�ӱm۶ ��2y��6mZ K�9*ņ�sN|�_��;w t��EU���      ��_�~�`������ �cɒ%t<�;�1c�Ĝ9s�?�A @G8�SbРA      ���xG<����� t���HX[YY@��C��7o^<��S��� ���;,?��      �|PRRg�yf|�ӟ�^x! ���x�1x�� :��r\�8;묳�3��L�_�> �=6,���      䓪��x������gc۶m m���1s�� :����/ζn� �/jkk��s�Ͷ�     �|�����zj|��_ �HMMM�dɒ :��	�Ā��UW] ����ʲ����>       _M�:5�x���� �***������t.�;�C9$�8��; �ƢE�b�ȑ      ���O�5k�ĪU� ���ŋ���t>�;䙅Ƴ�>�<�H ���5kV̘1#      �t��-����O}*ZZZ ��QG��t�;䙲��8��ⳟ�l���7n\�t�I      ����6�=�������رcG ��=zt,X� ��#p�<TYY\pA�ۿ�[l޼9 ����/�9�(--      (4Ç�N8!���� �޽{�ҥK5���m�.��2+�xS��_�(�G�      ���#��5k�į~�� ��Q^^�}�{���&��%p�<6bĈX�xq\s�5 +]x-[�,      
ݢE���}�ڵ {���$N?��<xp ]O�yn�����K/����� �6��묳Ί�C�      ����x������g���% `w͛7/9� r��
@:�n޼9~�� $'�tR|��      Ť��.�?�����Kc۶m ogҤI1w�� r��
��'�7n���? (n�gώw��      �h���q�gƕW^��� ofȐ!q�gDIII �C����4�.]�]vY<��@qJ�e��      �,�v|��ƭ�� �+�{��.� �w�@n�CI'ڴ�ֿ������? �1c�XU      �gΜ9�~��X�|y �UUUŲeˢ��6��#p�SSS����K/�6 �aذaq�y�E�n��     @�C�v�i�y��x�� ��V���������PP����㢋.�"���� ��80����GEEE       QVV�{n|�s����~: (nm��F�@��C�jll�}�CY�iӦ �0555�>��l�,      ��UVVf��.��X�~} P�.\S�N �	ܡ�����/�V!oٲ% (,}��/�8jkk      xs555ٮ�)r߼ys P|fΜGuT �O����9�@���?[�n 
C}}}\t�Eѳg�       �^ �lٲ�����^ �G��~�)���P��~\~��}��  ���)n�ݻw       �oȐ!�| ���/P$<��8�3���$�� p�"1z��,r��;v� �SUUU\x�ѷo�       ���������j( 
ۘ1c�sΉ��� ����رcc�ҥq�W�Ν;��RYY�Mn8p`       {�-x��+4 �mAS�nRY�7��B�9蠃���O�k���@Iq{�*q���      �<0�8㌸�ꫣ��5 (C��:���� ���дiӲUi_������_ r[UUU����aÆ      �~�N����^{���@477g�E&�'�;�ɓ'g'�~���}��  7����E]�]|      �o�����k��7� �>}�ą^����/�;����g۰|��_�.� �-={�������      �q���wƖ-[����~ ��z��u����7�;�Q�F�?��������J �z�>766   �-�رc��}�{���  @~�7o^l߾=~�� ����..��⬷ ���!C�d+׾��/��/� t��}�f�����  @�Ν;�)z)"O1y�ұu���{���j�1}���g?���?���f?�>�}�~����+�L:v���RRR��<�����]}��������O����ʲ�����\^^���+**������ا寧m�Zڞ9}���
   �����]��v�m@~HQ{�,(w 3hР�������?---@�8p`\x�QSS   �b۶m�y��?��)VOQz:R�����������):o;
͞��)�o���t�ħ�-�O1|����6��G�QYY�}La|:z�����  ���p�	����o�9 �m)j��?(n���3�g������q�e�ņ�Εv���>��,  �Ui�?��Y���+�d��H�-To��S��>���s���.$H�wW����I��c[���t��b����/�ӑ�  ��fϞ�����|ǵ-@�J�[��^WW@a�%�d��⋳�}���@�5jT\p���  �Ζ"��7f��7mڔ}�"�4a�m��`�]i�}H��ۤߛ��65>M�O�H���t�§k����,�����~  �+̜93[�{�u׹�1��/�0���;�wz��Mr����㩧�
 :�Ag�}v�0  �=�����HS�����i�)H��UڦƧ�����V�b�tݜ�����)�Oӹ��� ��2cƌ��ꫯ���F�˖-�& �I��Rz8�&����g���@ǘ5kV�|����  `w�M]O�_z�l�z�����q�6�7���w<���J���"�4>�'555ّ�u655Euuu   �C9$�ָ��+�]� �:�F��.���(pw�M������}q�-��m�� ���ϝ;7�=��   �[)�}��c���Y̛&��p�m�q���ߋt��'iǂ�������S߽{���g������eccc���  ���8qb�w�y�|E��E&L��}�{�!@a�o)m�{�	'dx����lR ��[�nq��ǔ)S  (^)T߰aC��	�i{[��A9�����?�n�����#�<��_�L������uuuY ��ܜ��  @q7n\\x�q��g�� t�ɓ'�Yg��ݿ
���-3f�Ȧ]u�U�m۶ `龜�iw��e  P�^~��l
{���D��y
kS��	���o����Y����{���o߾��  ��0r�ȸ袋�K_�R�� ����ŋg�Z�� pv���G���i� {&톱lٲ��7  P8R��nݺ,do�طnݚM��C�x��==\M�{eee���D}}}455e���  Px���ǲ���� :��ٳ��㏏��� ����#i+ޏ~���E�ڵk��3|��8���  @~j�ƞ\��5}�B���-�Ȑ��#-tI�N|���{m����o�l�{�>}b���Y  �4�*	��W��=�X о�@�E��G@��{,=����?W^ye<����[�>}z�UV�n�z @>x�����"���]
ٷmۖ� {ꍓ�7l��?�x�}���C�4ݽ��*jkk��}����W   ?TWW�E]���7�7��M �>***b�ҥ1q�� ���
�+i�������w◿�e ��҃�M�1�  @nI�z�ľnݺ,dO�_}��,d��u(E��H�C�W�ξ��'���)|�ٳg444D������>  �ܓ�\�}���{��o�= �7i�\C�	�x	܁��.�N=��l;���ر# ��4�!�&;vl   ]+E�)f_�vm����iӦؾ}{���@�I�{Zp�����O<��雷��!occc6�}РAv� �PRR,��}��u�]�����K���-[�{�����	�3fdo.��կf��]�q�v�hjj
  �s������3�ĳ�>�MD~�W���bv��;6lȎ�+Wf_K�{Zh��E�E�555  t��;,z���i�& v_ x��F�=@����Ç�'>��"��'��b5q��l����   :N�p�~��x����---ٴ��u�b�v������W��_���QZZ�ݛ�������)~O_  :֘1c������/����Ҁ�E�EYYY $w�ݤ�%_|q|��ߎ��+ �Iz@<��8�c�- ���&�=��ӱnݺظqc6�=M1`��b�-[�dG��"I�+***���6��{���!z ����k�E�k׮ v-ݗ8餓b֬Y�Fw�]����i���F��믿>�n� �.m�����i  ��IQ�3�<�=�}�bӦM�}��hmm �^zM�ґv�X�re��{�)zoll�"��  �������h|�[ߊ�˗ ���:�9���Kw�CL�6-W\qE6]�P�92���ٳg   {��_�5k����?---ٴa1;@�H��iG�6dG�������l�Φ��>|x��  �siA�g�����[n�%[�@Dsss�w�y��� �"p:L�~�������7��{��B�&��-�.\eee  �������g��B�W^yŃ]��^���u:����+�{��_6�2�9C���ݻ  ���s�ٳgg1�UW]���(f�'O��N;-***��܁�&����&L�뮻.����Բ�O?={m  v-��<�L�]�6�ξiӦx���Mg�C�����cv�^�:����֭[���fS��i�;  �k�ƍˆ~�+_�u��@�I��ϟ�sL���܁N1mڴ<xp|�k_�n�ѣGǙg��m�  �EKKK�Z�*���H��
ێ;⥗^ʎ�+Wf�{��My4hP6̔w  �i��'>�����w�uW �4H�Ί�c������_�~�},n����; ����s�̉y��YI  ���_�'�x"�8����۷{�P��[�lɎ��i���Q^^�MyO������a6  ��>���N�Q�Fŷ����
@!9rd,]�� A`�܁N�.�N>��1bDv��v ����8��c�С  ��瞋'�|2��&����� o%�:iAT:~��(++�"�4�r����=  (VӦM�����W\6l�B��̚5+.\�� �w�KL�4)[�w�5��C= �*�XZ�hQTVV  ��;w��ի㩧��^x!^~��l2/ �tٱcGlܸ1;y��Awuuu���7���=i=  (������o|#x�� (UUUq�g� {C�t��5�e���;�o�1�n� �"M[�d��-  ��k�����O?�t6e7�&h���sMZD���gG
�{���{�����l�{�ne P�Ң���??k'n��l'$�|6t��X�ti444��rW�R�Ō3bĈq��Wg��ڸq����O��={  �m۶ţ�>�]����K�� ��R�Y�c͚5�|��lW����6lX6�҄w  
Q[;�y~�k_�g�}6 �Mz-�5kV,\�0���`_܁�Я_���G>?�я��?�q�U-@gK[d�x�1}��  �B�s��X�zu�Z�*^x�x��W r]
��9+�0����<M��۷o�92���  
I������x�|��q�w@�������>;�^hw g��{�{lL�4)�����;@g?~|�z��E  ��{.{�X�n]����Y$ �,���9���ώ4�}����>}�Ę1c�w��  ����<N>��l����_���J ��z-^�8[��^�@�I+��4����gq�-��&�Pij�	'��m�  ����%�׮]��9Mm�B��u�6mʎ��gϞ1`��;vlv�  ���ɓcԨQq��ƃ> ����2.\�� :���I�AđG�=���7��m����M�SN9%jjj  ��k����|O=�T��⋱}�� �b����7f�C=�M�L��<8�"�{��  ����6.������;��o��[�@.H�L�y���� A��~��Ň?���{�������v����-����  �;vd�W�^��h�[K��֯_���{o6ѽO�>1bĈl�;  䃒��l:rZ�y��Wg�� �JZL>��lpiz}�(w �7CӦM˦��t�M�|�� �iw��3gf[  ����%��Ӕ�M�6Ekkk  {.�C� �'�|2;��ʲi�)tOCҶ�  �������G�g?�Y|�{�3� �tÆ��N;-X
���@�H��6ӧO�뮻.��� �]��SO=5ے  r�Ν;�)\�V�ʮ{�m�&j�����ƍ�㡇���7���  �4�+MM�8qb\{��裏@GKSۏ=��8�裳�!�� p���������w�qG���?�*xK���1w�ܘ5k�-  r�k��+W�����	����q:�#�C����&Ӎ92�w�  �KҢ�}�Cq�wƍ7ި� :̈#���MMMЙ�@^J+gϞS�L�[n�%�/_ o�Dv�a1���o��  r�s�=�E��֭�W_}5 �ܑvTy�����{�=zD���c�رѫW�  �\PRR3f̈ѣG���_������TUUł��"�� t6�;����3�<3=�и���g��Q���;}������Ir��@¾( ⾡�(�-ڷ��u{z��{k��<�5U��>������wf����]^���Kk7����l�����dO���"\�n[� Y^/�S�sN�]b��������]���/bٲe  S���H�2��ѣq� `�K;���Ç�TTT��ʕ+�;�c   7]js������O���������C<��C���Q__ 7��;0#������x�w�W^�7��g������<_l �ͦ� f����hooϓ������˗�]wݕ��  �f���{c͚5���/��o��k|)s�w�w��fpf�Ԝ�e˖x����^�m۶��̗n��_�U���?����  ����ɓq���8w�\ 0s��Pooo�۷/O�X�%K��}�ݗw �-�7M;]�_�>������� �&�,�y�x��d.�)C��q�[jp~����׿�u�޽��d���Л6m������5  7���D?~<:�C�Z��522��Z[[s!KKKKn�[�ti  ���z���?���Ď;b�֭��� �w���?��X�hQ L%����`���������/⥗^�#G�03���Ń>���.  ��R�=]k<x0:::,� �&������ӧ�{SSS�~��  7B���aÆ��{����w�ɟk$)W������{�7 �"w`ƻ��������y���q�ĉ ���z����+W�  �QR#�}������^�v ���^��������X�vm��:�P  �S]]]����a�_��q��� f����x��b˖-yA6�T�;0k�P���_�+v��������`����[�g?�Y�[�.  �FH[7��q������ �*5fvvv�����>����X�jU�y�Q,  ��T �?����O>�$����3!0{�]}�������FCCC Lu����N�z衸�����W_}�ELq��rK������y  p�uww��Z[[��ŋ p��a��0�q�ݻ77k.[�,o_[[  p=��ʹ���wߍ������ f�T
���ݿ�ל Ӆ�;0+�����?7n�?�0^y���0Ť��-փ>��  ��r�,;u�T��� �����i�����s�=5�����  L����x���G�!���{/����Y�,Y���w�uW L7������6l�[��޽;~��Ĺs��y�/_?��O� �������>�� L9)��O>���<W��iS� ��T__���>�l�������>&&&�ޚ��r��M��P(�t$�P�B�=�PԦ�������8�W�������7�  �zHA�O>�D� �V�¼49�~��w��M  ����������ǹ�=�����2gΜ�`%��\YY әO� �"�S�6��Ç㷿�m? �G�o.m��V�z�  �mdd$���G����^7� �i-��|��Ǳw��ܶy���wܡ� �I�dɒ������Yگ��8t�P S_]]]<��39�^UU 3��;�7X�fM��G��믿�oB��H+�7nܘ/�,X  0�FGGs�i����  3M��:��?����裏���1֮]��v��;  ?X�}��������lꩧ�駟���� �I��E����������.�{ｼ%,�ݥ-�7oޜ/���X  0Y&&&�/�����7���"�uvv����cǎ9�~��w�1 ��J1`*�x���a�lfw�k4������=�\n�y��7��ٳ|��˗Ǐ~��ذaCno ����P{
u��  �ٕ������������sO,^�8  ��J�������Y�?��?������R�`
�?��Q]] 3��;�w�N�x�x��������o�>��GR�������  L����ػwo���� |����8}�t��Y݊+���"  ��m������?�{�7b�Ν>�� �r���?�y�b� ���;��TVV��w_����x��r+N___�l�Z����{,���  &C�ٳ'Z[[cxx8  �v���q�ȑ<i��U�V����n ��-[�,���/���ױm۶��H���J��=��3��#�D�P��ħV �`޼y���?�i\���C�iug�H7��b��Zxݺuy  �P��)mw|������u� 0	��>�;��϶��޸��[  ���*��_�"g%R!�R@��R�⮻�-[��w� ���;�$J!߇~8OWWWގ�w��]ttt�D�/��7jk `R�<y2>��hoo��1 �u��ϱS����}��ʡw  �.���ڵ+�x�hkk�ڥ������'?�I,Y�$ f;w�뤱�1�t>��q�������w�-�^]]]��jӦM�|��  ����ߟw�jmm����  ��ˋ�TWWǚ5kr�{�X  �V)��aÆ<iWƷ�z+>��S%�455œO>�?�x�c p��;�u��Z�n]�����sn!����������Aeee��*}q�}��&  ����F_|񅭋 ���������yZjsO�m�~��  �ŕ�Dwww�ر#�~���/Y�'�x"x��(
��I��@)$��xM��}�Q�ܹ3�=�����$������֞ښ���  &CjM�ϝ;�Z `�J�i)��}�����c��9x���  p�Ңɟ��'��3�䅔��=���\�٨��!6n��7o���� �L��&����[�I7	҅\
x���Y���S������O `2����ȷ��-��� ��#���>}:OMMM�^�:�X,  �Ej�N�i�����C^L�>7��,�ݿ����������o'�0466�m��������w
�sݥ�P�b���{�'���  &Kڱj�޽q�  `��E-����m�i��e˖  \��;��~���������������H�L�p��x��cӦM��� |7� SLڎ(mE�fxx8��S�{
���;L����JS{
�WUU  L����سgO�kk ��.]��w'}��7���2V�\�<�Vw  �YYYY�q�y����s��������|��9s������Q��
��O�`
K��+[t����]9r$>���܎s�ԩ�k������[sC{�J  \�� f����8|�p�[�;  �G]]]<��Sy�B��螚�O�80���)׳aÆ\4XQ!�	0|7�&R@���n����<����СC�����{�����?����ijkk  &��v  ��� �dhll���~:O[[[�ڵ+>��hoo�
�5�]wݕ��w�}�y �w�i���>�(�I7R���r�=5�\�x1�]�E�ڵk�"��*���9  �z�� �_�ǭ�>�`,_�<  �H;����~�O��A���}kkk����r��ӹ������: �~�f�����u[�l�x��/��{{{��%5�_	��cz  ד�v  ��+��۶m�� ��dɒ<���Ν�ݻw�'�|ǎ��0��{��-�h0]� pc��@_�?��S�����8q�D��I�S��CUUU���n��I�v�  �(�� �_muoii�͇.  ���y�O��<i����}
����/^��{o�իW� 7��;�,���M�N��t#!��Ӷ]'O�̏Ϝ9����͕��R�=mכ��[oͫ��B  �����w�ؑ�\'  0�R�f{{{���Q]]�=x��� �����œi�g�i��������?����_2gΜX�n]nh�뮻r���O�`�J�&���i��ӧO��4)�����/��mjjʫ�.]���)؞V��� �͒�v��n�  p�ŧ�~�}�Y��tÆ���  �}����r����/����{
�wuu�[EEE�Y�&��<+V���0	�pU:�O'�i�*m�B.W�Y������٩����i��4�-ʓ��͚���  ��mbb"��I��t�  7ZZ\�>~��s�}����Y5  |W�������I����ȑ#9�~��ᜃ`f+��p�J�=S���M��o���J[Ħ���I!�+��4.\������3+�
�EUccc477�c
�/X� �׬� `*Ja��;w������=  LiWѷ�z��N��<�]/ ����C=�'I��ʡ��G�ƩS�|V:ͥ���zk�Z�*�\V�\��^|��{K7�4��9ccc9�~%����J�nN\y�&�j�T>���������;�ܹscΜ9W�ijj�Gv  ��Ԍ�k׮���ٰ( ��itt48�;bnذ!�U  `���G}4O2<<���q�رxO� )��Ԕ�멝=گ���ϟ L� \7�B"5���9�~�&�䇆�b||���tA��U��k�&կ���ɍ�W�UUUy;������+�^ ��$�?�ݻ7o��έ `�H�2�"�_|1�ׯ_+V�  �l)+�v��<W�C:M��'N��ٳg���`)ױt���Ⱦdɒ���[n��0C����q%\~��x  �ۥ�v�ܙ��l� �t�v}뭷���2V�^�<�Hޑ  ���cX�fM�+R1ߙ3gr���Ǵý�����-�b�r�%�]�   f�tCe׮]����
  3���h8p <��.6l���  p#������R�=���?>O{{�������ei���������㦦�(++ f7w   �"5��޽;}ҍ  ���bδ���_�y��Ń>+V�  �R�}�ʕy�XZ��
I�����4�q
��݊Ҏ��]
�ϙ3'�9z:���tL��t�;wn �_"�   0ͥ#��=�W���  �F)��[oE�X�;�3���(
  SA
~�݇�|���n___�������ϡ����̏�1=ʏ��I�'###1666)������\���:�s��~z�����D]]]>���_�\O� ~(w   �i*x>����X��+ �����?�8>��X�fM�_�>**� `�+//ϭ�i�/_����|O�}&�%�_��W� {�g ���'9    ��ٳgc�Νy;[�v  ��R{��СC�hѢشiSn� ��L�: 3��;   �4q�ر�裏�ִ  ��I�iף�[�Fssslܸ1�ϟ    LM�    SX
��ݻ7>���  �����W^y%����G�e˖    S��;   �422���:ccc  L�K�.Eooo���Q]]�֭���?    ��   �����رcG?~<��  ����P|��Ǳo߾X�zunu/
   ��#�   0\�p!v���O�΍�  ��3::�;(�X�"6lؐ��   ���   n����������'  ��+�vSJ��/��7F}}}    p��   �ǎ������   ����R�]��_����x�Ǣ��9    ���   n��ƞ={��ŋ  Lm)����/��r466ƦM�b���   ��#�   p� ��������J����ƍc���   ��p   ��R�}׮]144  ����{{{㷿�m444�   \�    �lbb"����}�Y���  0��믿uuu�aÆX�lY    ��	�   L�+��O?�4FGG  ��R�{l۶-jjjb����jժ    ��p   ��R����>�������X   �K
���~��عsg<��ñz��    �p   ��R���?��;  ���P���{9�~�}�ŝw�    \;w   ��hdd$7�<x�jc{YYY   \��҂ؽ{��{
�   ���   �Q
�l߾=�9��  �&�:��?�����<�֭    ���;   ��Ha��ؾo߾���   �E
��ر#7��_�>V�^    �)w   �o���)|�F�  �CCC����Ǯ]���G�[n�%    ��    �g�}�w��-�   �-��}�ݼ[�ƍcɒ%   ��;   ��8p 7)��	  �����o��f�����?.   ��L�   ��/���;w���`   �H�.]�A��^{-cӦM���    ���;   0��8q"�o�}}}  p�uuu�+��MMM��}޼y   0��   �R[[[|����ӓ�  ��t�������ob���y�樫�   ��@�   �U�������}�   Lu��^�E��F����    ���  �Y���#��Qc;  0��k�3g�į~��X�ti<��Q,   `&p   f����x��w���-   ��tO�6���/cժU��c�E�P   ��D�   �������C|��� �%]�9r$Z[[��;�3    f
w   `�ٳgO�ݻ7��  f�t���Ƨ�~7n�+V   �t'�   ���}ǎ144   �E�z�w���.6o�---   0]	�   ���ӧ��ދ���   ��.]�����ꫯ�{
���;   �t#�   L[������o����  ��A����x�b�ҥ��OD�X   ��B�   �v���rc��'rx  ��K�Jmmm�����w�>�`
�    ���  �icbb"v����y~  �_���������z(n���    ���  �i��>�]�v���X   �݌���|�|�I<���x��    ���  �)�ȑ#�}��
   ~����x��ף��16o����   ��D�   ��.\�۶m����   `ruuu�o~�X�|ynt/�   0�   S���H����q���   ��:y�d��?�c�}��q���   ��&�   L{�쉏?�8���  �#]��ݻ7<�6m�e˖   ��"�   �t�O��w�y'  ��chh(�m������SOE]]]    �h�   �M��ߟ���Ν�K�.   7_ggg����bŊؼys
�    �Q�  �nbb"v�����l  ��ҵZkkk�򗿌����ڵk   �Fp   n��?�<v�����  �Ԗ�ݶo��~�insoii	   ��I�   �!.\�o��Vtww   �K��꫱hѢx��'�X,   �� �   \W###���Ɖ'��   LO��̙3�����w��ׯ   ��&�   \7{�쉏?�8���  ��abb"���G���{,�/_    �E�   �tmmm���.  ��ihh(�z�hll���z*���   ��p   &M
7���q���   `v��ꊗ^z)V�Z���B    |_�   ��سgO��U=   �˥K��ȑ#yG��<�-[    ߇�;   ������%���@   0�Ƕmۢ��9�l����   �]�   ����X�������   �U����u�ָ����{�   �k%�   |g��y�ر#��  �ϙ���={������'�����    �6�   �5����[�www ���(�]��,.Ey���𤋮����ңKQ(���2��~OMMM��}��先�?�ߚ�T�.]��|hh0.��/���h��\�M�cc1<2W�9���c� �����x��WcѢE9�^,   ���   �*�������-� 7B
�� z��cDMU1j�����*��������X�������ʊ�����b1��K�����beeT/?���,���4�QV������(��,��f�ti"�FF�>�A��O��������q������X����p������|�q�}�C�������qpp(.�fpx$�t�zKגgΜ��[���?k׮   �?G�   ���;��^��� |_��2�����p9�^S,Ɯ9�QW[uu�cMm���Du���zu�Kϋ��L�Sz^(��l������W|��dI�F��r ~xx$7��c鵡��.�P����?0�}��S������o |ccc�}��طo_lٲ%���   ��  �?��ŋ��o���� ��Ԭ^,/��,*J�k�����>�룮�&���Ŝ�ڨ)=����buMT��U�c��:7�s�
��.�{J�]������P^,�;���`i��b�_����x1zK_��틾�{�@���/��R�Z�*{���    q�    �{��ɓ]�}�eQ����XQ�ڪb4��ż��Q?gN�ח�nN���Eu����%-R�-��H3����?>1C�����w9��ן���7:�����?�zz�b�= �|i�ӑ#G��ɓ��OĲe�   @�   ���ٳ��[o��U f�BYD��<������be4ϛ��^���������S��)�\QY��򨫛�g�_x���H���F�Ł��닞��|����=�q��+�GF��a��}۶m���[�l����    f/w    ���r��ĉ��V^V��<5�Q_SM�Rp}^�K����������!���(+�����X��������DoOO���EWww\(M�����s��14< L/����[�n�x ���    f'w   ��Z[[�wމ�Q-� �EE�J��<���PW-�͹����1�4̍چ����vf����<-��_����N�����t���������	 ������裏�������F}}}    ���;   �Ri������ L-eeeQU��W����ǂbol����b�ܹ1�a^�WVU�uUUձpѢ<lhh0߻.tEǅ�����;�t��� n����x饗��;����   0{�  �,���o�ccc�͓zի*ʣ����幕}������%�����)7��k�U5�L���X�(͟���GggG�?��:���s��8���.]
 n��}w߾}q�رx�駣��)   ��O�   f����x��7�ܹsZ 7P��,��s������X�2?̟s���~^c4�+�P(��)VU��%K�|U
�w]茎��8{�|�>{.N�k����w^p]��/��W���{�t�T   `�p  �Y�O>��>�(����룼P��QWY5��+VDKsS,X� �5��ܦ�h(M]}}��	f�t���/�s�W^����=5����S9�~.�/��;��:r�H���ŏ~��X�xq    3��;   �p�����oDggg 0y*R���<�)VDS}],Y�(���4�DCSS���f�bUu,]�2��J�.��F���ўB���ƉSg�����{�!����5�ҥK㩧���   3�;+   0��ٳ'���D ��e9�>�X���X��%ZZ�������9j��@RV�5�an�[V������pt�?gϵ��3g�ę�q��#F���%�w�k��g�&��>�x�X�lY    3��;   �@]]]���G___ p�
eeQ]Q�f�,����X���Fc˂<��GyEe |W�UU�xي<|����htu���z?{6�N��ֳ�h4ƅ������ضm[,X� �~��(�   L�   0�|����'�h�)�^[Y����^U��2�9���7�,��M�R��~����EK��u�����;ݝq�T[�:s6ZO��g����� �����غuklذ!V�^   ��&�   3D����o���@ 𧊅�h���2�^����/\��_ifof��B��ۤ���˯ƅ�sq�̙hm;�J�����@���X��������3�<UUU   LO�   0ͥ��w�y'�;���K�B�I��U�cE4��Ăŋ�y�hZ�8�,��� �.����+n��ࣗ_����Ϟ��S��h�8q�\����D �V���������o�=   ��G�   ����������P �V兲��,�9iR;{�����/�����ļ��(+��I�����u�x����h�\舳�ڢ�d[n=�}�d<&,�f��������������Fuuu    Ӈ�;   LS۷o�}���l�����1��27�ϫM��K�)��/X�[�+�U0�TTV��.�s׃ǥү����8w&�N���'�TGg���؄�;0�uuu�/�7n�U�V   0=�  �4�nп��kq��� ����hHa�bE��sr�}��%_��/�B� |]ڹbn��<��'~Tzmhp :Μ�S�Nű�q�ԙ���q�w`f���{/��?���Q,   ���  `����O>�K�������<7�7�c^Ue�k��2̞Z��ļ���໫���e�n���Ãq��\�=}*�;G�NG��h���L���[�n�'�x"V�X   ��%�   �@������ 3͜b��v��U����e�}i�,^����QUS�Wޚ灍���{Ǚ�q�T[o='Ξ�����8:a�%0�6���~;�-[O=��]�   `�p  �).5��ڵ+&&&`&�/Vļ���[]����0wn,X�<O��e�]��#ޗ�Z�g�C�q�T[�i;G�����=2���������矏'�|2/^   ��"�   S���@�������� �Ϊ+�s�=Oue���F��e�p��XP�����Ԕ-_�6�#OF\�뉎3g�ܙSq���8}�;��Fcx�bL`z�7�x#V�X�7o��   S��;   LA��۷������BYngO���h����%KsC{
��76EY� �OZ��f��u���~=���v2N�8_k���C�72��`��t�R���Ư~��زeK455   p�	�  ���^��8w�\��0�ʢ�x��}^Ue4��y��h_�tY4-Xee1f��Xi^sK���=O��EǙ�q���8z�X����ޑ���q��688/��r�~��aÆ    n.w   �">����v`�+��E}UE��2Ԟϩo��V����ce�* �]��+�π4�=�9����q��X9v4��^������(�v�ԩx��g���>   ��C�   n����ضm[�8qBk;0eUʢ15�����TUV��ũ�}EnjolY �U�5��r�</MDwGG��:'����'�kh4���bd|" �����x饗��{���?   �O�   n��'O�[o����0����E]e!������U�Q����E�WFEe1 �Z���b�4���P���q��h=z,:�rؽw�nF�͗��ݻ7�;?��O���6   �G�   n��������_|���2*
e����4M���*��e+r�=Mm}C �d���������x��j�3�����cq��B\����p��<�����/ģ�>k׮   ��p  ����;^}�ոx�b �l����\S��U1��2�kkr�}��[��pC
�WS=���q��'���9��#�32�#�p���۷o��Ǐǖ-[J߳
   \_�   p�۷/v�ؑo���ee�PU�[���������@����b^KK��~��RW?7��}�G����8}�H?v,.E��Xt��rw�F:s�L��?�c�ϟ??   ��G�   n�h����ԩSq�$pcU�rK{
����ʊʘ�xq�/�uM���	 ����kb��uy����q��X�;g�z�sh4���b�96p�+��w�yg<���   \�   p��;w.��Ӎp�%5�7�TFSM1�UWFuuM��Y�lETTV L'��W�=�ēq���8}�h����sp4:��bd�nI�����hkk��{.���   �\�   pm߾=�������幩���"�VUFM]],�eu,�uu�,Yee� �� �L[�ty��6m�������#q*��ϵ�f����v .�  ��IDAT������կ~�6m�[n�%   ��#�   ����@޶���' �������,�P��Ҥ�{��h_��X�d�P; 3^Y�Wc˂<w=�1.��ę�c�v�p�8y2������`2���Ż�Ǐ�͛7G���   &��;   L�Ç�{����p=4TU�@{K]UeQW�KnY�V�M� �Vu�sc�����j����S�98]C��3<�X&Kkkklݺ5�}��hll   ��p  �I211۶m�7�&S�,����5��T��B!�6��M��V����� &���H\����xi"�FF�����t���/�����<^��x��cc��mtx�k�/�~��|��+�7)��GEŵ}��vq��,���ߓ~oR����g����/�^Q,�]"���+K�w**��+K���ǅ���π��a����h;�Ei�����04�����d��_~9x����{   ���  `ttt�k���ohL��Ծ��*Zj�Q^(����X�zmin�9s��R}���xdd8FGFJ3c�#9t�B�iF���|<r��ޛ�c�D��+/��BEy�U��9_���)9_����=�yeUuا���b�ZX�"��\���y�{{.�ݏ|���5<v��]���.]��w���S�{�X   �p  �h׮]�w��|#��Hm����_S�uUQY(�a�h_�f��vf��A���H��xh����/�P���3.ޫ.�߿r����TU�DUMm�X���t,��ǜ������yz�.��#����Cq��+�h�������[�n���z*�,Y   �w#�   ����H���q��� �!j+�cAm1Ω�b�,j���@{jkolY0SLL����`ib(����p�8<4�/�K����.)$�f���OZ�B�Ś�|��������{u
�פ�5QS[�)�?���)�Z�!υ��rн�ȡ���C�����266o��F�\�2�|��    ���;   |i���~;߰�>R����X����(���Ukr��y��(+���bbb"�.�������+K�����_̡�^O�0��"��/L\��򊨙3'�k뢦�.k��DUm�׎�����Բ0Ͻ��3���������1�;Gcpl" �U����^�����Q[�9   |;w   ���o�����*|gU�XPW�QSQ����޺:��,Yee���&��^�X��+=���)Ȟ����S㺟�L��c��ӝ�/�,�nW��W��7D]CC>
��li�Y��yx�Gq��8q�`�>v4���s����h��߮�t���/��͛cŊ   �e�   p�FFF��_���� �V�BY����9Ŋ(
�p��X�v],^ykn��)~SX�b_OiJ��t�-��{��f���y��ȅ�����I;o��{m}×���W�5u���=3C�P�f���#_D�r�{ϗ����؄�>�7�;��\�2�|��    ���g   pN�>o��F�����)��ESMe,����ұ��ZCSs��m]������itx8�sp�4����@�qOOne׾�]Z������?���Kǜz��C��q�c}Cng���,�-��ʓv�8u�p;�?�:�G��x��ą���m�&�����K/�s�=U��   ��p  �o�}��ؿ�����cAmUnl�,�EMݜ�Ծ�u���p�\�4�ep�;������+�z�s� ;�iaI���<,�ޑC�s�E��ƨO��ω�yM9���~ί���<Ο����Ç���@t�������?�[:oۺuk��G?��˗   �u�   �R[�?��?������T�r�}aij*
��u٪5��ۣe�2�L����ׯ��{R��+�'&&���Ǣ��B�?VUS�E͙�)�^z\?o���)��ea�{7>gO��C�Ǚұh$�ӌ��>�����x뭷bݺu�裏   �/�  ��hoo��^{-FFF���ʢ��2�V�cY�����s[��[WGyEe��511�C�}]]��}��0{O��t���h 3���`�<�O��������˶�yM�ϻ<�kL�B!�ܲ*���@�8|(��=:�{x,�/�f����8�O�����U��    �  �O�޽;�����N��H!��bynjo�-Fy�yjӽ��;Jsg�Ω�.R�=��s�sg>� djc�3�c�����|��J?�jJ?�����mj�y�[r|�P�<U5�q�=���:�������Pt|���;< ����u��زeK,\�0   `����݇wTס����M�����@�M��N��o��%\�Yy�ɻlc�m c�cS%��*H��4}Fq�QT�|?���b��،�>���&�    �7
��z{{599) x��4����v�Ô�phs[��־iK���S��/��>�^���� ��� &_�����[�wk�UM4�H}�"u��QB������^��{�ɑ{Jds�N<
�g��^�\N��v�ڥ_��W    ��p    �hffF~���� �4E}.m
x���jcuڶc��tu���
�!�Ĳ�g5,/���!����� ֝���_����з�{|>��?�jc����ُC�m����sniﲇ�(a��n]�B[B-d�Jd�0�?5��d}v߸q�^x�ꫯ��v    �jD�    P���ǟ�9�C v[��Ծ)��4�r��ұ][�w*��$ౕ��K�Z��f�5��Ѱ� P��ɤ��F�����DU��-�Vۻ�6������h��~c7�[����=2�+z��hr9�4��@U����;Ｃ?��Ojhh     Ն�;    �j
?~\���ہ*��m�Vȯ��Y�v�Rs{�N�U�\6���3���������̞�� ��:^,~�YC��~�
�[A�hCc�Ѿg��g��[��ܦ��G�nZ݁*�-�~��G��/~��{�
    �j��9    @U���Woo��� T'�ӴC�߶�{<�ڽK��(T�S>������4�`�ne_Z�g!��d�J11<d�ǂ5��44*Z�h߇c�r�\³ki�ԍ������Vw��YǠW�\����x���)     �w    @չy�>��s��@u��v��L۾s�Z;�	�U�������v�}~fھ�`J�|^ ����`��;��s+��D����ZM�ֽi:�'
GT�=j�����mvvV�����^{M�pX     T:�    ��r�����@u��v�é��Nu����<��_���ķavk��9 ���.l��1��~�j�#�56�n�f;��Ddo�aV��͟�?F�;P��鴎=����C     T2�    ����d��sssPC���`{�����hL���m�9]n�r��	�NNhvjB���P{.� `�Y;%=�ݺn���x�oP�q�bMM�54�s�hi���K��k�mu/��TN��i���Zt �2Y���}������;     ���;    ����̨�����|VC���nۭ�v����vm۵[ͭ��V�������v#���};��{H� JH6���ب=,Vy(��彾i���U��⟅5�?���ud�:��4���T"�\���@���u���kr�Y�    �<�    ����:{�,!G�
]5��j�e�|��:��Ӷ�����ʑͤ5;5���1;eڧ�˲�	 ʉu|��-�P��6ہ�ئ&; _M����O���߼Sm5^���$3�XJ+�+@�v�{��w�{$     ���;    �b�9sF���P�b>���E�.�y]S�:��S��)���f����� *�r|������n���?�Ge�U������?fR��m��LN��&�PY���;��������     ���;    ��Xx�=j���L.�Ц���{��Z;��s�
���R�Y���531nߧ�	 �O&����=,�áh}�wB�V�R�F�
G�_�yL��i�TMAS�M%2�X(T�B�`�\7==�    �J@�    PQfff���k��T��ˡ��W~�LÐ��W���صW��c�������F5U&ƔN& �+�󚙼o�>]�_�j�вE�-�jl�"�ǣr��ީ[W.����:L��x�Z<�z��hb)�D�  �a``�>'��k���v    �rF�    P1nݺ�s��ie�6B����)�Q��_��7�s�~���4M�|�������};�>=>j7� �,���u�F�!\W���V5���-��./夥�k��c�F�����&�3�Mf��Y;ٽ��v�=�    �rU^g�     �gΜQ� T�i�)�-��S�á֎.;�n�Q�@���=Ӄ�q�L�W.�. ��g-t�{0m�����p{lS��7����EцFFi/����)X������_��i�T���匦��
,ʙ���ѣGu��uvv
    �rD�    P�_��Z� T��a�ڭa��.���إ�/�(_ (�������Fih l�|>g��ƍ�*S�kܤ��-�k�\�����N���Һ���ijk�W[j��Jdt)�t��;P��?gϞ����t    ��p    ��������!w �/�v�9�S��m?��jԱk��w���JW:���٧�P���E Pjr��7?�F���"�Xc�xohnU��^F��Z:��=���Y��o
���x<�0���RZKټ �������k��&��-     �w    @Y�u�Ν;g��(_�a(�u�9�Q��e��kP����ҵ�$[U!�sY�LM�-�V+���>� e'��|'����T�Ԣ��m�\.��,����kia^�x����e��LN��2v�@��v�{��w�{$     倀;    ��9sF���P�L�P�߭-5^��;�n�ɶ���Ꚛ�Ҳ�R�܃i; 8=>�٩I� *K:�����=�Ex����ukq��{�{��]��RP�v�&�T"W��g��(/��wG�Ձ���)     Jw    @��f�:r���7����q���n����.>6�vt�{��T�
�#�J���1;�>1<�TbY  Tkg���	{ܸx^�O��[��ҪM[�������w�L��1��TWا-!�&�3�Jd�+uʅ��v��Y����7���     (e�    e!����T*% ���0���WNӐ��U��Աk�<>���V����)M�kr����n�`  ���_�������ݭ�{��������g5�B5Z�/��X�um5^���Y��S�t�F__�r�7d����    �j!�    (y���:~����� ���۩�W�~���s�ϯ��{յw�\n���2锦�Gii �)X���`ָu墜.��m۪���[s{�����Re���p����l*��xZ�s6�������ӡC���0/    ��    ��v��5}���e&�q��Ƨ��e?�#�~�EmپC��6-�  ��\6k/���6Vg��7�mS�q�3���tt�t��1�0T�s�����tN�񴖲݁R����w�yG�������    @)!�    (YgΜQ� ���ץ�Z�B�G���u����K;�e��XoV�njlD��jr�ҩ�  ��Y���G�����|jڲ��7�l��ޟT��A�P��E��0+Zc1���bZ�{ �+����?��~�;utt    �RA�    Pr
��>�����@y���j��~l�۴��oj�J�}��	M���M�VS�r  �/�L�^�M{8N�55�a��m���?���1T�|���MM�pw����_��a�c�TY;:}��g�9��_~Y     ��    ���H$������ J�������֧��a���Ҫ]���b�M��Z�/؁���w4;5aU  @���s���ճgT��i�Vm�ڮh�\���Y��Ǭ�{Mԩx&��4Aw��ݾ}[�ӟ�$�4    �F"�    (����裏�-��.+���V��尟�tti��_�6V'�����f&����A{,�  ����Y{�]�,�F�۶�i�6�7�|.���V�{ryI�,�vhGԯD���xJ�I��@)�����Çu��!��n    �Q�    JB__�Ξ=�B�  ��0�z�G[j��9�[;�k�/)�k/��jr��h�V&�  (����\��.�[�Z۴yk�}o��_��J�w�����F��� ����%���;z�7�    �F �    �p�}��p_YY��c��������B���Z6������hjtD�<�\  Pɲ��F���jr�C�4Vн+�Skȣ�xZӉ���#����ѣz�W�u�V    ���    6���~��q���	@�q���n����v�v��y[�v����k,�N�j��؈
��  @���LK��T��1fGا�G�iM.tJ�����'�h~~^���     뉀;    `C$�I9r���@i��훃^;h�"ؾn2�&��j  U��4���W<�hl�Fw��@I�ꫯ4;;�?��    `�p    ����رc�d2P:L�P�߭�Z��K:�����P��ݒ  P�<V�{�X��
�ǿ	��F�v�{����׿�UN'    ��c�	    XW������O�BP2C��{�V��3M�Ԗ�;���_+�VWryIc�w4^�S|  �;��w��L2�1����;���7�T(     k��;    `�\�r� J���󹴵�/��ߍ�{^����aa�d�i����'G��  x�1jWا�G��f�Y�8���jr�ӟ����&    �V�    �ũS�488( �!�s��֧��a?oli�����±zau��9M��j�������   O��4��+�i|)��)���F)
:y����G۶m     k��;    `MY>�?���1�x����S��贐l�����o�_�������>>tW�,�+  ��*��:���i4��B:' ��:�s����q�۷O     �6�    �5��dt��-,,�ƪ�����Zϣ�A�MM����75�g�x{85����ӧt2)   ���S�cNͧs^Li9�N9�F���/�s>���     XM�    kbiiI���R�� l��rK�OQ��~mh��~���-�󙝚���~��P*�   �W��T�>���tO*�+������/�i�    `5p    �������(��
���j���ﶟ�D��������)�xóI./id�OC�ohia^   �x�SaOPS9��SJt�����>�������I    ���]    V��ȈN�<�B�@�<S[j}j��e��5����ߪ���`�3�e3�;�{��5;y_+++  @i��}c>��^�������䙗�eaaA���:$��/     �w    ���q�>��s�p��ZB^5�|*>���U��_�k�~��Cx:+��éI�뻥�;}ʱ#  @Y0����b�:�K�����i噣�"�J����z����F    ��"�    X�Νӭ[����Q�ǣ��>��N�:������\n��t�jlp��'�  @yr������\v��T"# k/�˩��G�����,     �w    �s�׿����AX_u~�l�92C[������ˤS����ۚ��/   T��TGا�A�F�i�&ٙXk�BA���?���/���[     <-�    �gf]�<r�fgg`��x��V��-�������[�?)��krdHC�ojjt�~  ��e-
�����ix1��l^ ֎�������E��׿     O��;    ���R)���{J$�>�.��j|vs�%ڰI{�;�7����ZZ��ȝ>ݺ���   P]j=N��M���R9:k�֭[������      �w    �S�.L>|X�tZ�a��r9L����\�߸P8�ݿ����;���;�s���&��4t뺦���&A   T��ϥ�ש�DV#�)�9F���ؘzzz����4M    �s�    ����z{{�ϳ�;�����A�Zk�r|��$�Ш���d�~��̴�nߴ۳�   ��d���n��\_J�~qs����]�p��!��n    �S�    ��ݻwu��i
l��%+ʾ)�Q[�_.���v�!�������h��u�=�   �s��c��n��}&��շ�����{O����+��/     ~w    ��u�Ξ=��m�T�ǩ�H@��{���r���K�>+�n��G��)�%�  ���u���ks �������\��L&���_o���jkk    �!�    �YW�\��˗`�x����j���V�-�]r�����l:�{}7�`{|~N   �j��[�L*�{Ie,�VS.�ӱc��ꫯ���^     �7�    ��t��y]�~] ֆ�0�R�UK�'���_�u�.��v   �=�x�^�s)�uj,���rFv4VM>��G}�����jmm     ���;    �G�>}Zw����������?'�(��I�*��ibxH׮jvrB   �z����x��wih!��tN V��ʊ}�������     �p    ���ǏkxxX V_��T{دZϓ���ڽK�U���yݾ��[7�I�   l�ӡ]��p����\^ ��r?{����v�b�2    �#�    �Q(t��1MMM	��r�������>��F�뺺U-VV
�֝�W5=>f   �R�8��>��DF#���U��p��%�R)���    ��;    �[V�������ܜ ��w�1���Z�\󩿾�m�|��*]*����ۺ{�k%��   J�Q<�o
�U�sid1��d�E��*�~��������V    ��F�    `�f�z�w���$ �'�q�=�W��x�ﱵ���i�{0m����  @�p��:�>m
�5��T<���300`7�<xP    ��E�    �d2�w�}׾�:|N���^�w?�����ڴe�*M����{���K�NM
   (W�bֽuA=Hf5��R&_�g7::�?�P����     Չ�;    T�x<�Ç�[@x~�!��������ںw�4MU�T2��[vc{ryY   @�����85Oib9# ����:z���|�͊�    �w    �b������Q.���W�q�3���X��ٶ}�*��̴�޼��������  @er���������|RKټ <���99rD���I�    �	�@    �Rccc���U(�u:��S푀��U���MM��DU�V����{v[��ب   �j�w��[ЃdVË)e+���<��[o��^�97    �tp   �*t��]�>}�p;��Ц�G�a��Ըڶu�R9�f����Tb).   �Z��\
{���� ����L&��_��W    *w    �2�n��ٳg��B{�<Bn�:#�<ksz��r��c��I|a�����V>�    �e�������bJ��́��N�u�����
��    T6�    PE���k]�pA ���4�V�SsȻ�����e����܃iݹ~U#},�   ~D�ǩꂚLd4O���3�Tr��zzz���+�
    P��   @��z��.^�( �.�s�+��a��{m۱[�l�x����W/ivrB    ~�aHM��V��BJ�iv>�F>�Woo�^{�5���	    P��   @�r�= <�ˡ�H@��4���E7�
y����//*>?'    O��0�3��\*��Ť�y�܁'U(��G����    �<�   ��}���ꫯ�陆��oq�����jo7�~��$�Ʉ�޼��׿V:�   ���:U�j|9��Kis��r?q����?���I    ��B�    *؅���_�ӳ��;����u}_�0���[�biqAw���[ו��   `u9�� �Q����bJK�� �<+�~��I<xP---    T�    P�Ο?��ׯ��q����}j
z7���ڶ��h��NM���eMie�I   `�\��5����bJÁ�e�WO�:�����jmm    �2p   �
�駟���O �N��VW4 ��ܰ�ö����`��//��v    ���ѩ��V����BR�ivQ~�r?}������jkk    ��p   �
��'����_ ���4������߇��Wc��_�_)�&���֕/�pzJ    6��ahgԯߴ��s~�r?s�8���    �w    � 'O������Ө�[��A;��ںw�4ׯ=�
�����K�8�P    JK�ϥZ�CC�)=L���+�~��Y�1!w    (o�   �B�8qB����'�q��*�u�Tl�޵.�S(�5zg�nl_Z�   ���.�]�#~�&����Y�Ν+�{���    �<p   �
p��q��i
z���al|k�cu�6+���{�Y�뻡����\^   �����=N��ӚJd��YM��ϟW.��Ν;    (?�   �����j||\ ~���PW$�p	��?�u�ڵ�g�)ݹ���\��~   �<9MC�^E�N.$������K�.�a�]��g�4    ��!�    e�p;�d������j}2K���1�˭����:=�L�m�C�����    *C���uA�.�5���!^ �e���B���|��^    �|p   �2T(t��QMOO�O�ꎅt;T�Z;��t�^�|:�P��_ڭ��\N    *��4��ƫ�ץ�I%s��������߿_    ��@�    ʌn�������q�!��������l���;Vg�t��   @�	��W��RF����]V��ڵk�9�_|Q    ��G�    ʈu!������� ���۩�h@Aw���#�6nz��A�   �n�a�-�Q����\R�<m���B�ׯ_�i�4�   @(���     ���v������ڭ���Z��(�v�.�����J�   �
�z�>�1��}9c�z����n�^x�    Jw    (���z��� �0�ӡ�j=.�����O�u�   �k��87r��|Ri�܁oY�>���k{>�o�>    Jw    (===�������=��,����6om����_O�   ���u;��.��xZS�� <b�ܯ^�*�ө]�v	    Pz�   @�����߿/ ��u:��̈́�hk��]H�������ו�l   �d����Z��V��BR� <r��e���;�~g5    ��*ϫ�    P%N�<���q��:�[ۣA;�Q����M[�~���Yݽ�n]�X|L�"   �g�:r5����TV 5����cB�    PZ�   @���?����!�.�i�+���l�]2��Y>����v�=�L
    ��5���4�tjp1E�;���/��r���C    ��@�    Jп��/
�w��=���r�*wm�w~�B��ᾛ�y�����   ���t;uw>��LN@����Ϟ=+�0���.    ��#�    %��O?�ݻw�ߜ��ma���^U���f�o��o�wt��9--.    ֒�ahW̯�DF�S���r7MS[�n    `cp   �b]H�����x]��S��m۱˾�����t��y-��    �S�߭�ǩ���♼�jf5�[�N�S---    l�    P"Ν;�[�n�� H��5xد͡�hm��r�y[���G�����   ��b-&�hl)��xZ@5��˝:uJ$�    ��;    ���/�ƍ����Ю��.�*M(�g~���q   @)0��5�Q��T�\R�|A@��B�O�֟��g566
    ���   ��t钮^�* �4<��0U"�   ���ˡ}u-�4��
�V�BAǏ�_��544    ���   ��ꫯ��p9Lm��    �N�PWا�ǩ���
+�����8�^__/    ��!�    �
�_�xѾXT�Z�S;�Br;L    6^��e7��'����FV�����_]�XL    ��A�    6��k���_�vFql��iK�O�a    P:|NS{c�/�5��a�>����o��p8,    ��#�    �l``@.\P�<�nm��pz    J���%�����'�)rG���r����[o��`0(    ���
2    ����}��'4��������i�    ���ǩꃺ3��\:'����y;vLo���<�     k��;    ����I�8q�p;���4�	�!��`    (7��nGԯ�匆S��M&�ё#G����Mn�[    ��A�    ���̌z{{U(T��ǩѠ|.�     �)����Jd��I*�ROO��z�-��L    k��;    ����e{�bkc�����W[�~    T��Ԟ�_��)M'��I<�C�    `�p   �5d5:���{�f�Ћ��r��*�u	    PY���Z�"��.$�+��sss:~��^}�U    Vw    X#�LF���r�Q�ǩu!yl�    �,�u���>�D��P=&''u��)<xP    ��C�    �@�P��Ç�H$T��W��C    �*�s��hh1��;١z����ܹs:p��     ���;    �������E��i����    �����������BJ����Ν;�x<��/)    ��#�    ����W>Pm�n�vՅ�u:    �^�>��.���J�
��͛7���={    x>�   `?~\�MSЫ��_�a     ���޺��Χ4��
�t+++�r��~����    xv�   `��={V������0��!�     �ɚ3n��4�p��bZ�����>���VKK�     φ�;    ��˗/�����thw}H~�C     ��F�[A�S}s	�������z��W���     ��#�    ��ƍ���/T���jn���     �9��}u�]H�a*'��
�8qBo�����     O��;    <����?^+l��*aRg$�MA�     x�⤲;���rF��8��J�����ӣ��zK�`P    �'G�    ���ȈΜ9C�U��rhg,����	    �g�p+P�c�%�)p^��q���ߖ��    ��pE    ���̌N�<io7T��ϥ��ݶ    ��q;�B}P�sI-dr*U:��|�����2MS    ��G�    �R"�бc��&�������'� �    X=�"�1�F�i�/�T*�|���~��!    ~w    x
�\N�V6�P����hPu~��    �k)���G~���)VVT���9�:uJ    �p   �'T(�p�ոT:�ˡ��!��    ���|���T�\R�|A@%Յ���/    ���   ���������J���[�    �^.����?��B&'�������F;w�    ��p   �'p��MLL�t�5>m���0�    ֟��zg̯�xZ�Ki�feeE�.]R Ж-[    �>�    �3�\����>��a�U�w    ��d-�����4uw!��ʊ�Jb�ܭB��^{Muuu    |w    �	w�ܱ�@%��]���     ����*�UM��%��T�B���Ǐ뭷޲��    �F�    ~���>���Q	�T1�[ݱ��<     �&�rh_]@�sI-dr*I.�ӱc����o��fW=    x��;    ����E����MJ@�j��ik�O�A�    P��E�;c~���_J�$�tZ===v��i�    p   ���d2z������T"�i�;T��f0    @y��fo	y�w�\H)ώ{� �x\'N��_��    �   �wX�����ݜT"�ˡ��5�9i    ��:�˞�ޞK*�g�=T���)}��z�W    Վ�;    ��#G�؍I@%�x]�Y���    e,�rh_]@�&��e>T���!�B!�߿_    P��   �7>��#����DMA�:#�     ({.���X@�I=HfT�k׮)���S    P��   @����5::*�uDjy    @%1�3��ij4�P	VVVt��9;�i�&   @5"�   ��Y�Hׯ_Pi����!E�.    P�Z�����̧TXYP	N�<���zK�PH    Pm�   �jccc�pႀJ�s:��!d�    P�b^�<1S�&�-rG�+
����?��9�D;    TfA    �V<׉'�m�JR�qiW]P.�)     �E���޺���Z����L&�cǎ�o��    ��p   P�r���9b��dSЫΈ_�a    �j�q���B�	ͥ9�򷸸�S�N����   �jA�   @U����L&T��Z_q�    @53iGԯ�xZ�Ki�nllLW�^����    Հ�;   ��s��	���
��Pw4�:�[     ��-!��NSC)VV������׮]SMM����    ���;   ��b5ݻwO@�p[[�ׇr3�    �5�\��η����|Y!��g�*+�
    *W�   T���!]�tI@��B�V��
�    �r;��.���J��ʕr�裏����]^�W    P��   �
sss:u�}��~��cA��     ���:L���7��b��;�W.�SOO��~�m�&�    *w    /����ѣ��x����=�A�    �'�4��uw!��dV@�Z^^�ɓ'�ꫯ
    *w    �P(�ȑ#J��*���_�5>    ��g���>���F�/B�����_|��^zI    Pi�   �h������;�|w,�z�G     ���=r���ZP�n߾�h4���N   @%!�   �b]�xQcccʝ������z��    �Z�.{�}g>��
1w����ϫ��V���   �J��q    ��ݻ�ꫯ�;��Ԟ��]    ���:�+�׭��rB�(?+++:~���~�m��~   @% �   �������������\�m���a
     ����8����Ä����r���u��1����ir	   @�#�   ���R)����P�b$�[��Ү���!     ���S�c��%��������_]    P��   �V������d2�Yc���Ѡ��     ��ihgį����R9����:{��~���	    �w    ���WKKK�Yk�O��~    ��g�#���BJS	JP~U__��۷    �w    ���˚��ٻ�/����㯻�]f�aeSDC�|�6mOlN�tM��&��6�Q������ *"3,�,�ܹ��&]�����<�|��0?���~���ʕ@7{tC_��   ���C����\�=�&�V+'N��ƍ�iӦ   t#�;  ��>����W�
t��:��M�X�	   ���UR.$ߞN������^�O~�T*�   t�;  �����s����C�F�R1On�@�+:   t�ͽ��|���������Di4���~���~:   ���9  е��f����m���Q�\ʁ-��W�   �i�ZΓ#}936�FS�N�h��=z4O=�T   ���  �Z�=�\&''ݨ^.��[S-��  �����v�>:��;]�ټys��   t�;  Е�z�\�r%Ѝ�+��<0�9   ��7�}mS;r���\3�-N�<�M�6�?   �@�  t��>�,��կ�h�֓'7�T,   �.��ڑ�ٱ�L���A��ʡC���3Ϥ\��   �ϛ  �U�����/��@��W��@��   нz�z�bco޿1���;�avv6?��O���O  ��	� ���l6�a�F��l�汑�h�  �����<9җnLelz6���!ǎ�w��   t2�;  �5�{�LLL�̓�����+n  �5����؆z>��|9%r�;�?>�6m��?  �N%p  ��[o��+W��͎�zv�   X{ڑ���zz��|>q7�N�<9��  �N$p  :�g�}�_��W�n�gC_�   X���\L>���Z�V:�g�y&�l  �<�T  ��6>>�_|q���E�P�c����   `}x���R�����}ˢ����������/��/  �4w  �c5�����?M��t�R�������^	   ��<�ۓr!���T$�t�۷o�رc��w�  �N"p  :�s�=����@�(�yrS�j=   ֧M�����|pc*MK�t����g���ٷo_   :��  �Ho��V�\��=�b��e0}=�    �ۆj9�o����ij��p���/�#��7  �� ��s�ҥ��W�
t��b!_�< n   ��P��'6����̩��`�V+�3�<�rYF  �>o&  @G���ɋ/�8�ݠ����^q;   �TJyrcoΌM�!r������СC����   �6�;  �Q����m�0�A��q{]�   ����o���c�����������5���o  `5	� ��q���ܸq#�j�RlH�,n   ~��_G���t��n|��lݺ5   �E�  t�O>�$�Νt��,����    ܋����FzszԒ;��^�O~�T*�   ��;  �ꦦ�r���Z��|���?�:�JI�   ܟ�w�'G���g暁N�h4r�����?�s   V��  Xu?��O�M�����r`��   X�z��'6����d���P7n�ȉ'��o;   +M�  ���_~9�n�
t�v��uq;   �ڑ��#�9=*r�s�;w.=�P�o�  ��$p  V�G}��?�8���+��<�q;   �D��v�ޗ3c�n���LG�ɏ���j�   ��;  �*����ꫯ��j:Y��[�S,   `)UK�<��7g�&3%r���������я~  ��"p  V\����~�����d���r�`J�v   `�T~��>:�I�;�֭[y�������  X	w  `Ž�����Ɇj=��恔
�v   `y�o�{b�/g�&31k����f۶mٹsg   ���  XQ|�A>��@'����M�v   `��G�{sF�N�:v�X�lْ���   ,'�;  �bnܸ��G�:�`��'-�   �������щL5��N�l6�����_��_  ���  ��h~<��s�?�ST�9�yP�   ��v���H_N���@w�ܙ1yꩧ  �\�  ��8x�`&''����oL�(n   VW�ȝv�<��Cٽ{w   ���  Xv�O�ΥK�����4����   @�hG�O����wrw��$���Z6oޜ���   ,5�;  �������o:UoO)_�:4h   �I*�K���K�w�,��9������?��O  ���  ��ir<����?��˥|}ˠ�   �X�R!Ol읏�g�������9v�X���  `)	� �es���LLL:Q��?��J�   �NV+�䦾�w}"�"w:����cǎ<��#  X*w  `Y�6.^��D�C�v�^�   ]�V*�ɑ��%w�;����m۶T*�   ,�;  �䦧�s�ȑ�Z��<���[���   @ש��ٿ�7g�&E�t���������~  �� p  �ܿ�����h:�|ܾup~�   �����#�3c�i���cccy���o|#   �%p  ��ɓ's�ƍ@��)���z�   �n��#�9�;��w�͎;222  ���  K����9u�T�������-�v   `��oG�zs���D�W��ʳ�>�b��  ��	� �%�l6���|�:I;n�������  ��e�R���#ro�.G���ɑ#G�W�W  X(�;  �$���LOO:I�Xȓ��W��   �M����G'"q�|��g��㏳gϞ   ,�~  `����\�|9�I��B��4���W_   `m���w���nM�a�����g۶m���  ��r�  ,ʝ;w��k�:;��l��   `=�T��\���ܲ��k6�9t�P~��  �~	� �E���~����@'yl�?�{�   XO��V2;��gw�Vۭ[��_�"��  ��!p  ��ѣ�}�v����З���   ���}�:�����L`��;w.;w�̖-[  p��  ��|���y������z��   ��=2XK��ʵ���jj�Zy饗��3Ϥ\��   ���  p�fgg��/:ɶ�Zv�   �d�p=s�dtZ���jO>|�p����.   �B�  ܷ������)��V�w��   ��;\�܍Vn�mV�_|��g�f���  �C�  �}9u���at���<6ҟB�    �K�P�c�9;6���ji�Zy뭷�cǎ���  ���  ��Ν;y��7�b�Z���k   ��J�B�Л�F'2�hVK��̡C����O  ���  ��g?���!t���R��y0���   ��)ybc;r���9��X=����#*��ַ  �� �{Ҿ>���ہNP�)������Y    ��J�8���̌ȝUt�̙�ݻ7���  �m�  �t�ƍ���ہN�>�������    ܻZ���7�sfl2�f+�Z:�g�y&   ���  ��~��ٴ���k/������   `A�zJٷ���c�Ѹ�Z�����������  �	� ����ѣ�����b��'6���    n�R�ޡz>�5�VK�������{��lݺ5   ���  ���]��s��:�c�2\�	    �7R��L��������_γ�>�bэ�  ��  �U�����-8�vo�͖�j    X:��*�;�̕���j�����E����n   ~C�  �V�����&V�C�l�   ���s���f+קf��O>ɥK��}��   �	� ���}�p��j��[����    �|��2;�ʭ�F`5���y��gS.�X   �;  �4�ͼ��K��6T-��
   `�<����c������F��W^y%����   p  ���fff&����R��<���   `E���<ގ�G'sw�Xi��y>����ٳ'  ��&p  �Ӆr�ҥ�j���9�e`�P   ��S-�#r�L��
��'Ndǎ�T*  �/�;  0ovv6G�	��R���mH�\
    +�����6����T�-�;+��h��_�?��?  X��  ���~>r��R($OlHū*   �j���g��oNV���hΝ;�}��  X�T  ��a�իW�����P�	    �oS�'�s�|6~7��Z�VN�<�;v���7  ��#p �unzz:���Z`5�����    �9��W3;���ə�Jj6�y�����0  ��#p �u��K����v���`=    t�]C��4�����u��ͼ��9p�@  ��E�  ��ٳg3::X-j=ytc    �\���щL��VҩS��gϞ���  X?�  �N����7���ޞR�o�O!    t�b!y|co޽>���f`�4��>|8?��  �w  X�<�Fõ¬��b!OnH�X    ��R,���9=:��V+�Rnܸ�s��e߾}  ��;  �C}�Q�^�X�B�����{J   �{���g��nLVJ���ɓ'�k׮T*�   k��  ֙���ǎ����2T�:
   ЍFj=�1��g�w+��]��������   k��   ֙�fvv6�vֳ��    ����j��\�򝑕s�ڵ\�pa~�  X��  ��\�t)�/_����Jv�   ��g���F3wf�+���_ώ;R.�]  `-�?  ���µ�jVZ���#�   `m(�}�yot"w�|sde4�9r$�7  `�� �:��K/��ݻ��V)��恔ڧ�    ���>�7���щ�5E�-���J�o�  `m� �:p�ڵ|��'���n��q{�T    kO�\�c������cǎ��g�M��#  �Ew  X��f:�V˂+ﱑ�T�z   �e��r���Ӂ�0333���_�e  ��Ge   k\�#���$V�#C�l�   �����J��|19X	/^̾}��u��   k��  ְ���|�ᇁ�����G�z   ���k����\n��V�+���g�y&�b1  ��!p �5�^H�����J)���   ���PH�m��{��j�.��{�nN�<�o��  ��;  �Qo��F���+�Z*�k�Sj�f   ����Pϻ��i���>Ⱦ}�2<<  `m� ���O�>XI�B!OlH��:`   ���^.���z>�9�VK���j�����K��  `m� ����ϧ�t0+kT�f   �l���P_%���,����������/  @�S  �s�ԩܼy3�����j    �7��W2٘��t#��ڷ��۷/}}}  ���  ֐������[��4X-g�po    ��3T�Tc�Ǎ�,�V���_~9?��  t7�;  �!/��b���+�R*f����    ��V*��p=��&�h���ƍ��㏳gϞ   �K�  k��˗���VJ;j����TK�    ��R/��?�9=��˥��u�ĉ�ڵ+Ţ�  Э�  �F���+�XQ{7�e��   �?lC����*�t�n`95�?~<O=�T  ��D  �5��^���d`�<8P˶�    �W��+�l�el�XN/^�O<����   �G�  ]nbb"gϞ���j9{6�    �מ�Z��_=��ri�v�ꫯ�駟  �}�  ��<�f�a+�R*�̓)
   ��U*��p=��&�h��e||<gΜ�_r  ���  ��G}�����JhG�_�<�j�    X�z��݃�|xkz~i��/���ݻ7�J%  @�� @�j��;v�+fT�F   �xk�<����;3�����~�ȑ����m  ��L  �.��+�dvv6��e�@-    �T��U21;��w���ʕ+�϶m�  t�;  t�7n����0T��ލ�   ��T(�w���F'3=�,��G���g�  ��  Ѕ^xᅴZ��r���yb�@
�    ��+ylC=�G'3�'�dzz:o��f���o  �|w  �2��Nn߾Xn��}#��;    ,��r1;����t`��={6���O___  ��&p �.2;;;�2+ᑡz6�+   �嶹ޓ�ٹ\��,�������J����  �lw  �"����\`�m�U��Po    `���eb����(�ctt4/^�Ν;  t.�;  t�+W����ˁ�V)����    �J*�G��ywt"s�V`9����y��S,  t&�;  t��^z)��
_=�7�G�    ��j�Bv���ͩ�r���������SO  �Lw  ��E��):,�]�2\�	    ���Z9��=�bj6�.\��dxx8  @�� @�k��gΜ	,������    V�ΡZ�4����,�#G��G?�Q  ��#p ���K/��l�S�\��    ������p=�Nd��
,�۷o��?Ξ={  t�;  t��W��ʕ+��T($�7��X    t�j��=C��c2��Z�VN�<�]�v�X,  �w  �`/��r`���П���C    :�p��m}�\��	,����������v  �Ρ`  �u���ܹs'��6�V��@-    Щ����\�g�K�>ȁ���  �3� �5����XN�r1�F    ���ճw��wG'�h�K��j��ѣ�����   �A�  �W^���l`���Sj�    �Z*���ZΎM�ڵk�r���<��  V��  :���xΟ?XN{7����   ��1T)硾J.O��R{��رc��O~  `��  �ü����a�l�f[-    �m�Ts{f.�s��499�w�}7  ���  �A.\������ri_���H    ��z�P�;�'�h
ai������\��  �j�9  t����\
�B�4�r�    �V�b!�����t`)5�?~<���w  ��;  t�7�x#��dX>��3\�	    t��ZOn�����l`)}�駹u�V���  ��;  t�����9s&�\�j=yd�7    �V�����\���Ri�Z9r�H~��  Xw  � /��b���ˡ\,f���    �ZR,${��9=6�f�X*�����g���  V��  Vٵk�����ˣ�R-    kM_O1��+�t�n`��W�O�8��;w�X�m  V��  V��Ç�?��r��_˖�j    `���ۓ[w�5�L����l�z��ɟ�I  ��%p �U��{�e||<��=����    X�
�B�������6���tΝ;����V��  �J� �*i6�y��7ˡPH�����    ָ�b!{�jy��T`����9r$�w  `�� `�=zt��SX���2P��   ��1\-�ޞ\��ݕ�s���\�~=�6m
  �2�  �
�����G���z%��   ����Zn��e��,��Ǐ�G?�Q  ��!p �U���/�_m
K��T̾��    �zT��yt���F'3�j���۷s����ܹ3  ��� �
�y�f._�X�R*    ֫z���*�p�n`)�Z��<yR�  +D�  +쥗^
,�����+   ��nko%�f�26�,�������{��׾  `y	� `]�t)ccc����Sʮ��     �a�`-�3�m�K�ԩSy�'R,�E  ���  V�ѣGK��ճo�?�B!    �(�5X�7�Kann.���/�g�g  ���  V�ٳgs�Ν�R{x�7�՞     ���Z9��z�O7Kᣏ>�7���j�   �C�  +��lί��R믔��`=    �o�s���ىܝk������^�_��_  Xw  X'N����L`)�<>�?�    ����Bv�r��T`)\�t)7o����p  ��'p �e��Ϟ=Xj��{�W�Z    �P����=�br6��?����  ��  �ّ#G277XJ��r��    ܛ���uw.�s��b�����իy��  ,-�;  ,�;w��O>	,�R���7    �w�B!{�j9=6X
�����  ���  ���Ç�j�Ki�p_��b    ��3P)塾J.O�kbb"~�a}��   KG�  ��ڵk��/KiC�'�j    f{57g��m��7�̞={R,% ��"p �er�ȑ�R*�ٷi     ��
�ޡz��H��,���lN�:�o~�  ���  ���r�֭�Rڻ�/Ւ     X�z�8�������b�>}:H�,� ���?k  XǏO�e��������}�     Kc[oOn�m���\`1��f^��<��S  O�  K������T`����ytc_    ��S(�g��S�'ҴW�"]�x1������   �#p �%�^ii����R*    XZ�R1��r��t`1ڷ����k����  `q�  ���|������ʖ�jF�     �ckoOF�gs{f.�W�\���x  ,��  �H{��̙3���S*fφ�     �k�P=�\�H��
,T{���������   'p �%���[ogI��ЗJ�    `y�J�l����Ÿv�Zn޼����   #p �%�h4r�ܹ�R�W���    `el�dt���ٹ�b�Wܿ���  X�;  ,�cǎenΡK�T,�ё�     +��ճg��wG'�jlttt�	  p��  �H333���Keφ�TK�     +��\̃��\��	,F{���?�a  ��'p �E:r�H��f`)�z���    `ul�f�n#S�}Y��7o�/��֭[  ��;  ,���T>����R(
ylc    ��S���3T�{����x�����O  �?w  X�W_}�z;Kf�po�=�     �����m}�\��	,���x.]���۷  �ww  X�;w�����0P-g�`=    @g��_ɍ�F�猜�p'N�� �}� ����+��Y�B!�F    t�R��]C՜�
,���d>����ٳ'  ��� �ܾ};��y
�B`�����    ��U���ۓk������/)p �� p �x��K��RΎ�z    ���p57��ef΍�,���tΝ;�}��  ���  p��_��/��"�X� �؟��     �c������܍��B����w  �Gw  �O���j`)<4P�`�k    t��rFj=��,���LΞ=����  ���  p�����Ū���9�    �;����L#�f+��N��_q/�  ~7�;  ܇#G���rx��=:ҟR�    �;���_���w1;;�w�}7�G  �w� �=���Os����bm�W2��    t����\�j���\`!Μ9�Xq ��C�  ����_,V{�}�H    ��S(�k��wG'�h4�� � p �{����֭[���9ܛj�2    t���b�������B�>}ڊ;  �w  ����Z`��zJyh�    ��=�_͍�Ff����������  ���  �\�v-7n�,֣#�)    t�R���k���T`!�  �	� �8v�XZ-+<,ζ�Z��=    ֆM�r���rkf.p�fggs����߿?  ��$p ������,FO��]C�    ֖]C��s�N�6RX�w�yG�  ���  ~��G�Zog�vo�OO�    `m��
y���Kw�����LΝ;�}��  �/w  �n޼�/��2�C��<�_    �6=�_���l����j��� �� ���ꫯ�������     kW�;�#ռc*p��������G  ��  �[����/�,Ǝ�����    �m��rFj�N7��ԩSw  �o�  �[���[�V`�j�b�    Xv�rkf"��o�ܟ����?>�w�   p ��cbb"��y`1�n�O�X    �>���_���Ӂ����o� ���  �9r�z;�2R��?    ���@oO������\�~��w>���ر#  ��	� �i_z����B����    `}�9P�����:y��  "p ����W_��΢l��^.    X�*�l��s}����+W�d۶m ��L�  �6===�',T�T�Ã�     ���Ռ�m�iO��t�ĉ�˿�K  `=� ��;v,�f3�P�7��T,    X��c�U�ٝ����իW��  �+�;  |eff&/^,�`���}�     �=�_͗S���3�����/~���� ��J�  _9~���v�P(d���     �F��Ǉk���T�~ܾ};_~�e6o�  X��  �{�����z������+    ��X-g�����F�^�Z������ ��H� ��w�ĉ����T,d�Po     ~�G��5�H��g7n����x  �� �u�ܹs��j��R1     �M�\��z%W'g����������  Xo�  �k��^ff*�0�=�<4P    �ﳽ���ӳi4͸s�^�:�Q�T  �� �u���,Ԟ})    �{�����������j����������  �z"p `ݺp�B&''1R�dc�j    po��˹6U��l3p��g�g�b�  X/�  �['O�,D�PȞ�}    �W�B!;k9=jx�{�l6��;����F  `�� �.]�~=7o�,���z��R     ��@O)#�rF��{u��Y�;  �� �u���ぅ�)��`=     ��@57�6�l�I��ȇ~�G}4  �� Xw&''s�ڵ�B��؟R�    �����y���Kw���;�#p `�� ��=z4��i�_��-��     ,ƃ}�|19�Y3�ܣ�x��˗��C  �:�;  ����l>���B��M�`�    X��%�;�9k:p��z�-�;  �� �u�7������Sg~��_��g8
IX>���wk�)W���S�����ڿ|�U�hW�lY�@� 3�l�ȑ% �������K��t�G�;��n�i]��.    ��p�V���vl�{f�ɼx�"���brr2  `�	� ȍ,l���	8�l�=[o    8K��VㇵV�I]�~=����=  `�	� ȍ�7o���^�i]��c���	    8[�B������ĳg�bgg'��j  ��Rh  ��}�]�i�Iį&    p>��w��������;�����o�  0��  �������	��ǣ���     8�R!.U
�|g?�$?~�n7�Գk  ��� �\�������*��d�     ���F+���6�9�l���o��/��2  `	� z������pZ��ע�&    p�*�4>���ik/�$��k����ي;  CI� ���ӟ�pZ�b!��T    �"|4R�������q�x���q�������  ��� �����+++����z���v    �bd�I~8R�ٍ����s�� ��$p `����G�z�n8��J)��+    p��k�Xj����g{{;���bzz:  `�� Z�n7fggN���     �h٩��Vbf};�8��ύ7��c  �0� 0�n޼�N'�4.��1^-    ��p�Z���B4�<��x+++�����SI w  �֝;wN#������    �ٯF+q{�pׯ_����:  `X� JO�<�V��N��h-�%�I    ��5Z.�d�k���y��qt��H�4  `(7  J��N#M">�    @?�d���N�z����t:q�������  ��� ���-������G��(��     ��^�V���cŝ�ݾ}[� ��� 0t���?Y��T
i�Yo    ��ߍVbmg?<��8;;;������  �N� �P�v���ѣ����z;    Ї��4.�J����6��ύ7��c  ��� 0Tn޼�N'ऊi�V    �}<R��;��ur)�XYY���ݨT*  �L� �P�s�N�i|2V���v    �OU
i\�c�eŝ�]�~=����  �A&p `h,,,D��
8�,l�h�     �죑J,o[q�x�?�n�ij� ��%p `h���g�i|:^�B�    @?+�IL�K��x�N�w�ލ�?�<  `P	� 
�r���J�Ie��^�    � ��Q�g���Xq��o�� 0��  �?��O��P�S�t���v    `@�$>h��ɖw�ngg'���bzz:  `	� x�n7=zpR�z�t�z;    0X>l�c���]�/-�q�F��  Dw  �_����t:'��Ɇ�v    `��$�5�1���6+++������  �� ��w��퀓��
q�z;    0���˱�lǞw�q������  �� ������V+���D#     U�D|8R�ٍ���y��q  � � 0в��^�J'3Z.��z9     �t�t�������������>  $w  ���~,--�ԯ&�    0�V��x���6�o�� 0p�  �o��6�]�4�L��~�f�    Wk�Xh�Yq�^�x�f3�F  ��� 0��ݻpR�Zo    �H�D\k��w�q�ƍ��o  �� ��������'�(b�z;    0dVܷ�����277  0H�  ��ׯG��='�	G�    �'�V�G*1��p�N���ߏ�>�,  `� 8�v;���N�^*�T�     �h�V����س��[ܾ}[� ��� 0p����;��n�I��x-�$	    �a����(���n�Q^�x�f3'� ���  �{���D�X���J     �j�x�lǾw��ƍ��7�  �;�;  eqq1���N�Ӊz�n    �]!M�z)��G���  w  ���ף׳@���4���    ������9B�Ӊ����g�}  ���  �v�KKK'�w��H��    @>�w��Iӊ;G�}��� ��'p ``ܸq#��n�q*�4��     ȓ�x�jG׈;Gx��E4��h4  �J� �����	8�O�k��   ��)�IL�J�p�lP�o�	  �Ww  ���b�Z���d/p��T     �>����~t{f�9���\  @?� 0�_�p��׭�    ����\��b��8L�Ӊ����g�}  Џ�  ��v�KKK��^�|h�    ȹk�R,��aÝ�ܾ}[� @�� ��nܸ�n7�8�ף�Zo    �RH�J��Z{���؈f��F#  ��� �{333�)�I|d�    ��G�J,����s�^�w00��7�  ��;  }�ٳg���p�Gk��    �W���T�+�V�9ܓ'O  ��� ���������$I�[o    xՇ����#������\|��'  �D� @��v����p��F%*�4     �?�b��b�h�����w  ��� ��u����t:��d�     ��Ñr�X�s�������45" @�� з��8ΥZ)�B     ��r!�B4���^�w�܉/��"  �_� �K�v;�����w���    ��Z�3�������  ��;  }��o�=X��-c�R
     �6U)�\!�ݎ��l\�F#  �� �K���8�'�     ��$�F%f7v��%��_�5  �� �;ϟ?�V��6�b!��+    ��֊1��D������w  ��� �����瓱j     p2�$��z)�������ӧO�ڵk  �� ����ɓ��)�IL7�     �q�Q��V;�F�9ĭ[��  ��;  }eff�`%�棱Z�$     8�l<�r��Z�������v���i  ��$p ��d� �6�1��Xo    x���X�ޏ^ό;?���w�ލ�?�<  �}� �7��v������H%J�1     �VLc�\������	� �w  ��_���1���Z     ��>l��jss3Z�V���  ��E� @߸w�^��\iT�V*     �n�\���][�N����׿�W_}  �� �kkk����6��    �Ƶz9^���c�;  �� �������h�c�0     g�R��B��n��vwwcii)���  �u  }a~~>�m>�     g#I"��J1���[�n	� xo�  �w>�v�p�R!�+�;    �Y����Is7����y��Yt��H�4  �	� x����p�i     ��b�ĥj)V��^��t�>��  ��&p ���?�8JvL���     ��Z�,p�Pw��� �^� x�~��ǃ8ʕz%*G�    ��F1��r!6۞��s���CEi�=  K� �{������G��     ��L�Jw������~���  \$�;  �M�����p��r1�*n[     ��T�s[���t^u��=�;  N) �{s�Ν��8�G��     �|%I��Z���j}}=����X� pq|� ����R*�q�!p    ���R<i�F�.����|��  E� �{��}����Ñj�I     p�i���X��x�����  \(�;  ��_�������p��k�6j�    �"]k��ass3��v���  �� p མ��	8��z%*�4     �8�b��Bl�;/e�E�oߎ��
  �w  .\����ŋ��|4f�    �}�����ѣGw  .�� �w��̓�8�H��R     p�j���j�n��R�ٌ����V�  p��  \���Z     �~$���K1���R6\t�֭���/  Λ� ��j�bcc#�0�4���r     ��\��b~k7�ʫfgg�  \�;  ��͛G�n���$    ��SJ��,cuw?ढ़����܌���  ��$p �B=|�0�(�Fk    �����yU�׋۷o�W_}  p��  \�lգ�jf�Z�F�     ���BTi�t�/���	� 8ww  .̍7�=�0�F�    @��R+��V;ढ़��X__����  ��"p ��<~�8�0�4���r     �?���1�l��^u�֭��o  ΋� ����������Q�B�     ���&1Y.���~�K  �I� ���y�f�Q��V    ��3�(�������a����  �� p �B<y�$�0�R�K�     ����Q-����dz�^ܾ};����  �� p ��mmmE��
8̵��     ��J�s[퀗�>}  p^�  �����/�)�iL��    @��Z/�|��^�����������  ��&p ������F%
I     ��R��d����/ݹs'��_�%  �	� 8WقG��8̵�j     ���e�;?3??/p �\� 8W�n݊�3K9�D��R!     ���BTi�t��V�u0tT�� �l	� 8W>8̵�    ɕZ1���l��~�?��  gI� ����ߏ����ו�$.�+    ��Z/�|�n�G�	� 8sw  �͝;w��uT)o�nT#M    ����L���������<<*%H  ��. 87���8���v    �At�^��3?��c����}  �Y� p.�������׍��     �g�R<Xr���2<� p�T%  ��l�=���u�T    �����\+��f; ���~�N(M�  �� p �\d�Q��W�     `p]��^�w������&  �,� 8Ϟ=x�T�|pt-     ��^L�־�\�333w  Ό� �37;;�N'�u�#�     `�e+�����  ��"p ��ݹs'�u�4�K�R     0�.�J�xk7z���᣹����O  ~)�;  gnqq1�uӍj�I     �R��D�k����w�
� 8w  ����R����n�Q	     �ǕZI��O�={  p�  ��[�n��^*�h��    �0����&���t:��!����  �_Ba ��ZXXx�#�     `��IS�b,m;ٕ���?� ���  ��f�;;;�J�$�6*    ��R+	��ɳg�  ~)�;  g��x�D��B     ��r!��4Z�݀l��jE�^  xWw  ���Ǐ^��H5     ^�k�x����w�^��?�c  ��� p&��n������&q�^     ����We�Hw  ~	�;  g������^u�^�4I    ��UN���c}w?�ŋ�Hi�  ��;  g";n^7=R	     �_��.p'�"���ŧ�~  �.�  ������WU�i�WJ    ��"M"�{�o�߿/p ��	� �����boo/�UW���    �$1Y)��+�D,//  �+�;  ���۷���W]i�    ��r�$p�@�ݎ���  8-�;  ����|���B���n     ��x��4���Q"~�����/  NKq �/��v8�UW��    �N�$1Y)���^��'O�  ��;  ��ݻw�׳���	�    ��r�$p������PR��  �!p ����	x�h��b!     ȟ�r!Ji{]�8y�$=z�(~��_  ��� �_dyy9�UW���    ��R�K-+�Dܿ_� ��	� xg+++�����;    @�MUKw<�<  ��  ����.�U�RT
i     �_c������N7ȷ���X[[����  ��� ��^u�z;     s�R��-�;w�ލ���*  ��  ��v��f3�$I�J�     p�V���� �I  ��� �w����G��xi�R�r!     h�
Q-$���.!�Z�V���G�(S �d|s ��<x� �UW�     �����x�l��&�������  ��� �NVWW^J����;     ��r�(p����� �� pjϟ?�N��ҥj9Ji     �R�X�z��=��nmm-  ��  �������    8�TE�N���^lmm���H  �q�  ����B�Ki��T�     �Z9��333�?�!  �8w  N������F�K�b�$     �u�B�b��n�oO�<� p"w  Ne~~� r����+     G���e�=�^�x  pw  N�޽{�ʎ�    ��\���=�:�N<�<���  �F� ��,--�4^-E��     �Q*D���n�	�y�)	� 8�� ��v��l6^�R�     �R�O�V��nqq1  �8w  N,[���z/M��     Ǚ�܉���:TJS�� p4�;  '������F+Ũ=�    �x��4Ji{]C:y�)-,,��  p�;  '�����e��     �P�$q�Z��������  ��� ����9����J     �IMV
��
rnyy9  �m�  ��ݻw���L��F�T     8��r1
I�r��j���~��%  �"  '2;;�ҕF5     �4�$b�R��;�A�=|�0~���  F� ������4U+     ��T�$p�`XI� �Q�  kcc#���2�Bc�;     �7Q)F�Dt{A�=�<  �(w  �����G��I3��r�     �.��}�\��]+�y�+���D�Z  x�� �c����t�^	     xW��{�e�J333��_  �N� ��^�x�)�i�WJ     �j�Z�d#�ٱ��,	� 8�� ��Z\\�N�����"I     �Y)Mb�\����y���  p�;  o�	/M�+     ��d�(pϹl`��lF��  x�� ����!��g��    �/5Q)��f�c�^/�߿���  �*u
  o���������     �T�X�j!��N7ȯ���;  o� p��������L��     ge�R����=ϲwQ  �:�;  G�w�^�Kw     ��d�K�� ������nG��  �G� ���<y��Ҩ�
     ge�\�B�D�����Ç���.  �%�;  GZ[[�L�+     g)M�-b}w?ȯ��9�;  ?#p �P�V��XH�\��     ��d�(p�9�K  �N� ���ݻ�I�����    ��7^.�����n7�4  �� 8���|@f�Z�B�     ��j1�Z���� �z�^<~�8~��_  d�  �����K�r     �y�(������� ��;  o��ۋ����̥Z)     ༌��x����J  �Kw  �p����L�T88     ��d��ͽ����|��ގn�i�  � xCv$d�j�     ��$��������bqq1>���   �;  oX^^�L�J     �m���	r�ѣGw  � ������H($I�W�     ���#��_nF�P��   /	� ����كc ![oO��    p�j�R$흿������V  @F� ��<|�0 s�V     �(#�$��^$�Wr);e����155  �� ��YZZ
�LV�     \��F�Zތ��� �<x p @� ��5�̀Z��b     pQ��5��pA��c��  �� �������0Q+     \�4Ib�T���ݨT*A�lnn  � �Iv�#d&+w     .��1��E\�z5ȟ�����ىj�  �� ��<{�, I���
�    �xY�~s�iLMME�P�gvv6~���  �%p �'/^�)�TH     .�d��b!677cbb"ȟ���; @�	� 8�����`�    ��%;etz|$��������Z  �ow  <z�( #p    �}�6>�W�c{{;j�Z�/��;  �&p ����\@�$1^�    ��d��{u�݃����   ��  X^^���&     ��h�#�r4���t:Q(�|���� �� �[[[U��     �L�������܌��� _�={  �� ��P`R�    @�9�766�9���  �� �x��a�z� �
I��;     �_�����ۋ����jA~���F�ۍ4M ��� �����R$     �_�T��F-֚�+���y��i|��G @�� ���Հ���v     �����A��l6���D�P�cnnN� �Sw  ��jL
�    �#�&F㇅���z���A~���  �$p ȹgϞE���RH�^r{     @��:6i�D�׋���{�lmm  ��` ȹ��ـ	��     ��b!���z,o4coo/����V��������(�� @�� rnqq1`�"p    ��d+�Y���V����5����  �E� �skkk�    �GW�?���lF�ӉB�����  ��  9��vcww7ȷb�D��     ��+��H�$z������A>���  �#p ȱ�X��a0�6^)�     �~S.b�^�������i�Z @�� rl~~>`�Z
     �WW�?�{{{����j5~�i��j���h  �w �{��Y�X�m     ���X#~|����Y�,pϏ�D�/��"  �% @�e�ɷB��H�m     ������~��ڊ˗/G�$��3� �?J ��ʎt̎�$�F+�H�      ���ʥ�Vbsg����G�ٌ���`����  �"p ȩ'O�D���m�Z
     �wW�?��Z�{>���  �"p ȩ,p���[     ��ձF<x���ϭV+:�N
�`�e��Y�^�V �|P�  ����r�o�߮��w     �ߕ�7�ڳ����`�e'����o~�   �  9�����h��4	     �wc�J�ʥ�n�����=?�  9"p ȩ��N�m��v     ��qe������s�ݎ��ݨT*�p[[[  �C� �C����9�o�R     ���2���=���܇_��  �C� �Csssc�;     �cz|�ϲ�}jj*�$	����^t��H�4  ~w �Z\\�^*D)��    ��1Q�F�X��~�ϲ��jE������R\�v-  ~w �Z__�m�j�    �����_m�����>�V���o~~^� �w �j6�A����
     0x.���ܳ��N'
�B0�VWW �|P�  ������C^�m�b�    ���-�fkk+��ǃᵱ�  ��  gfgg����UL���     �A35R?����M������  �A� �3O�>�m�\�$I     M�X��Z%6�;g�s�ݎr��l�i}}=&&& ��&p ș�ϟ�6Z)     �K#�7�L��>55���y�; @� rfkk+ȷ���      ���z<Z^{�����}�-//  �O� �#�n��xN�m��6     ��55R?�������ىj��/^  �O� �#O�<�^��W��F��     �K#�H�$�����V��ë�j  �O� �#Y�N��VJ     �,��'�x��f��/_�S�ӱ� �w �YYY	�m��     ��wy�~h������Q�Ղᴰ����� ��n ȑ��� ��*n     |S������d+��ᵼ�,p r� �Ɏl$�FJn     |S#�#��/_�$I�ᳶ�  7u @N�������k�\�B�a>     �o�V�r������v��j���h�'�  7�; @N<}�4ȷъ��     �l����桿�"h��p���  ���  '�|-��    ��x[��l6���E�8�t�d�����r9  N
 ��X]]�m�R
     S��#���Y�>22������O ��$p ����moIz���|�dI����K���Z ȓY�=c�߻�lk3�̮mI�DuU� �)e��BT������A��� �:      ?\�}������� �M� P��b��b2��    ���hg�qܯ7_����H۶QUU��_�5  ȗ� � ���v��u>��    ���?�}3p���qA^�u~  �r (�O?���|�?     ��>��~���w!��=?��2  ȗ� � w�Fu     @n���{�E4Mu�<'���ݫ��   ?w �|��1(W5�\�    @���揾���>޽{�c��?<�ۿ�[  ��; @>����ۻ�     rs6�d4��v������	�3���?� 2%p (�r��uf�    ��]�g��͗o�{���mۨ�*ȇ� �%p �\w`�^��r�O|�     _Wg������������˗   OJ ��Y��|�k?     �z6{�=���V�   OJ �����wP��Q     ���'��"��}� ����&㪪 ��� 2g��l���Q�`    �|]ΦQ����|O�w����Y��O�>ŏ?�  �E� ��ϟ?庘�     rVU���O����w�w/p��_��W�; @��  ��k)���     ����ٓ�n�}0y�� ȏ�  s��:(��H�    @���G�Ӷm�V���/i���	  �#p ������	庘�     r���i�z��D����  ȏ�  c��_�r�*&u     ����E������?y�n� @~�  ���cP��q     P�Q]��tw��w��4����t:���d���b8�@ �ķ; ��}��9(����}     �q=�=�w�w�{�������  �x �ؗ/_�r	�    (���,��G���>|� p ȏ�  c��"(�|X     ��j>{����ml6���A�nn��  �"p �Xw8K��#�;     �x7�<��݊��=n4 ȏ�  S���~��4�QW�     �R\L'QU�h�ǟ�t����u�>7 �G� ���~�I�^�ٰ
     (I��O�q�\?���z��.�C�L��h ��� 2���?�:��    @y.��'�n����2H[�4ѶmT�� �\�^  2�믿��     �Ҽ�M��?o����b!p�D�\�Ç @�  �����5�    (��|���.�����1��}��Q� ��; @����5��    @y�=#p���.r���A�~��   � �L���L�j��    �Ҽ�Mٻx�)����p�1 @^�  j�6��	�t6�5    �2�*�&��[m��~7���� �� @�>~���e�3�     �z7�>9p��v��lb<�r�1 @^�  ��矃r�-�    P���4�߯�O~��-pO[��
  �C� ��_~�%(�|T     ��r6y�������*HWw����]���  �� d����A��F��    P�w��޿\.�mۨ*2)�n8� �A� ������Lê�q�     �r]�=/p�t+���}��)��?�#  H��  C��*(�|$n    �l����x����?#pO���M  ��; @��ۧؒ�����     p9�>;p'm>C �|�_  2ӭ�����L�Q     P���$~�����o�&��uL&� M�� @�  ����SP���     �b6}��t��tm6�   w �����A�f�*     �t�����>����4u+�  �A� ������\ӡw     ��=�}�^?D�u�=U�
�|>  �&p ����]P�I]E5     ��l2��`���Y?��A�����  �� dF�^��Ȣ     t�A��x��ͳ~n�\
��������  �M� ���j�i6�    �o.��g�݂;麽�  �'p ��f�Z�1V     ���lq�i���Y�x<��c �<� 2���2M-�    ��:��/�K�{�,� �A� ���j��>(�l$p    ��\L'�\I_^^�q�1 @�  ��_�r�,�    ��:��w�ݠ�`0Ҳ�n ��	� 2"p/װ���r�     ������.n_��1�N��4M  �O� ��ϟ?e���      ��hX��o�����s��.pO�b���|  �K� ������L�Z�     ��|6���ų��������t7� �&p �Hw�J�f�:     �?��N����z���m��̤�������� �t	� 2�]�I��#�;     �����������Z�,�'�˗/ @��  �l6A�,�    �?��M��nXH������   mw ��4M�if�     ������}�Xć����  }w �Lt�d�m��b\     ��������n��ƅ���LJ��u  �6�; @&>~��i:�b0�    �?��GQWU4�uk����A:��m  �6�; @&>��iRW     |��d���V���q�1 @��  �����4
�    �[f����b�e���f���x  �I� ������L��     ����C��n��6F�Q�������� �4	� 2�Z��2Yp    �o����ӗ˥�=1���w ��	� 2��R��Ђ;     |���nd�ݻwA:�E  �.�; @&6�MP�qm�     �e>9~������  �� db��e��    �������n��e6��� �6߼ 2��R�z0�a5     ���&��j����� �� @��  �h�6(�dX     �m�aú�]s����r)pO�z�  �%p �@w�����L�U      �7��vyx�l<-n> H��  777A�Ƶ�     s6�o6�h�&��ͪ)� �M� ����۠L�;     <j6�;��u�����?F   ]w ����e�    ������r)pO�~���m��<G H��  �rM�f    �1g��ѿc�Z鸿�����   =w �,��L�a     �����/����e��`�����  Qw �X)פ��     �����{�w�df�Y�_�|	  �$p Ȁ��L�`ue%     s69~��#pO���]  �&�; @v�]P���z;     <Ũ�^ۦ9��,�˸���o�X  i� d`����w     x��x��q��[u�� H��  m���    ��M�]&�>�w���X��1�L�~�>'  �$p H\���4�     <�t�2��r��'��  �� $���&(Ӹ�     x���e2��j��v�  �$p H���]P&�     �t/��^���s2 @��  �[,A���*     ����F/�{v���k8�����  ]�i $�5���     O�R�n�]��o��>  H�o�  ���k\�     <�K��󙳳���,� ��78 ��	��e�     ���鿻�����
  �"p H��2ՃA�w     x��^p�����  Aw ��	��4���     ���0�jm�?�w����l61����  i� $�;<�<�     �y&�a,7��]����ߺw  �#p H�v�2���eTYp    �皎^.p���/..���� �&�; @⚦	�3V     <O���t�u+�  �G� ���n�gT	�    �&/�o6�h�6*g���}F  �G� ������k��     �\/������t���  Mw ��5M�gT     x���W����Ƕ�m  ��; @�,��iT�    �^:p_��A�v�   =w ���V�\�     �y&���N	� �$p H�b��T,�    �s��/; ��M�Dm����  i� $���>(Ө�    �s�^!D�V���΂�i�6  H��  a��2(�`0�Z�     �6�|*�^��=��� ��� �X,����     p�q]����w�ɂ; @��  	��^�Z�     뇛R_r�[��o��&��q  ��; @�V�UP�a���2     P�Q]�f׼��k���U�u�?�`��  -w ��u��gX�p    �C�������l6������  �!p H�n��c�     7z����z-p�)�Q  �� $L�^�ڀ;     �[pi]�N?m��   -w ���m�gd�     6~�w+��� H��  a��44�     �^'p���18���  �� $�i��<u�p     5z��N�O&��_F �G� ���m��*     �Ì�����k�{Yp H��  a'�Tp    ����;�#p H��  a��4��     {�w��` @z�  	��iX�p    �C�ւ�����  �� $L�^&�     p��+-�����n�1���h�&  H��  a�A)��     ��R���V���"p H��  a�2��    �p�+ޔ��l�~� �G� �0�{y�AT�;     jT�^��-��/w ���  !��    �8��Ҷm  ��; @���8���     �y��}��=,��u��  =w �D��L��     �RW��6$��n�=���  i� $j�Z���     p�nPf�J��f���t�w ��� ��R�     p���b�J�g8�"p H��  QG�T�p    ���A�_�wo��   'p H���LU      Ǫ��;q��_��}  ��; @������     G{��}��E۶QUfk���,  H��  Q��(�w     8ְ~���*�L&  <��  Q�&�$p    ��_y]}���{b��
 @r�  ����Ay*g�     p���;��� @z�  �j�&(Ome     �&p ��� @B*�;     �~�+S��m   �� $ʂ{�*};     m���]���c`��ڶ��?s  ^��  Qݡ(��     ǫO�(�E��$x{w ��� %p/Sm�     �Vׯ;o6�{Ot�;  �� $�i��<�    �x��4�;�`8
  -w �D9�+��     �w�=��v��( ��� %p/���;     �7�Zp��; @Z�  �j�6(��     �w�A��� @Z�  ���^*�;     ��{��E��(x[�� �E� �(Ke:Ţ     �:�y���<W H��  Q�&�$o    ��2p��5M  �C� �(�;     @�	����; @Z�  �rW�S-�     @�':o��v��3 ��; @��     ��N�[pi �t� e�     ����� @Z�  ���^��DW�    @�N4��Vw��u]o�s5 ��� � �T>w     8����2݊���mYp H��  Q�2Yp    ��:p�N���� �E�       @QN9'��  ��	� UUU      �|Չ�y[u]  �� $�Wg���     �6��p @Z�  ��     �����y� ��; @�,M��,     �7�6Mm�z���  �!p       �Wԭ�O&�   'p H���2���      �Ӟ��]����C� @J|{ H���Lw     H�n�ގ�j  i� @BZ�;     �����&  ��� $��D�ڶ     �8��1Ղ�۪�:  H��  Q�2�-�    ��N}�.p[w ��� 5��w     8���� H��  Q��Դm      �i���m�>�<�y��  �"p H���2�-�    @����x��?,  H��  Q��tq��e      Go1(#p;áD
  %�� $���,Mӄ�     ��{2]��۰� ��; @�,���;�~�E     ��[-�  �� $��Dy��     p��8m���n4�s5 ��� � �<]��
�    �h��a<  =w �Duk���7     ��V�  �%p HT]�AY,�    @��  �4w �DUU��;�v�&     �-eڶ}xy�  �'p H�p�\i���     ���jP�������   -�( �D�F���A{��w     H�����  �� $j2��x���f׶     gۼ�y{�sZw ��� %p/�o�w     8^�
�KQUU  ��; @�\_Y��ܛf     �q��� ��; @�,���w�     p�]�6�2�ӳ� ��; @�������~oѻw     x9��Q�u  ��; @��M���}��    �X����v���x� ��;  $��;     ���}�r�'p H��  a�� ���9����	��     p����w�{]��i��  =w ��u�������     �X����� H��  a݂;e�-pߺ�     ��ց;�3ʣ  R� @ºw������b?     m��K!p H�op  	s�b~�ݴ�      ��{�A��n���i  �� $̂{��[p    �c�堌�Ӳ� ���  fq��?�~�+S     o9(#p?��h  �E� �0�{����,�    �Q���]�~Zw ��� &p/����     p��ݿ����I��( ��� �0�{������     R�Xp/�x<  �"p H���������òL]     x>�{YF�Q  ��; @�\�X�<�����+�=     bۼm���t�6��1�S� �G �0W*��������Wy     8�f�{��g���Nc:�  i�M  a��$��?�]w��    �C���{g��	�Od6�  i�M  a'��]Qڽ~��     �����i  �� $́\��v�����;     ��C2��QUU  ��; @�\������C��֡7     �C2_;���u�;  �� $���,�����V]     �`������Ӱ� �&�; @���σ�}u�}'p    �C�a��1fsu]  �� $l:�y�z����     ��m�����OC� �&�; @ºk��C�|}�][p    ���aHƳ���F @z�  �A����?�߶�-    ��m,�C� �&�; @��F𜭯po-�    ��6۷_p�l�4�  i� $n8�v�����}-p    ��m[��� @z�  ��w�e�     ^�~���9���4&�I  �5 @�\����povw     8Ķ�GX.p?�; @��  �����M�~�`     ��mv�苦i������f�   =w �č�� _�Zp�O��|�    ���4�YN��_�t:  ң� H��=o���;     <W�ܿ���3�� ��(b  7�L�|}�p{�k�<     ����l���uvv  �G� ���l��{��mf      �M�כ�	^�t:  �#p H��=_�������l     x��?���_�`0��� ��� 'p����[V�    ���tC���uu�;  i� $n>�y����҂;     <�J�^��  �� $�ݻwA����7�me�     �m%p/�p(� H�or  ���fW,~/�&M�;�^	�    ��V�b� �� @�+��	����m      ϳ���|�x��L& @��  �(���n����     ����c��g5]�����i  �&�; @F�Q��� /�_p�    �s���^E�m۟�>G��<  H��  ��8���ٛ���n㡯�     �}��[pUggg @��0  ��fA~;����     �4��� ҥ� ��t:�����r��w��     �dݳ��m���\\\  i� d`>��y�`�o�     �g��ryy  �I� �yz�`{��     �4�r��� @��  ��鱃��F�     Oշ����\9\UU @��  p�b�]p���      ��o7�Zp=w ��	� 2��ݻ ?��[�;     <U����g4  �� d�[��^�����{��f     ���x3j�l������ @��  �����}��    �S�q8Ɗ��L& @��  ��(v��-�p���`a��     ��vMۿ�\��:��i  �.�; @&�C_�r�ءvw���b2��    ��,��[o︝�u���   ]J �L�f������Ֆ��F�     ���魨�_���y  �.% @&&�I�����ϭ�     ��,6�\p���; @��  �p�b~�r���+U    �O�=�۶^���e  �.�; @&,Q�婋-��^�
     }�<�,ggg @��  �x��]P�;�     �����?u���QUU  �.�; @&�����,zz�*     ���r�r( ���F �����?,RX���S?�Ū��3     �ݙ�b����s��7� ��	� 2�]�ؽ��	���+U    �/V�]�B�b�f�   mw ��tW.
����w�ӑ��     �5�M?��;�_�|>  Ҧ� ��d2��z��9�݊��     �n��o���;??  Ҧ� �H�Hq{{��;���     ����+�/���2  H��  #)���w     ���%y��}  �6�; @F...��,�     �M���_���u  �6�; @Fؕ��     |���PL)�ATU  �M� �W.��9�-�    ������[pY��(  H��  #WWW�C�r�^     �Ϻg&��.(�x<  �'p �Hw�b�j�&H۳���h�6jWn    �tg�mk���$  H��  3�Ջ��t1�b����C[     ��/�~߂�Vޗuvv  �O� ��n�b�Ze���     �G��MP����   }w ����󸹹	���Ŗ/�u�u      �c��,��� @��  �q�b��~@     o��yY��� ��	� 2��ݻ }-�     p��D�YpY�׮� ȁ�  3�)�0��~4     ������y9UU=�  H��  3>|�sg�     �`���v�D�=w��o��:  ȃ�  3�������,ˮmc���l<
      ��O�/g<  y� d����ߋ$|�!��A��     ��n�	�1�� �<� 24�Lb�Xe�[��O��     Hc���sqq  �A� ��n�B�����-�     �oR87?�y _wuu  �A� ��n��ӧOAY,�     ���n>�?��c  ��; @�����/�KP���*     ���[[p/ɇ �<� 2��?i;�@ۂ;     �ݮmc��e��*�C @.|� �п�˿�Yow��51�     %�[�1
c��e���   w ������~����n����<     �dw�MP��t  �C� ��n�b�Nc���#p    ��<��݂��8??  �!p ��l6��v�
     (���yyI��� �|� 2uvv�?�t�b���5     ��}������Ç   w �LuK��_�����2     �t����?  �� d�A^�n����_     (�r����	��=��� @>�  ��ӟ����@}׶q����t     P���:Ra��x��(  ȋ�  S�����ݚ7e�Y,�     �f�
�1{& ��; @Ɔ�al�� =�,�t�~     P��e:���㝟� ��ٻ���3��/ �)J")q�,K�▇�޻�\��]՗�T�S��$�'�<E�e��'� �igQ'qEX�y��w�<�������� ������sh�2     9��W������d  �_�  }l||<vww�lJ���v�����j     @^m[pϕ�g�  �E� �ǒŊ�ϟ�����w     ��lF� ;��
܏off&  �/w �>f�"ۊ�b�Z�#���f��clh0      O�*��I��x��'  ��� ������u�Ֆ��}�;     ��]�V�n��xJ���H  �	� ���=ێs���ۏS     y��d���x��� ��#p �c�bE�\�l6��9�Q{�R     ț�j-����񌏏  �G� ��FGG�\.�s��=cO�    �Iض��+gΜ	  ��� ��MNN
�3�8G�-�     �L�Պ��zd������� ��#p �sgϞ��O��s�gI�덨5�1<P
     ȃ�j-��vd�q������  ��� ����l�M�]nٮTc���     �<��ۏ,��~<� 066  ��; @�[XX�鸇�M�;     9��ųD�~<CCC @� �����(�J�l6�l9��     �"kw�d��w7>>  �'�; @���D�R	�币�Fe/      /6-�����T  П�  9p��)�{w�e�\�V�Er     �\����Fd���x��� ��$p ȁ3g����r�-�=l7[���ۏ���     �~�����q�n�nnn.  �Ow ��������:Ȗ�Xn٨T�     ������]��nbb"  �Ow �XXX��$ۛ彈ٳ     �l��Yc���  �K� �ɂEK��� ;N$p��b     �fe/�Ƃ��  ���  '���c?{�%yv�-����    �(�V��D�XpwSSS @�� �D��.pϖ�8l���;��ؐ�:    �O�k�Y|�V��� ��%p ȉd�buu5Ȏ�:lo��b���     �~��W�,������  �	� rbff&��� ;
��:�j,�    �S�l�R)8����s��  �K� �.\����+{     �j��Yd���  �M� ���Ӈ��V�dC�@�����c�:ɂ;     ��䆾���;���݌��  �M� �#CCC������J���f�X���~-�V��    �/���7�,������  ��	� rdllL��1'�'�5��j�L�     ����^d���ݜ;w.  �ow �9s�Llll�qR����/p    ��l�ewاT*G777  �7�; @��?>�߿d�I�ɂ;     ���޿���Gg� ��	� r�ҥK����qR��z�     �o�L����y3<<� @� rdbb���f�d�I.�7[�(9�    �'���_oD���ͩS� ��'p ș���(��A6�ԁ��j�F�3��     �`m7���&�D�ٳg ��'p ș��)�{�����nY�    @�X/�EVYp7��� @�� ����L<~�8ȆB�pb���nv�     ���|��]�Ʌ ��'p ș������d�I��v��T+     ��V���jd����J�R  �O� �3�����v;H��<p��עVo��?     �m[��h�Z�U��  �A� �3��tdd$��쮚��I��v+�p�t     @����E�%k����T  �w �����g��     ^�^�D�Yp?����  � p ȡ���XYY	��\�2�h     �5��  ��  �����޽{A�ub�     ���l�N�Y&p?�B��N�
  �A� �CKKKAv$G�f�y"�V�ވ��ZL�     d�zy/��vd���hFFF ��� ������O�^��$���NE�    @f���E�	܏���� @~� rj||<�����+�'��m����ٳ     Y�.pϝ���   ?�  9u��Y�{F���{u�     �U�l����[XX  �C� �S.\��w҇����l��t���     �i{�ß,���w �|�  �.]���y�~�ћ�vlU����X     @���f{�=a��h���N��  �M� �S���V��['����    ��Y/��&�N �|� ����X��� �:q�^�.�{s3     Y�����5�Gs���   _�  9v���{t��͕m��    ȖV��sgnn.  ��; @�%�G��։Cw�v���852     �k�{�l�#��o�P(���R  �/w ��v�Z��w�ҭS����S#��     ��uR�����K�  ���  �&&&���f3H�d�$�i�Ov�fe{7��
�    Ȇd�������d  �?w ������ ݒcw��8�_s�O�n     ���zy/��������  �#p ȹ���{t"p��ۏZ���     ����~4��EZ��ۻx�b  �?w ��[\\�����֩c���n,��
     H�~y��X,���
���P  �#p ȹ+W�į�� �:u�N��    �v�;��������h  �Ow ��:�988ҫs���x    @[�����ӧ �|� �������W���h4[1P�*     �S�E���``@����� �|� ������\�ޭv;Vw�175     �F�;������]�t)  �'�� ��/ƽ{����䓥+�w     �ke��B��v��EN�:  �O�  ���b
�h��A:u�ོ�?�7     ��U�{�  ��S3  Q,ctt4����tJ�u�?BX۩D�Պ�_~     H��A=v�k�/�o��ٳ @~�� ����)�{�%�q6��u�VlV�1=a    �tY��WH�ogaa!  �/�� 8t�x��i�^�ѻ�{be�,p     uVv*�O�1~���b  �_w  ]�z5���?��ɣ��v9n/�     H��>
ܓ!�B�������  �%p ��ٳg�X,F��
ҩ�ϖ&�{��vX     5j�fl��G��䝿�LLL  ��3  s�ԩ���	ҩ���F������x     @<��9g���3==  �O�  �M��.pO�N��m�
�    H��[��'��s�ҥ   �|r �o�~ҩ���[����     i�|[��7�B!fff �|�� ���r�J����{�N�>|/o�F�ՊR�     �K��A��k�O�lxx8���  �=�� �������a��_�~�t��v�ݑ_���_we�sS     ��lk7������;w.  �'g  ~fjj*����t*�J�h4:��?���    �sϷ��o�lii)  �'g  ~faaA��b�񻣁���_��B     @/=߶��GW�\	  �� ��y����C�N�>~o��Q�7bx�     ��ʋ[u?�����!��  8�S!  ?399��p�]�T���n�Wq.M�	     ��[������M  ��O�  ����ӱ���O7��6w�     ��3�{.���  $|z �%sss���J�އ_     ��v;Vw+�o�7�z�j  @B� �K�]�_|�E�>��w����b|x(     ��Vw*�h�����,��cll,   !p �%�ϟ�b��V����[O�>�܉�     ��y��2*p�ӧO  ��� �W������� }�Ƚ�ht��H�@�    �m�;��G�7�p�B  �_	� x�d�]��N�ܟm�     tS�ٌ��^��B�еZ���ի  ��3  ������ }����������FlV�qf|4     ��o���jG���Y�T����  ���	 �WZ\\<\i��u�:�'+�w     �ey��(������  ��� �W*���r�?��Y֭����v�^<     �O�v�	���  O� �k����S�[���N%��f�J     ��S���_~����ͮ\�  ���  �֥K����ҥ[��f�϶v�⹩     �Nz�ٟ��	���%/
���  �=�;  �u�������v;H�B��R)��f��'�w     :N��O���  �H� �k���HT�� ]�7���oG�     �F�����W�כ��	  �Gw  �hzz:=z�K��j���>Ճzl���쩱     �Nx���>}M6��'/��j�/_  �Gw  �hiiI��B�\{y��#p    �c�;t����zI����  ���  �����㷿�m��t9%��ŗny��\�     �	϶�y422�b1  �	� x��8<<���Azt3p_ݭD�ь�R     �IڬT�R�G�������  ^E� �/J�>ң��{�ޟ��_�=     p��l��z{B��zW�^  x�;  �������)�JQ(��nx��#p    ��=������5Y�|Ǳ��  �*>E ��nܸ���o�S�v�՗�����^ɂ{��?98    �I8h4c}w/���W;u�T  ��� �E�b1��ǣ\.�����Vo���^�L�     ��d�����:�k��/���  x�;  o%94~��wAzt{�%Yq�    pR����Yo��ׯ  ��� ��r��5�{�t�0�xc;>�<     p\�v;�m�F?
^��ڟ;w.  �u�  ���/F�X�V��C����^��bl�A    ��Y/��~��L��j���  o"p �%ǭ�� �P(��t˓͝�qa:     �8�n��z{B��jKKK  o"p �-,,�S$�ۓȽ^�w��|��%p    �؞llG���K�Yq���  �7� ��n޼_~�e��q�����͝�7�1X*     ��J� 6*��g����5���  ��'i  ������1��h�����f��6w���T     ��x�����CCC��Ξ=  �K�  ə3gbuu5H�^<o�����    �w�h}+�����.^�  �K�  Irx��G/���[�l��T,     �~���{���/+
q���  �_"p �Hnݺ����t�E�~�h��v9��L     ���h�����/���  �̧F  �d||�� Y�Ղ�K�N�cp����������    �#{��yЋ������	  xw  �lzz:�<y�Cr$�zྺ����a`     o��L^ݍ~����/�r�J  ��� pd�/_��Hr$�V�]�=��X�݋���     ���dc'��v��������ii)  �m� 8�7n���v����W+0�6�     ��Gۑ��_6>>�b1  �m� 8�dydtt4������ա�ǵ��立     ���nǳ����/���  x[w  ����\ܿ?�^����جT���h     ��<�܉z�y p�{�  ��  ��[�n	�S"yҳT*E�_$+�w     ~���ȋ^ӤU����L  ��� �Nb`` �F�{�L�Z������Vܽ4     �:�v;o�D
����ٳ  G!p ��%ɕ�����5�^j��kqjd8     �UVv*Q��c0G���+W�  �� �w�$���˃y��~{�|     ��<Zߎ����ڵk  G!p ��ݾ};~���>-Jo�4p_�    �z�7�"/���x��N�:�$  ��'H  ����`���G�\z+�wQ(z���T�zP�ѡ�     ���QދJ�y!p�����  ��� p,��7������j����IT�pm3n��     ��V7#Oz��j�$�<�n�
  8*�;  �r���{J$+��?��    xُ�ۑɝ�X,/�J����
  8*�;  �2==}x�����hZ�rfe���A�[�    �������8/���\�  ��;  ǖ(�={�V���3�w�     $�mF�?�z�j  ��� pl׮]��@����;     ���v���y2d��o
�B\�r%  �]� 8�[�n������X<00�F�'��zy/v��19:     ����r��{s���?����b�  �.�  [r���������u�^��W6���      ��l�=��$�ᅅ��  �w�5  'biiI��Iྷ�׳����M�;    @ε��x�����z��ݼy3  �]	� 8�oߎ/��2��v�;I��K�{��Y�ƙ��      ��n��A�y"p�I�]���D  ��� p"���bpp0���u���ae#�\��(    @^=\��z{"������	  8�;  'fvv6?~�N�T:�i6{�����F|$p    ȥF��7�#o,���ƍ  �!p �ļ��{�HVb��j�~���A��Vbzb<     ȗ'��h�"O
���+���g��` ��� pb�^���o��V��i��{�'~X��    ���խțdx&	��8}�t��  ��� pb�����Tlll���{������ʂ�>    @���x��y���|Z\�x1  ��  ��d�]��[��ý�K��A=V��q~j"     ȇG����+�###���~  �q	� 8Q|�A�����v�������~��_"|��!p    ȑV7#��0<��N��f ��� p�crr2�����I���j��׶�]��B!     �o�z#�wʑ7�BA���[\\  8	w  N��˗�����I��ܓ/3�n�����    @KFOZ�������s�N  �I� p�>���{���9����w    �x��y��{|�������X  �I� p����xT*��7�rP���F3�J    @��ۏ��^�Qv���  pR�  t�ŋ㫯�
z�X,���@4���u4[�x�����     �)���a��ܹ  pR�  t�ݻw�=��{�'��|]�    Ч��v���yT*�bpp0�nhh(N�>  pR�  t����᳜���Ao$�J��뿌Xۭ��^5N��     ���v9��G��_�p�B  �I� �1q����7�tX���_Y     �˃��ȫa�����?  �$	� �>�@��Cɂ{Z$_p|ty>
�B     ��f<^ߎ�J^�ͻ������  8Iw  :&9h&��z=�O��Z�'����A��Rb�vp�L���D     ��oE�Պ���133  p��  t���\���Ao�%pO�_^�    ����W��O�T���u�V  �I� �Q�o���P�S.�#�n����C�    �u��Z��V"���G��XXX  8i�  :��ŋ100�F#�4؛�V<\ۊ�    �l{��������H����{?  �!p ��fff�ٳgA�%O�
�h�ۑ���     }����ȳa�q���  �N� �q7o���Prd��ߏ4X�.��~-&F�    �*����"��a����b1�\�  �	w  :.Y���o~�V+辡�����q��\     �MV6"ϒ�{����ӧ#w  ��;  �8ϝ;���A��mE�����.^���     ��V<Zߎ<���v�Z  @�� �7n�{$m��J� V��q~j"     Ȗ׷��lF�����͛  �"p �+n߾���o��nݕ,�F�^�������     ��lDލ��F�MMM~�   �"p �+�C�����NU��pm+>�7bx�I     �b�Z;|�3ϒA�R�y���  ��& �knݺ%p���r9=_:4[�x���/�     ِ�Ιwɽ=�
�B���{  �$p �kn޼��y4�͠��xp��ٚ�     #Z�v|��y7::yv����W{ ���  tMr𜙙��ϟݕ<�:00�F#�b{�+;嘝<     �ۏk[Q�����+#9_pOƌ  ���  t��۷�=2<<���=����    ����ȻdLfpp0�*2�r�J  @�	� ��ׯ�o~�ԅ�y���T*�H���������G    ��ک�be�y7::y6==}� @��H  ����Ǔ'O��J�Ӧ�jŃ��xa6     H�/�d�����  ��;  ]�O��O�H�MM�UZ�V�ɷ���     )�j����� ��R).^�  �w  �nii�0����Aw%�2{{{�&�{�çmgO�
     ����V��Ȼd@fhh(�jff&  �[�  ����\���Aw�.pO|�lU�    �B^^^����۷  �E� @O|���H�4z���֗bx�Q     �b�Z;|��|�R)  �E= @O\�p��)σ���{���P(D�ݎ4i���`e#�_�     ���k�����Wɫ�  �Mw  zfqq1<xtW����G�|�lU�    ��v;�_��p8&�/�vï~��  �n� �3~�a|����[�w�3�iܷ�����=}*     譇k[Q�7��^Gͣ������	  �&�;  =3==}[W�ՠ{Ҽ2����    z���������W���  �&p ������K3i\����֗bx�U     ze�Z;|q����<J�K�s�N  @��F  詏>�H��e�A:�����#m��v�_^�ۋ�    �����Z�BrS�k�>44�Ν  �6�;  =555ccc���tOr�Oc�����J��0{��     �Uo6���F�BrO/��G�+�  �w  z����q�޽�{Ҽ6S��㍝X:w:     �+q�h/���F^}��  � p ��>����ꫯ��n�1<<|�8�j�"��z�,p    �o��?�k���}OLL  �� ���ӧO���V�=I�^�V#��o��V�S����     ��m��N���Ť�E�N�v�Z  @�� H���?~���ݓ���5pO|�t%�ύK    @w|�t5�I^���B|��  �"p  �ܹ�����V+莴��<Xވ�./��?�     t�n�v���O��OMM����<  ���(  ��<�y���x��Y����Q*���lF5Z����z�Y<     tַ�ע�n?�k��� @/	� H��?�8��_�%�dŽR�DZ}�d%n/�>�
    @gԛ�x���$���I���\�  �Kw  Rcaa!����V�ݑ���R;��;�t�t     �I�~�H�k��266y4??  �kw  R�ҥK���ݑ��U�z�,p    �o��?���y'ܽ{7  ���  ��'�|�}�]����F�^�GZ=�ڍ�J5����e    @'=�܉���U�Q����3g�  ��� �T����S�N���n���:́{��+�n\
     N�7��_���/��|�r  @���8  �w���������;��=��A������B�#    �II�۟m��>�ccc�Gw��  Hu  �������h�ZA�%�{�5���^^�;��    ����h���ύ��F�LMM���P  @� H�b�333���t^��;9ZD�}�d%n/�F�P     ���lƃՍ�ey�oݺ  �w  R飏>����#9֧=p�����v,��
     ����F���熇��a�$���v�Z  @Z� H��/���`�����FFFb{{;��ޓ�;    �1������Z𲱱�ț����.�  ��  �V�߿?輿.ҴZ�H���Xۭ���x     �n~\ߎ�j-xY��B�w��  H�;  ���'�ܻ$9`'+�{{{�v_>Z�����     ��|�t5xY2����dhh(fff  �D� @jMMMũS��\.�7::��������e����     �h��ˇ/e򲼭�'.]�  �6w  R�ƍ��?�1�$pςv��/���q1     8�{OV�W�c�~���  ��� �j�a������f:�T*>Ezppi��嵸{y>F��    �m�Tk�lk7x���122  �6j  R-	�gggcyy9�d�=�{�Վo����Ks    �����A��HB�d&On߾  �Fw  R��O?��>�,�$p��ގ,���J�Y<�b     �fՃz����Z��ۓ��ƍ  i$p  ������j�t���p��h�Z�v�z#�/�����     �;~�-����}qq1   ��  dµk��/�:/��	*�Jd����Ǎ��(
    ��՛����z�jɚy2 �'}�Q  @Z	� ȄO?�4�ݻ��e��R�^�?�Gk[qi�L     �j~�~��jy[o�������  ��� �	���133���Ag%�{�|�xY�    ��V;�y�����x���۷  �L� @f$+�}�Y�Y�b��)�Z�Y��[��[�qa��    �?�am3*�z�zY~9�R�׮]  H3�;  �1??###���tVr��J������    ��~j��M�{x2��������  ��  d�����/�:+9�ommEV<�؎����	     ^x����j�zccc�'}�Q  @�	� ȔO?�4�ݻ�V+蜡���gJ��fdŗ����s�r     �½'+���)p���8� ��� �)���133���Ag%+��r9�������|�    @�m��by;;7�^8|ɋ;w�  d�� ��IV�?�쳠���7[���x9>��     y��cC1�d||<�"y��ڵk  Y p  s���cdd$�����I�
�h�ۑ�>[�;Kblh0     �j{o?o�o666y����b1   �  dҍ7�O�S�9ɡ;�ܫ�jdE�Վ�/�'W     ���G�35^���K�i^|���  Y!p  �>�����/��j����d)pO|�l5~�t!��q    ȟ��~<Z��l||�0rσ����  �
�  �444333���tN�k�V�{�]�    ���ӣe��o!	������  Y"p  �>�����ς�)�J1<<�Z-���+q{a֊;    �+����qm+x�d�=y�4�;����  �D� @f������H��������������%+�    @~|�x%Z��Q�zi�X�<XXX���+  �C� @�ݸq#���?����5_?]�ۋ�c�T
    �~W�����������G^|���  Y#p  �����9���h[�阁������ȒZ��<]�_-]    �~�������R^�����  ��;  �688�����ɓ�s����//ǭ��(y~   ���ޝ>�Yh�>��-�؀1�;lll�l�Kg��d:==�n*5U���n:@��8x��]�*˖dk�۷�3�tX$Y����qT��*��`]��9/(�����>/��ͩ���?�y�  @%� P�������]X>E�>44�JS�����'}(     eu���L�Xo�����T��e�'�x"  P��  T����tvv����ayK�������J�)Vܷ?�&u�V�   ����ʩ�7���.�@� @%� P
�v��|�Oq�_�"(��-.w��    �l������������]ʮ��f��  *�� �Rعsg>���LLL��Q��{����e]�w    �TƧ���/@[[[���u����  �Tw  Jc˖-9r�HXŲM]]]���SiF�'r�ʍl[o�    (����f��l�j܋���{.  P��  ����?�cǎe�S�˦XqN%��lYכښ�     T�"l?y�z������X5oooOwww  ��	� (��p�xv���?,�J�G���Vܷ��    @�;r�j&����W5���~��  @�� P*�/~�<���R[[[�+�8?���Xq    *���T�Xo_�bټ슅�͛7  *�� �R���Igggn߾�^MMMZZZ2::�J426�׳��5    �T�/]ͤ��y����p)�'�x"  Pw  Jg׮]�����hmm����P��oYד���     T���9i�}A�a���)�G  ��  ��Ν;���gbb",�b����6333�D�����ky�ч    Pi��x%Sz>��TC�nݺ466  �@� @)mٲ%G�	K�X�)"�J^q���@���MC}]     *���DN]�毾�>���)��{.  Pw  J���ϱc�*ve|�kkk���}|j:G.]ɮ�    �R������Ά��������tww  �B� @)544�=�����^��^[[[� 8z�jv<�P���    ����z3,L5�O?�t  �L�  �ց�_�",���֌���RMLM����ٳ�     �t�����>MMM)�b�g��� �2� PZ===s�r�����Vс{�X���|dmZ    �R�˹�Caa�;��۲eK  �l�  �ڮ]�������ܜ���LOO�RMM�����o�     �T��d�z�������jjj�{��  @�� (�'�|2�|�I&&&��kmm����������1     +����\�q+,Lcc��W��_�>���  �ǿr (��y�#G������V����L�p�r�o},     +͗���}���w��  @	� (�����رc���	K���infjj*���������t�6    `��6<����yP��www�} @	� (�"�޸qcΜ9�^��~�Ve?�;;;�C�rpǦ     �_�W��444��jjj�o߾  @Y	� �
/��bΞ=;2��Z[[+>p/��v3?ذ.��Z    ���Wn���+�z{KKK֭[  (+�;  U���z�\�|9,���ƹ%����T���_���kOm    ������8eܟy�  @�	� �Ŋ�����Yq_mmmJ��pchn顮r_~     +[�����ݰp��ͩ�/oS��lݺ5  Pf��=  �'===����͛7��*K�^����yg��     <3�����H����;v8� ���  T��>��կ��*�p�՘���T��Gs���l\�*     �۱�k�S�����.O?�t  ���  T��{,����s�NXZŊ{�B�⾡�;�55    �_&��s�╰8����զM�R[[  (;�;  U��g��o~󛰴����7o�F�&r��Zv>�6     ��.\���Y�2�����d�޽ �j p ��<��S���2>�ץT__���挍����kW����M    ��+�7N\�S��K�e������1  P�  T��۷�СCai�e	��'��޳�     ,�/�dfv6,N��^[[��z���  �B� @U���Çgz�S�K��3[�K����d��k��d    X>7������a�:::RV===�^� ��L� @U*V\�x≜<y2,��	���֌����gf��������     ,�b��ū��OKKK�j߾} �j"p �j8p �N�*���JQ<[���p��`v>�6=�    Xjn���[�a�ʼ�^���Y�&  PM�  T����<��ùt�RX:��X˙��J�����y�m    XJ���W筷߫2�{��	  T�;  U�^�����3,����ܺu+eqyh8�7o��U�    X*���֝��x��JCCCʨ��6n�  �6w  �ڪU���ӓ7n��S<�Z����Y����=;SSS    �{55=�?\��M��۟z�  @5� P�^|����K���>MMMOY����+�ٲ�'     ���+�;1�$)Wʨ8g߱cG  �	� �z�֭�[xK��T(S�^���<�fU��j    �Xw&&s��Z�7mmm��-�y��͛K�� ��� ��ڿ���1,����fvv6eQ\:�x%�l\    ��:t�r��g½)�kʨ۟{�  @�� ��ڴi������hX�|���w����y]Oښ    �P��w�wu0ܛ����3�2�� @�� �������{/,�2~h`zf&�����;6    `�~�w�T/_>(e^o߳gO  ��	� ��mݺ5}�Q�޽�FKK�܊���t�����l[ߛ���y�    ,���n���r��<(e�7nܘ�F/� P��  �<��s�����)V�o߾�������ճ;RSS    ��353�/���{���T��8o޿  ��	� �?عsg>��3+�K��������ȝ��|=�֯	    ��9|�JF�'ý+�z{}��  ��  ��ݻw�w��]XsK:)�/����5����    �#c�9�5ܻb�V)���z���  � �/<�������3>>�Fq�088����ʡs����G    �m>?۟��p����RWW��y�G��b   �;  |�]�v�O>	K��o޼����]�뿚-�{���    �����p.ܸ�FgggʦXo?p�@  �#p �o�{��|��WVܗHq8_�ꌌ��lffg�ɩ�y�m    �����ߟ�K���>---)���ק�و
  ���  �œO>�/��",����R�[`ʆ��     �щ����FWWW�h���  �D�  �b�޽���399�]cc�����D���������    `bj:__��F�Rh1�R6�֭�{  ��;  |���ڹ����*,���������s���`ú     |q�?�S�aix]]]ʤ��8  ��	� �;�۷/����T�wE�~�����Φ�������!    @��9z7���s��A���L٬Y�f��  �sw  �Ŋ�����"w�]�FS�쌌�����g���Kyi��    ��gg.�v��A���OKKK�f���  ���  �G�<���ǭ�/�����+7�m]o�vY�   �jt���\�U�3����+e���[ʟ  ���  �G��e˖;v,ܻ��ƹ�����է}����s��    @���W���*�S��?�a  �o&p �yx�r���LOO�{W\Fܸq#eucx4'�g��k    T�C�rgb2,������եLV�Z����   �L�  �P__�'�xb.r��������MY}~�R6�v���!    @�����������J�8p   ��� �<�������jjj�"��������t~�w1wl
    P~�������z<��LKKK��z;  |?�;  �Sccc�mۖ�G��{���Q���p��`�X�:��.��    �'���ȵۣai�q���^  ���  � Ŋ�ɓ'355�M��kbb"eV�6�������    (���|yn ,�b(�L֬Y�իW  �nw  X�����ر#_�u�w��č7Rf�w��������p    ����̥�OEYjmmm���K�8p   ��� ��߿?'N�(����P\Pfvv6e��������jm    P�n����`Xz]]])�u�֕�g ��"p �*Vܟz�|��������E�###)����|r�|�|f[    �r(��>��^CCCZZZR&/��B  ��� �"�ݻ7����d�7�����C�9{mpn�    �|G/]��ѻa���e��#�̍�   �#p �E(Vܟ}��|��'��K<���K�}z�b^ՙ�z�   @%������W��Y����y�� �¨*  `�v�ڕC�UE���:::���xwb2_�Ⱦ�    T���.fjz&,�"n/Ff����y  �O�  �`߾}���½immM}}}���Rv���eӚ����-    T�����XeZo/B����  X�;  ܃;v����}�ܹ�M��~��͔���l>>}!���>�4-    P9�ff�Yߥ�<�1���ƔŦM�J��  ��"p �{T����?�s�7���������hN\����    �89��aytuu�,�������  X8�;  ܣ͛7�O>���HX��ֶ����=~q�?��v���!    ��74z7�������0��^[�lI}�,  ÿ� `	����?���T���r��쬚�}bj*����W�|"    ��V��~�w133΀�K������  `q�  �{�ttt����a񊅞��挍����~3��-�    +ױ��v{4,�����3��عs�ܫ�  ��� `����������{S\bTK�^����<�՞��   �J4:>�C���)^�,K^__�ݻw  X<  ,����g�������:w055�jpwb2�?s1/l{<    �������	˧���駟��v  �7w  XB�/����Ά�+V�o޼�jq��<�fu^U�K    (�SWnd`h8,�b����1eP�E�  ��;  ,��kצ��7׮]���ޞ��������N��}��4��    x����8��WWWW�b���  ��  �ث�������W��/^�|k[[[FFFR-F�'�����ۼ!    ����鋙��˧��an��ZZZ�cǎ   �N�  K���;6l������uvvVU�^8�-{WemW{    ������0x+,�2���߿?  ��� �2x���������LX�b����9ccc�����N��O�<��ښ     ����t>��WMMM:::RE�_�   KC�  ˠ��1۶m˱c������n�ˡ�y��    ���]���TX^�+����)�_|1  ��� �2)�O�>���ɰ8���sK���;<|�r��NO{k    �����휽v3,�b��z����  X:w  X&����ݻ�駟��+V|nܸ�j23;��?��zv��T    `�MM��Ӿ�a����ύ�T����<x0  ��� �2*����:w�����֖���LOO�����#����    X~_�����DX~eYoߴi��K�  ��� �2+�[���1���a������Ƚ�|y�?z����    `�\�=��W��%����%��ͩtuuuٿ  ��'p �e�q��tvv�֭[aq�����Uۇf�����sy{����    Xz�9�G�.�H����ݝ2xꩧR_/� ���_�  p����������8���ioo���p�M�u|�Zv<�6    �����@n�˯��1����t�ϱ{��   �C�NU�  ��IDAT�  �Aooo֭[�˗/��)V�1p/|�w)�;��Z���   �JRL����ٳ'  ��� �}��k��o��o<s�H�S�mmmM����ɇ����۵#��5    ����L>:uޙ�}RWW7�Rg�+~�m۶  X>w  �O�C�M�6���/,N��^��{����x%O?�.    �����K�}w<��z{MMex���  ,/�;  �G̹s�2==���1���K5��|^Ց���     �704�SWn���Ë�J�z��_�>  ��� �}T�O=�T:�����}ff6�9q.�����V��    <(�������p�tuu���6���_  ���  p��۷/Ǐ����o���e��FC�w�չ����H    ������ܙ��O�W�G}4  ���  �b����?��ð8Ŋ����S�_��GVw�.�)    �o�쵛��)������S�s�^x!  ��Q�A  @�ڹsg��⋌����kmmM]]]���S�fgg����_�>�����    �����puww��mݺ5���  ��;  < ̯~���p555s+�7oV�����x~�w1�o},    ����ԅ�OU�hƃR��466����ū�  ��#p �dÆY�vm�^����=�n����L���ky��+���
    ��N]��K7o�����{��Im��4 �~� ���o��?�yUGڋU\(�����})����_�>���   �7���g�����Ԕ���T�����ر#  ����  ��x�u�֭9~�xX����gvv6����d>9}!wl
    �犳�ߝ<����p�Z�*����&/��R  ��O�  Xq@~�̙LLL������[q/"�jv��`����5�}a    K����\�5���ƴ�����[�.k֬	  p�	� �����������������HU��>:u>k�����     �}w,_��_�����  �`� `ؾ}{����ܾ};,L��^,�{5���G'�絧6    ����l~s�\�gf�����0��f%{ꩧ���  ��� �
��(��n�/�/F��>::Z���7�r��Z�?��\    �ۗ�28z7����^���>�l  �G�  +Dooo}��\�p!,L}}���Y߅��jϪ��    @5α�k��+�j;::R����  ��� �
����g?�Y�����+��dzf6���O��L]mm    ���ON�w'��K�F����^�:�=�X  �K�  +Hccc�y�|��aa���>::�jw��X>뻘緸�   ��|t�B�NL������kjj��+�  x��  ��<��s9~�x�ܹ�Xq��������l��
    T�c��rq�Vx0����"�J���Wt�  e"p ���_ί~���0imm����g�=;���    (��U�/�����.����T����/  X�  �mذ!����~�zX�b�]��o�'����y����    �ezf6�9q�_�;�J_o߻wojkk  �w  X��x�����?2;;毱�1---�{�nH����+���u   �2�����u������H�jkkˎ;  �w  X�:::�e˖�<y2,L�$p��/��g]wGz;�    erq�VN]��J_o?x�`  ��E�  +��/���g�frr2̟�?73;����O��LC}]    ��NL棓�ÃS[[����T����g�ڵ  V�;  �`����������)�������x>>}!/m<    P�fgg���3>5�b��8ǮD��]��   +��  V�;v��/����p�����477gll,���+7�pwG�x�'    PɎ\��˷��>HE ^�T��۷ϝ#  +��  *�o��w�}wn���+.W��S���ٞ�7    T�#wr����`篕����ؘ�{�  X��  Pz{{����̙3a��w+�njz&;��wmOmmM    ���[�=q.33�@�"l���N%����K/�T�q>  T�;  T��_=?��O399毸d�|ٚ�t}x4_��ϳ�	    T��O_�����*�]+5_�vm}��   +��  *DqY��/�׿�ufg��WSSSZZZr����'�p9������    �'/_��k7ÃU�UwuU�b���k  V6�;  T��[��СC�W�		���oO��O��L[Sc    `%�9z7�?��U�VU�z�3�<��F�  ��	� �¼��[�ۿ����̄�).,Z[[s�Ν�'�S��Ѿ���m���)    �orz:�;�ig�\]]]Ů������  ��'p �
��ё;v�ȑ#a��w��_�~{4_���s�    �D�;y>#c���[�zujjjR�^}��   �A�  ���������X��������ett4��#��dmW{��    �$G���[������`�D7n��� �� p �
T[[;�6�_�*��W�gggß����j��_�   �����h�<�V�J]o������  T�;  T�6d����S,+�###��MNO���}y�����    <HS�������X�2+q�����΍�   �C�  �7��_��_gzz:�O��>::j�����O�.f���    Jqv����+C��^����[�  �,w  �`���ٻwo>��0?�s�����D����h��    �×�f`���J���8w�Zi����^{-  @�� @�۵kW�9����0?�jO������>:u>��[���    ����ɡ���Q���۶m��0  � @)���y��w��T[[����ܺu+������h_�yvG��    ����T~{�s����)mmm�4���o߾   �I�  %��ۛ�7��ٳa~��}xx8333�/ݺ3��N����    ˭�ڋ����dX9zzzRijjj��/��   �I�  %��(?��O39�h>���>44�ٙ��y��=�֯	    ,�C.g`h8����iiiI�Y�vm}��   �K�  %Q�����|��o߾m��;|z�Bz:����    X�7o��ūaeY�zu*MqN�ꫯ  �lw  (�;v����߯x����+7o��lzf6�r�t~�gg��		   ����oO����lX9Z[[+r��駟NSSS  �ʦN  ��y뭷���V�穣�#��Ù��
߬�d|�h_�xz�܇    `)L�����g2>�ln����I�iooϮ]�  T>�;  �Ll��?ȡC���+�����\�~=|����|q�?{6=    X
�;y!��w����ٙ���T�����_  Pw  (��>}}}	߯��mn�}||<|��/\����<�fu    �^�t5��+K��^]y�۶m�2  �A�  %���8���������ˏ+W���������Ҝ���    �b\�W���S����ե�477ύ�   �!p ��*Vv�՚cǎ��W\������]O"�陙�����ɞ�ij�'%    3:>�O����lXY���W�_{�   �F  �{��s���ܹs'|�U�V	�硸�|�h_�xz�ܓ�    0�x����d|r*�<�hJmmm*ɦM��f͚   �"p �+.#�|����̬E����А��������604�/��gϦG    ��ѩ10�g�����$���s#/  @�� ��֮];�b����_�������.gu{K_�:    �]�^����n�����'�楗^���y  `~�  P^{�\�t)������ե��+CCC����Ĺt�����%    �M.��saejnnN[[[*ɣ�>:�  ���  �@�b��������+�����t�nS�3���O�'{v�����    ����|x�\f���b����������_  P^�  �Ś͆r���jjj��ݝ7n��W\R��/o<�u�w    ��ټ�L�'�����ޞ���T�^xa.r  �˿� �����[��O�����݊��۷o�]��@�����<��    @��28r7�L�X��իSI֭[��<  @�	� ������W^�����7|�U�V��իa~�p�rV����5�   @u;r�j�������+�uuuy��W  ���  �̦M���C�ʕ+ỵ�����9ccca~~{�l�Z����%    T�?����U��tww�Rk����Kccc  ��� @z����,����+�a~��g��_��_�ٙ�r   T��w����3������Y��s�b�R��m�  T�  T�b��������w+~Wmmm�3:>���T~�k[�kk   @u���ο9=�_V����tuu�Rk��z  ��!p �*�s��=z47n�߭X�s�Nfgg����o���+;�    �733�����[pge��驨u�ݻw���5  @�� @{�����<333��O��FCCCa��]��C�yf��    Pn����˷�����Ғ���T������?  P]�  PŊ՛�{���O?߭�H���T��/�����)�֮    �t��՜�V����T�be�G?�Q  ��#p �*W<���ח7n�oW\��Z�*׮]����"�ގ�    P.�7o狳�a�+F<S)v�ڕ���   �G�  �w����s��ߣX�onn���X��陙�w�t�yvGښ*�   ��v��X><~6���ae�����Օ��bwww�y�   �I�  �E�/��B����݊K��~�Tuwbr.r{�����   ��6>9����ebj:�|Źf]]]*A���  ���  ��}���8q"�/_߮��a�Y����0�#w��3y��'RSS    *���l��h_F����W�ivuu�����{M  �^w  ��y���������d�v�󸣣����	s��P�8۟=�	    ��S�s��h�������Z��   �M�  �?Œ�+��������l�f��E�>88�����ܘm��   ��r��@�\u.V)���*f���.?�я   p  �̦M��裏���uttddd$a�>9}!�-�Y��    *���C9t�r�555���I�8p�@   p  ��[o�����g�nժU�r�JX�����������t�4   ��mp�n~{�\��+�ū����G�O<  ���  ����y��������577�=�{�Ν�p�S�y��鼽k[��y
   �Rݙ��{�Ogjf&T�����������W^	  �)  �o�裏f���9}�t�v�W��ݻw3;;nh�n�;җ7�ޚښ�    ��L#�O���d����sC&���_���  ��_  ��z��W���?p�͊%����ܺu+,Ε��|x�l�x<5"w   �cfv6�;����+I��d{{{*�ƍ��V   �#�;  𭊅���~;��������Օ���LMM��9{m0mM����,   ��⣓�304*K��^	�����  ���  �w*.Cv�ؑ�G��oV��www����a�_��֦��|dm    x�>?s)}WCe)^�ljj�JW�����ks#+   ���  �^/��R.^���akMߦ��-###��Y�Ŵ55���    �`���#����R��W�N%غuk֬Y  �o"p  �����/~���̄oV\dvv6,N���ؙ���֬�l    �ץ�����b�<===����J��ښ���  ��� �y�����ݻ��矇o���0��[���M��佯O���;���    ��w���3*PSS���d%x�7  �]�  ���ݻ7}}}
߬��+������
�7>5���d�yvg���
   �܆���ޑә���c%Z�fM*�~���1  ��   �w������df�E�7�����իs���poF�&�"�?�=�u�   `y�ON�ç36i���x���� {��	  ���  ��֖W^y%��^�f---imm͝;w½)����Ѿ�������   ��553��������Py���jժ�tuuuy��7  0w  `��lْ�'O��ŋ�+�ccc�����[����غ1    ,��������\����7��+������ύ�   ̇�  X��������ܽ{7��b��xr��͛�ޝ�����<���    �4>�7n��T�ŋ�+݆�y��   ̗�  X�b���λ�;���_������h&&&½��l�\����    po�ȉ��2���̭��t���y�W  �w  `ъ�ݻw�/��l��չ|�rX�;y.-�yxUg    X����9tޙU%[�jU����o�97�  �w  ��<��s9w�\�_jjjJ{{{FFF½���Ϳ>�7�ޚ�]� ��ٻ�/9�3��w眣��X�!
!$�P ���?p�Ú��0��$�s@����\������P���:��>�խ�9����} ��|:4��,_I������ʅ�   ߖ�  �iO?�t���G����%�8�����f��������������Z_    |3�����";7,_�������-���   �.�  �M�����<>��do��c6��_~r&����h��    ����d�{�|d���嬡�!jjj"������ݻ  ��  �b�ڵ�~���p�B�����cbb"�����1�J�[G?���*   ��665�;�L&X��A�d�|��#�De��:  ��  �&�������Bn�Qkkk���Ɯ��f|z6���I�U��   ����T�u�lnX �[�'����ƍ�[n	  ����  �7���{��K/��l6�����hll����`��LN�[��ƞ;7GyYi    �T:~�ə����������b>�����z(   n��  �W---q�������555�&ܧ�&fͧ�c�5ۻ���%%   P�R�Lnr���L�����Dggg�d�ɓO>   �A�  ̻��;.^���%�Q�*����`~����{��ǎ;6��  ����f���chb*X�������2�Ur����?  `>� ��o߾�����F*�
����:���c||<�_WG�w�/�C��   �b���ůN\��1gO����"�53�%����   �/w  `A$/�J�W_}5���/K.����"����\�`T���}�   @�����:<�$/��m��9�]�  `>	� ��bŊؼys�:u*�����hkk����`���:5��mMw    �?��������Ԕ���v�����  `~y�  ,�G}4z{{cl�Ԩ�WSSuuu111̿#��&�o^�    ��K�q��0�B�D㭭��϶l���L   �O�  ,�����?�t:���jjj*��l0�~�J.r_בߗ�    7�T����J_P8:;;s[ �UKKK�w�}  ��  ��K&�?�����o���\�W�%U�_�~=����oO]��X��    ��l�`��ܕ�p444��T�U2]��'�  ��"p  �ڵk��n��'O_VWW����/�_&������wl�   �|�`�^�^P��ʢ��=�ٮ]����2   ��  X4�<�H������p�e������f����"r|��X��    ��������LGGGn�c����;���+   ��  XT���G�J���J&3577���P�0��������m����!    ����G�7�.FV�^P���s��U�o߾=   ��  XT���ݻw�k��f���ihh�����$wF:������]�6EW��   X~z����(���������"v��   �A�  ,�U�V�V�~��������EOO���3I�~.vo�5��w"   ��K���N���$nO�<棒��x�'r�K   ��  X��\�z5��*//����N*��_=���m"w    ���܈�N\�LV�^hjjjr��Q��{ߋ���   X,w  `�8p ~�����l�W���199333�M�s��w�m��   ����s��3�lPX��<��񮮮�6N  ��$p  �LEEE�ݻ7~���Ŝ��_���}}}~.l&��_~r&����h��   �|sml"�9v>�q{!jkk˝�棪��x�'  `�	� �%�����sO��O
����2���bdd$XXI���G��ɻ7GSmM    䋡��x���He2Aᩮ�Ν�d���={���4   ��  Xr۷o�+W�D�W�����T���k:7��l�{s4TW   �R��_=�iq{!J򮮮�W��{o���  �R�  ya�������s�������鉹��`aM����NǓw��Օ   �T�'��-q{A������L6V�^[�l	  �����  �����ݷo_��'?s���+��444,�\���\�^W%r   ���L�}�\̈�Vmmm444D>�����{,   ���  �ɴ�x ���௒ˮ����o|z6���L��֨�   �hlj:���lLͦ�����|TRRO=�T�5  ,%�;  �W�n��.]��W����===��f���\&������E�   �������(++�|t�����dy  ��� ���L	�я~db��H.�ZZZbpp0X3�q��S�����P]    eh|2�:v.fR�p�����Ѻu�b���  ��  @�IV�:t(^x��d2��˯$�������l��t.ro��   �ohb*�:z6f���
Y2����=�Q2���G  �|!p  �Rr��k׮x��7cnn.�\kkk����Q2���OƓw�M��   0_���<z6f�����3�����ػwo   ��;  ��֮][�n��G��K.����ڵk��N�㍏NŞ�6Gs]M    ܬ���x���H��^ccc���F�)))�'�x"��u   ��  �k<�@.����>�\�������D�xr��ǧ�m����.    �����x���Hg�AaK&����E>���r��  ��  �{����^��7�)���ӑɘ�fR�x��ĝ��]�   |=�c�މ�ɊۋA����F�I�g�~��  ���  @�K.�8/������$?���v���l:���L��vkt4��  �o���|d�sA�knn�����7�cǎ   �Ww  `YH.]v��o��f�͹ LTWW�~.7n��l:o~r:ߺ)��   �_�:�yܞu�U***r[�Myyy�ݻ7   ��  X6���[�n��G��kii����H����Jg���ѳ��6�;   ��.]�ߞ�(n/"]]]QRR�$y=O<�Dnp  @>�  ��<�/>��joo����`񥳟G�m�+[   ��]�6$n/"�������7��{otvv  @��  �΁�?��?brr2��eYsss����/���9v.ݲ>ִ5   �.��g.ǜ��h$�ѓ���&َ�e˖   X�  ��SZZ�^x!2�L�����ӹ/_&������wl�   9�{���_���ܲ��+�MCCC�ر#   ��;  �,%�2;w�z�%�ioo�����f���K֌�{�|�ۭ�ĭ��   �c���_.�ť��#���+�H^�޽{  `9ɯwV   �����c�֭q��� ���,����ڵk��H>l�ӗ"�����oZ   ���\�ǯť��1���#����Į]����:   ��;  ��=��100��"���6w�6>>,�?��4�S����U   ���?w%��ť��"�]1�|�{ߋ�.C  ��G�  ,{���G155D������L�R�`�����LܿiMnZ   P��ss����HP\�s����;�Y�fM�y�  �	� �e���4:/��Bd2�(v�eZ21���/79��s��Z�>��|h��~O��   ��L6~u�B��ŧ��-*++#�444�Ν;  `��  !��y�����u&�Tknn����`i]�Mr�qǆ(/-   �p$���9~.��Mŧ��6���"�����޽{  `9�  cÆ144~����3���1==SSS�Һ:4�?:��m��
o�  �Lͦ��c�bx��K1*++�����'�f�={�Duuu   ,gn� ��r�����`\�|9�|Eroood2�`i]�1o|t*��ks�VV   �|�O��[G�ƍ陠8uuu�"�|���F{{{   ,ww  ��<����/榹��-����729�x2vߵ9��   X~F?{��퓳��8577GMMM�-[��ƍ  �� ��t����������t�䲭��!nܸ,�d������w��u�u
   |�������1��-�XUUUEkkk�U�V�}��   �B�  ����x�g�^�LƅcKKK������l���fS��ǧ�񭛢��.   ���7r#�=q>ҙlP�JJJ���+�g������;w  @!�  +�Z�{��x�7bnn.�Yr����===E���3�t����x쎍���1   ��u��p��Rd��U�Yr�VQQ�"�q���(--  �B"p  
ښ5kr�y���?D�+//ϭO�C2���g����Ǻ��    ��ɞk��W(rɤ�d�F�H����z*w�  Ph��  
��wߝ��ϝ;�.��������� ?d���W'���䊸{��    ��Ǘ{?���[2�=�ޞO}��hnn  �B$p  ���?���q���(vmmm1;;�T*�]��t&�ݰ:JJJ   X:���?}).^�[rN��Օ���/����rK   *�;  P48�?�|LMME1K.咉S���Vk�Wbbz6ٲ>����   �I��wO������������|�v��\�  P��  @�(//�C��/��L&�Y�V9��n�}��<8o|t:vm�U޶  �b����w����������룱�1�ESSS�ر#   
��r  ��444ľ}��W^)���uuu1==�㦑��7&���'��5�3!   
���T�}�\LΦ*++���3�E2E~�޽  P�  @���z(~���}��������/�ˍ��x��S���M��P   �����:y!f�Ž��ϕ��DWWW��|PVVO?�t.�  (w  �(mٲ%�������Q̒K�������l6䗩�T���xtˆX��   ��;�?���lqB௒�|�ɓ�;wF}}}   �;  P��)����Ŭ��<����ڵkA�Ig��αsq��5�yeG    ��dϵ���O�����/���X�re   �;  P�����?�|LLLD1����]�ݸq#�?sss����1>3�_�*   ��������O�t���/$S����#_lڴ)��  ��� ��VZZ?����?�q���D1kii���٢�9䳣W�bj6ܺ���ݒ    ��d[گO]��Cc_H�	�����$?�\�����  �b$p  �^uuu<x0^z��d2Q��˻������l6�s��193�ݱ1*��   ��fҙx����6V����G���QQQ����>v��   �J�  ����طo_���Ew�����0��w�F��t�ܺ)j+���   ����t�}�|�O�^Ǘ%g�uuu����r�8���   �J�  �_��;v�w�}7���X���Dccc��Yӝ�oL�/����[7F[C~\�  @�J>,��c6��[IP���� >���(/�r   �ͻ"  ���iӦ�q�F��O�b���333�/���l*^��T<�y]��̏�X   �7g�����l�4�%Sғ�%%%K�Rr�婧�ʛI�   KI�  �w�oߞ�^~���(f����l6�_��\���ܚ��׮   �sɆ�/�ƱO��JWWW^LKO�Gy$���   �;  �WڱcG.r���b��D������܅0��K�165n^e��   �,���oN]��Cc_���5jkk��e���{�7֮]   |N�  �O<�����/���H����hii���� �]���عuSTWx�  @qJ��s�|�NN|�$lOμ���͛c˖-  �_��  �'JKK�СC���8����X544���l�������D�z�D�ܺ1Z�~
   ,��}�{'��t*�U***���+���5k����   �L�  �5*++�?�A.rO�RQ����I�|��&ff���N�#���5m�   �����ݙK���|���������Xj��ͱs��   �	�  ��de�����_�l6�(����쌞����,7�L6�=~>��[��t   ��/�~���u����@��VSS���   ���  �H&��ٳ'�x㍘�+�)`eee�Ƚ���h�M��t��ո1=�o�%JKK   
I��ߞ�WG�NKKK���-�ˈ���8p�@^L�  �Ww  �oh͚5������_��wUUUn}���p�|��c�������Q    �ar6�?C�S_'�И�XjIԾw�ި��   �9��   ��w�7n܈�?�8�Uccc�R�������Ň'�񭛢��%*   ����d�{�|.r���LL���Z�%%%��O�G   ���   �����###q���(V�ī�����Ǎ��x��S�����!   `9�pm8>8s92�l��I���������~<�@�   �	�  ��'�|2^z��b�\�uttDoood]&/+3�t��3�}��ضƥ*   ����\|x�7�}��MtvvFee�R�����cӦM  �7#p  ���y�x�bll,�Qyyy��?w����}�p5�����뢼li��  ��2���oN^�ޑ�DKKK���/��ȅ�w�uW   ��	�  ��d���>���'''�UUU�.������������[7F}uU   @>J>����b|z6��������֥~�f͚x��  �oG�  p���=�\.r����b������1>>,?�S��_N�#����-�   �$�p�g.G:��&***���k�_Ftww�Ν;  �oO�  p�����?�A.rO�RQ����r����L��̤���O�Ķ5�����   �Zvn.>���>���JJJray�yq)%���   |7w  �yPWW���_~92�L��򰣣#z{{���/G�����t<|ۺ�(/   X
��}�b���6�����ť���O?�t   ��	�  �I2�i߾}�ꫯF��f���Gggg������\�<]�_|x2�cc4�V   ,����x�ą����6Z[[sC(�R��1�ۗz�<  �r'p  �G�
�ݻw��Ç�2򮪪�����~�z�|%Sܓ�����ǚ��   ��p��p����H�� nN}}}n��RJ&�'�z�<  @!�  ̳[n�%v����^QF�Ʌb*�����`�J�3�α��mMwl_�2JJJ   Bvn.>���>�������V��TVV����   ��	�  ����333��e�L�J��111,oG���&�?tۺ�,/   �O3�t�������m����6*.���駟�}   `~�  ȶm�r���#G�����"��g��vep$^��d�ܺ)jL"  `~�O�{����l*��J��+V��RZZ�w����   `��  �=�����q���(6�%c����7����LN�+GN���ƺ��   ��q~`(~�Jd�ـ�+*++��5<��c��/   ��  `�=��C111�.]�b�L�J.����"��z�Ke2��o�#�۸:�JK   ��t&���|W������%}?�p�^�:   �w  �E�gϞx�Wr�̋M2I+�t
���k�5�;�l��꥝�  ��165����UCCC455-�󓭅۷o�6   C�  �H���/��rE��������6��Pޘ�W���o_�Z��R  �����P��ܕ�w��������cI_�w�۶m   ��  `����Ƴ�>/��B���E�I&k�R�
�L:o=[Vu�=�W�;^   �2ٹ��ūq��Z�ͨ���+V�&�/�M�6�=��   ,,�;  �"J"������8&''�ش���"�����p��:C�S�Ȗ�Q[Y   ����_���S7#9SK���ϥ�v��x��  ��'p  Xdɴ��{.7�}zz:�I2a���+z{{s�;���F��������ʖ�   ��]��\��t:�fuww��ԖʪU�bǎ  ���  ,����������ܓI[�����=���c&��_~r&�����V.��p   �Fvn.�\�'{�̇������Y��'q��]�  ��#p  X"I���$����(&�ĭ�rr`` ����r�J_ޘ�G����
G   �bb&�>y!�ߘ�����ظt�����cϞ=  ��r�  ��jkk��������Yt�{2y���%������;2�9���;�  �����h��R̦3󡮮.��ږ��ɳ���   ,>�;  �K.�I�/��b�E���L&���Aᙘ�����;o鎻nY%%%  @a����6y}r�ߖ6�MUUUtvv.�󛚚b�޽  ���  ����8t�P���ˑN���$Sܓ�}||<(<I��ѥ���o_5�  @aH>���S�b`�{z�Oyyy�X�"JKK���I�~���%{>   w  ������<�L���?�T*�$Y��D�SSSAa��?���x�u���)   X�._��^��t&`�$Q�ʕ+���lI��l�  ,=�;  @I��<x0~���bQRR������Aa�N�㭣gc˪����UQ�  `�Ie2q�BO��0���dr{E��l���˝ˉ�  ���   ϴ���.�~���U�\vuuEooo���p��:�[_���룱�:   X��'�7�.���L�|K΅���� �۟}�Yq;  @��  ����ؿ���?�l6�"Y?�E�^L�w1�1?���$�d�;   ��dϵ8r�jd���[r�D�K!��:$n  �#w  �<���{���^{��b�du����ǜK�������D��x�ֵQU�   �L�����K�3<�ZZZ���iI�����<�L��;�   �'ޥ  䱕+W�SO=���zQE���b2��ڵkA�|}$������GWS}   ����g.�L:���룵�uI�]UU���+++  ��"p  �s�V��'�|2��D�d-u:�������O���O���]�+���$   X��\����8���,��������D��  �)�;  �2�z��صkW���[E�'�3�L��Y�^���W��o�F<�e}�WW   �ktr:~s�bOL,�$,������{���6  ���   �����2rO�T'��'''��p��D��ȉ��-��si֔  ��C�W"��,����X�bE���.��+**rq{mmm   ���   �H�?���_���"������닙���8�ҙ����?z#�۰&����  �X̤��3��ӡр��D�+W�����O��   ˇ�  `�ټys����.��=YW�������J���q��z���÷����   `~���g.����,��|���;*++���3��   ˇ�  `ڰaC�R0�ܳE�6<����ٙ���d��113o||:���{6����~�  �9��#{�L���Ő�����,�s��   ˏ�  `�Z�~}�ٳ'>\4�{�J:��D���=�W'��&>|��h�w)  �]����N_��3����-�����I���3�Duuu   �|�  ��5k��޽{��^+��;��L"���������x�/'��]�+���4w  �o*����/���177�Z[[���yџ�D�Iܞ�%  ���  ���+W�����W^)�໪�*����ڵk.�P����W��o�F<�y]4՚�  �ޘ�ߞ�cS���x������eџ[SS��  ,Sw  ��L4?p�@.r�d2Qjkk�;r�8]��W����׮�������4w  ���|H��Ձ��rod�>$��ihhȝ�,�$n��g��\  �\yG  P :;;s��_}��H��Q���rS�������ȅ����h<tۺh��
   >7:9���>4>���3��j���������   ˜wu   $�8|�g�'?�I�D��4�dj���HP�F�s���Y�*6��  �bw��z����Hg��)���l\lIܞ�����   ˛�  �������0����E�777�&�����+���g.Ǖ��x`�ڨ��  �b313�������*������dQ�����  �;  @J��db�O��H�RQZ[[s�����bwuh4~������k���   (����>�T&��***bŊ��'�`����  �;  @�J&�?��s��K/���l����\�>99��T:�=~.6t��}�DU�#  �p%S��J��l��(//��+WFYY٢>W�  P���  �������gff�tttDLOO$�����u+c�   (4g��Ǒ=���d��=�ۓ�}1%����   �;  @�����E�/��bQD�%%%��ٙ��g�$���%��?8s9��ƿ�zK�UU  �rwcj&>8{9�G��J29}ŊQQQ���M�ݻ7   (Lw  �"PWW?��s����d��r���+z{{#�J$�����|<��veܾ�#�a  ��&;7'��Ǘ{#��X*���$n���Z���  
��  �HTWW�&����gLMME��"r���t:�H�3��sW����x�ֵ�T[   ����T����/���ߒ����;w޴�V�^�?�x   P��   E$�tL&����Kq�ƍ(t�����g2��/���+GN��kW���]��  y-��~�Ӿ8z�?7��R����3jkk��6l��~8   (|w  �"SYY���_~���BWQQ������E�|I&��#���k�����V���   ����x|p�r�M��������_��%A�����w_   P�   E���4�}��x��Ws��]�1�=�������x�/'��]�u+��4w   �?{����8~u �Lm'OtttDcc�=/�۷o�۶m   ���  �H%�������q�ҥ(tI����-r�+e���蕾�28ݶ.��  `������^���T@�H&�/fܞ�������[  ��"p  (r{����{/Μ9S�ᾘ����/r�+�NN�k��[��������4   �l:��g��䓶��hjjZ��%��y�X�n]   P|�   Ď;���>��|�^UU%r�k%�N�^������n�խ�w�  ������=1�J����hnn^��%[�x��&>   ���  ��{�'����w����>3>=o=kښ�lZuU�  0�Ʀf��D�ȍ�|���---������x��'���=   (^w   ��֭[s����[�{GGG���͹28��c�uMWl[�e��  p�2�l��?�^鏬���dj�b�����hhh   ���  �/ٴiS.�>|�p�O7������N�;�R��]���G��n]�u  �]]�MmO6GA>jjj����E{^ru������   �  �֬Y�����_�"��t�$rO&�_�vM�ο4<1�}x26t��}VGU��  ����MŇ�z�|�`@�J�����E{^�<x0*++   na  �J]]]��3��O��H�RQȒ�T�;�F�\��nY��숒��   �g����<�{=�*������E���СCQZZ   ��;   �TKKK<��s���/���L�$rO.p�_�.r��I�������q��k���:   ����T|p��gN�$6O ,����ػw��  � p  �k%��?����_���¾�������I��T��x�r�xܶ�#��[�e.� ���t&>���z}���W__������+V��ݻ   ���  ����:����=7�}ll,
Yr����md�sq��Z\�{7����-  ��Cq��՘N��]r��յh�۸qc<��C   ���  �o����#����(d��n2]opp0�ۘ���_��kچ㾍k���"  ��1:9�?{%����Ŏ۷n���sO   ���  ������s�=o��v�;w.
YCCC��M&�[%Ϸuep$z��b˪θsMw���  P�f��8��@��:Y�!Y&3n/))���/n���   �E�  �����Guuu;v,
Y]]]�O�;�E&���W����Pl_�26t�  PX����ǑWc:�X.��wvv.ʳ��=�X�^�:   ���  �<������|�AA��"wn���l����8�?�mX-u5  ,��������T�r��������سgO���   |Sw   ���[���Y���[��f�P%�{�J�ڵk"w������_N���ָg����p,  �Q�!�/�������f1��d�߁���6   ��p�
  �MY�vm<��3���<R�T��26Y�=00 r�;K~w����hܱ�3�X��%%  �L6'{��'W�"�)�yS�������mQ����IܞLp  �o˻I   nZkkk<��s��$����P��Ԉܙ3�t��bO��Ms_��  @��:4<%Ƨg��Ōۓ��'�|2JKK   ��;   󢾾>����_��}tt4
U�wuu�"�l��>n���t�}�\�nm��6����   ����t�����X�3n߰aC<��#   7C�  ������Mr?|�p|��Q����s�{�ȝy���h.�ټ�=��neT��  �tfә��ro��n��Z�u���eQ��}���뮻   n��  �y���~ꩧ�wމ���lPUU%rg^e?��r��Z\�>�ׯ���  ,��������K�1�J,g��'gA?�p�_�>   `>�  X;w��8r�H�$r���>�;�fr6�=u1N^�{֯���   ^�ȍ��121�ܵ����eZ�?���bŊ   ��"p  `�|��ߏ������]�xeee.rO&�g2���28>�?9+��ލk���:  ��7�������t<�,V�^QQO?���<  ��"p  `A�z뭹����_�t�0׻�'��E�̷d��GN�Ʈ��{튨��  ��%ۓ>��g�cnn.`�+))�����9�B�������D   `�	�  XpI�}�С���~�T*
Q2�L��B���ř��q��Pܾ�3��銊��   ���t&�}�'{"��S3nokk�}��Eiii   �B�  �(ZZZ�?�a����199�(��W�X����ҙl����㮵+bSW[.b   ��䃣�>���zc&U��(N��®���T��~Κ5kb�Ν   I�  ����������w����M:/D���I�I�>;;�&gS����q�Ӂ������%  �����8r�'Ƨg
I2E=9�H�\ڝw�۷o   Xhw   Ur������݉w�՝&���}߽bv�I�b�	�@�!��Lz�O�+g:�L���B;�m�b�1��}�U�kL�ɮ*=�9�|�RUI:ǖ�[�{����q���(GUUU_���'�<S�q䃳�?8��]͍  ����8������������u�{9O<�D�ٳ'   �fp  ��x��'���#�y�X[[�rs�Amhh(���6���t�z�����mۣ��6  `+��_�?}v!7�C9J;�m۶-jjj6��������  ��E�  �[f߾}������Z���D����������Ym�l�φ����Dܻ�7����jo�  ���/-�{��K�Q(��Ԑ������@�o����x��7�!   ��UN   n��6���������oY6���{OOOnt����l���x������Hܳ�'��苚�  �r�����σO_��B!�\����p{U����҂��>��   7��;   �\KKK����9����QWWWnV��WW������H������*�  ���j!N_΋<�VV�YCCC���oz���{�G}4   �Vp  �(�������x�7�̙3Q����r����X�Ͳ��'>��b(��������  P�R���K�yQ���9/����������+l��{,��   �[I�  ����3�Dwww=z4��֢ܴ���0���hY�|��/��^�v�}]��  ����<�K��޹��_Z�
��w===�nO����?�C�:   p�	�  Pt���������B�妹�9�܇���ܹ�f���ˍ��v�Ǟ��Mo  �U(�ŧ#��޹�1���U��GR�f������?�G466   w   ���ݻ�����������Qn�E㴵���PY��)~�s��ӟ������bwOG  @�I��?��?}v!���onߥ��=���6�k����O~��  @�p  �h����/~�r����r������ҥK���p+�����F�C�]���5  �|16�����[MjmO�����o�'�|2   ���  P�jjj���������ܹs�������~r_YY	�UF�g��?������mۢ��9  �V�81'>�"�f��z***���7��7oN���������   (F�   ��M�s�=G����{��B�)�?00�C�KKK����L��އ���-��=�M  7Å�x��`^|	[Qz����/7�kTUUŏ~���>   +w   JFj���#G�D�P�r�.0���CCC1?���[�<zۚcߎ����  �����>���s[Uuuu�᭮�nӾFCCC�����d!3   �M�  ��r�wFwww��W�����('W�!�����b049oL~��ͱo��;  #��ua|:�=w!�f,�ek���͋�S�}�������   �N�  ��������J���188�$��S�?]Ԟ��(CS3���Ggsc����{:  �U
�>:��bL͗עe��U=5�of�����Gy$   �T�  P�҅ߗ^z)�~��x����ܤ
��6� �b163G>8���;�bOOG^�  ߥPX�OG����y���b ��͹Y}��T齓ÇǮ]�   J��;   %��������7ߌ���('�Bw�=<<,�Nљ���ߟ�4�����z:�R� �o(��e>��Z?o�l�������6Kj���O~��[   �R#�  @�۳gOtuuſ�˿���|������*� ?�arn!����B����%� @�ri4���`�--pYjkO�a���fI���?�|^4   �H�  �����/��r���188央�.�ҥK��,Bq�YX�?|t.����w�DU��; �V��Z��/�Ʃ���R�=��7�U}߾}���   �2w   �Fj&{饗��ߎ��?�Iuu�W!���ŀb5��<s>����;�����*  (o��+q����ɷ���Z������7��>;w�   (u�   ����ƿ��o�P(D�H��s���\@1Km�)��qGog�7��  �%�������xp4V�h����&/ZO�͐B�/���6�  ��$�  @YڳgOtuuſ�˿���|��+ۙ������T@�[^Y�.ǇG���ط�/�7�� ��glf.>X?��th,
kk�muuu9�^�I;[������(   ʅ�;   e���5^~��x��Wcpp0�IgggTWW�;��z:si4�����o{_l�l  J�ŉ�8}a8ΏM�����o���<�@<��C   �F�  ���."���K�?�!���X+�f��Op###e�sQ�R(*���Ƹw{o���Ȼ  P��b�O�����brn!�����-���7��{���;w   �#w   ���{,�������B�墩�)7����j@)���ߟ�4���bܻ�'���Mj6 ��-��1>�4��_���� ���x���+�7C}}}^ȟ�   �r%�  ���gϞ���_��W��P>��uuu�m۶�t�R,--���������_���==QW�m+ �[e~i9>�.����J W'�"��766n������s�=��   �3W
  �R����W^��^{-���X[[�r��'���ᘛ�(E��+������ξ��o{o4��  7���|���p|:<�By̕�f����������
�o߾x衇   �w   ���t��/ĉ'����erO�{{{cbb"(U+�����p��8�m�q������  l�4������_��&�v���9ܞ�o����x��gs3<   l�   lY>�`�ܹ3~��_���b���R�.�����Mx��)���81�GkC}�=�w�wGuUe  pc�WV㓡����P�,,p}Z[[���;/:�hy��f��  @1p  `KK���_ƫ�����Q.������CCC���P���g�ǻ�.����ս�^� �Z��/��ǗF��9��K����My�{�����   �"w   �����x饗����q�ĉ�i=��������t�R,//���4����8}q$�ۚs�}{gk  ���gpr&N��G���Ƥ�z{{���i�_���*�z�رcG   �V%�   _z衇r ���^+�@xuuu�����c~~>�\���ŉ�<Z����;��* �����O���C1����K�������|����Ə�㨯�   ���  �/�0��/�����s(��f���������r35�<s>�=w1���̭���� �U��/��ǗFce���H��nO-����<    w   �+����ӟ�4�z��������Aggg����{��L�RC����ő�ok�A�흭 ��s��ə8�~>t~l2��������QQQ�������]�v   p��;   |�Ԝ�.0���뱲�堥�%o����M����81�G[c}�=�{z:���[a @��_Z�O.��G��1����koo�����4G��O~���  ���   |�;v�����կ~���т���144����lrn!�~�y;s>vv��]��1��  ��J[�G�#���P�Cl����������m�����SO   ���  ��H�������~;���(5559�>22sss宰����Z�o���aw�� @)Im�g��r[���b �'͛������vC_7��ӎqw�qG    �+x   p�<�/n��曱���.]T���������[Eju?��x���Z�����n����<_���������)��   PN�  ��ٳ'oO��_�*fff�����f���^(�
�� @1���F{{{tuum���޽;:��   ���:   �F�i���E����q�ԩܨX�R����@���r�V�� (����I��}�����>��q��w   pu�  �:<x0v��o��FY��S�{
��&������蛭�w��f���  �,sK��ɥ��xp4f����|���?jkk7�uSX��^����    ���;   ܀�;w��/�����cxx8J]j���������R���O>�cg�Ƕ��t��վ���"  nTZXwq|:>���c��K;�������F����{�'7�   �N�   nPjx��OǏ�'N�ZS����ϕB��B!`+Ka��c�y�&���qWwt�4 �����3C�qvh,WV�u��ۣ��kC_3��?���y�4   ���  �y衇���o�W_}5����544��CCC���@���j|48�G[c}nu���;�k�� |��ť8;<�\���� n�+��555m�린�/����   p#̬  `���_����o�ٳgK��=5ϥ����HY��a#M�-ĉO/ğ>��m�q{_W��n����  X-��c�qfh,���r��	�A������]�6JEEE8p ���    n��;   l����3��'�|G�����(eW��&''c||<��Ka���y��:��o�����  ��t^0<=g������X.� ����������܍�Z����hii	   `c�  �&��;r��������h������p7<<�B!���������X��t�}]�T�q� @�]\�O�����ј^X���׺��6�5w��O=�T    K�   6Qj����~G����{/7:������O!���� ����B����x��`����ή����� ����872��ڇ�f(NWv%KM����*:�v�
   `㹚   7����s�[js_\,�Fǚ��r���� �[Z�ra|*�ʊ��������TU P:�n-�Ǧr����T
����]]]]����y�F���^x!�p   lw   �IRc�/��x������Q�***���),���B!�������&󨪬���)쾫�=��? ��������L|24�G'��s�����DOOO��n��:�����?�A    �K�   n��5zjz;u�T��(�`xsss����R W/�宄ݏ~R;����z��ܘ p}R����t|6:�F�ce����a+I��lO�ՍR__�>�l^�   l>w   ����;w�W_}5�����������ctt4fgg�vK+�q��h���v��Ѳa�� �w[[[����8;4�����@i�������|�(�v�Ç��<   ps�  �-��K���G����{/jJՕ�����t/�n���7��Ʈ��������@	 \v%�~nd">��� JS�cwwwoX���:~���m��   ��%�   �������;�����_�7��-�SS���P�����[\�.��R_�����jn�� ש��C�3qnt"ΏN���r �+�wuuE[[ۆ�fooo��G?��&x   ��	�  @����m����⣏>*�� ضm[nr/��>���x���<�j�c{g[���-Q)� �i����q~l2>���e���&���7,����}�Ѹ��   �u�  �H���{�'~�����B�������D]]]����t`����J��4�G
����Ďζ���5UU D�����L|6:��L���j 壩�)7����FHϟ��<�   n-w   (2}}}��+�ěo�gϞ-�pxkkk�ʊ�L�)����xU��1���])���5��`kI���s#qa�XX���MEEEtuuE[[ۆ�^
�?��ñw��    ��+\   P���g�y&>�����oKKKQ�R�}۶m9�>??��Y-���d�|�y��6Ů������u� �hvq)>��/�����v�v(_���yQx}}���^sssnmOG   �x�  @۹sgnsO!��>�,JU
����DLNN�t+=����lhr&�cg�����꾳�-Z6& ����\^Е���Q�V������y~y�R�<>�`    �G�   �\j�{��⣏>������������=r�{)�PjR�}xj6��g�����ho]-���-��n<$ �i�P��RK�����[Z`kHa����hkkې�KA������   @qp  �q�]w��ݻ��^�K�.�lz]]]l۶-FGGcvv6��ofa)>ɣ��2z[�r�}Ww{4�� ���Ÿ81_�MŅ�(������ڼX:ި������'�   ��	�  @	I�_z�8y�d���g
�(EiK������>66V�?�����)<��Ϝ�������;�ڣ��9*+* n���ZM����ߤ�G'cj~!��+5��yc������Ǐ~�����   ��	�  @	ڷo_n�����܄^����s�`xx8��R[��󨮪��������;Z�Q�; lay%�������ӱ����VUU�����ظ!��cǎx���Bk   �4�  @�J���������ĉ�������:bbb"�x��r�0�Ԝ��ܘ��;:��o7lH�& [K���ӳ���ߖ/ƧbrNK;���._)ܞ�7*���SO��&   PZ�  ��=��Cq��w�o~�nsooo�m�###���@qI�hF�g�x����������-1��]-Ӱ	@�I��\���cp},�hi�.-�Ls����y��۷km  �&�   e���9�����{q�رX]-��P
��v�ԟ���x�v�+a�q!jk���9�[b[Gk4�� [���rO����}n�c�oSSS�[��|�F��l���	   �t	�  @�������_���RTUU�����166�[������4���{-Q[�H�r���#�s�����T�����hii����iZ��;�����   e�U%   (3��^�ӧO��o�+++Q�R�!�,��ñ��@i�YX��������ln�����oo����\��ҴZ(���l�M������_,J��;�;R=�Ӽ�F566Ə~�����   �<�  @���{bϞ=��o�_|Q�M�i��������� JS��3:=�������2��Zrؽ��):���X
��L����l\����X-�޹%P��ꢯ�/��nD
��ݻ7~��    ʋ�;   �����x���O?�#G��dzn~���m�###Q((m+��8?6�G��͍����U轪�2 �5���ٹ�����}6��܈4�kooߐ���������i�   ���;   l��v[�ڵ+�|��8{�lI���m�o����177@�HA��L#5��6����ii�z�h��� `s,,��]6��f���ͭ� %�������7"��?��Cq���   P��  `�HA�g�y&���_����(5UUU9133ccc�ܡL�Pe
Z�����|_s}]�v����[Mu����_Z���hj&��g��[�����]]]yNz��������   �O�   �����x�W�w��]|��Q��v�)�022R�A}���,,�G�i��[��r�=�����(�𷤝{&��
�M����R l�������ɻq݈������;�3   ��A�   ��Ԝw�СػwonsO��&�%RXzz:�����uL/,��ɥ��qMUUt47DgSC��6G_{K��x��zR;���|��\nfO��+p3�E����9�~#�^�=�\��   [�w   `K��_��q���x��J2$����U����b [�����v������|_cmMt67FWKc��6�������r��Z��ٹd��_�83�ف['�Sk{SS��N
�?���gϞ    �w    ���w�uW��7�����(5555100��������$sK�176��.�^����ֆ��ji�M�)������P�
��7��1:���=5�;��Ecccn\����ݻw��*-L  �-K�   �����������s���;�������-r��Ғ�R��Rtrn!�3_�WSU����Ҕ�񽥾. n���jza1�G�fcd�r�}�P�b���]]]���zC���O=�Tn�   �6w   �k����~�ȑ8{�lɵ�����6���>55ZM�ﲼ��&g�"��[뢭�᫦�|��"
l�o6��������Uav���Pz
�WW_�e����������    p   �J
'<��3188o��F���E)��������Hm����p�R�}tz.�+M��W�j���>޻��r�{CmM \��啘�_ȿ_R�=ڧ�-�JN�suvv��nDj~��g���>    �p   �U���+q�ĉ�ӟ����QJ���b۶m1>>����WjX�YX�����W�7��D[c}]-M����u9�l])�>���s��}�򢙙��_��(})����55׿�/�՞x�رcG    |��;   �w=���q�}��믿�[�Kɕf�������� �(sK�y\��^�h8�W]Um���P�U�=}�\_������L�/���|nb���|�\?����e#Z��k�~�����Geee    �-�   �UI-}/��R|��gq�ȑX\\�R��۷o��������Ͳ�Z����<�ReeE4��F{c}�75\�7����������A������[�;:��ف�`#Z�[[[��g�����    �.�   �5ٽ{w�򗿌w�y'N�:kk��Jm����###��� 7K����i���B��ښ��ޯ��;֏5UU�<K++1=��C�s1�����t��QR�z�C�Hk{uuu8p ��    ��   �5K!��ƾ}����_����(%uuu�m۶�䞆�p��--�qqb�k���TGs}�������߷/�k���3Ky��t^tr���# ����===9�~�v��O?�t�C   \-w   ລ�����ş����農��"�����H��E�6��� n��s�����c�u�_��S����1��������斖�
�� ����'L�-���j ��R���+Z[[��5�<멧��y   �k%�   ܰ��/o7�ȑ8{�lI5�������@nr���m�@�(�����2������ʊh������M��9��T[�o7��)U�)����w=�M����ا�����\�������������~<�@    \/w   `C� �3�<�������6fgg�����}�澰� �,5X��oߦ��:��Gcm�W�)������6��fJ7ҮWB�)����q
�ϯ�N��P� ;�ƪ���m�)�~�����駟΋�   n��;   ��R���_���?�=+++Q*jjj��?==���Q(�\�q�siQ��_}���"R �.�kr���.ꫫr8>�S@�^<W!��/,_����������]LA���ʞ���jii����r�i���Ç���7    6��;   �)�����{�ȑ#q��ْjZM������>?? [Q���ڳ�����������h���������>௄��ǵ�I�Uė�Z�_Z��F�W
�ǥ���K���_������ (*i�ojmOs��������   ��$�   l����x�gr#�o����Q*��������9���ۭR��pU!����Z�k�*s�&�禀|uUU>��k�/�_[U���iԬm����K+��c%ԗV�o�p�j�?���r`==���Ws��PB�� �������^YYy��M�v������   �=�   ��K��?��O�̙3��[o���B������������v�ƤP�\j����W�O����c��J𽺲2��t_���]ݗ��5_�_��c��</=��2��ؤ0���JnL_Y-��k��j��K���5O�IǕ��Ǥ�.�ϥ�/����W�})��b���SWW�[���Z���in�1���   �fp   n��o�=�'Nğ���X]]�RPUU�C )̑�ܗ��~C1 �#��WV�n��K�o�������7�V��W]��-���_o:_K��o�˯�`3���J����A�kU[[��n�-    6��;   p�=���q�}�śo��ϟ�R��ܷm����y��" �mq��C� �#�J������~i8���8p�@�   p3�   �D
����122���Q
R�a{{{�������|   ����loll���yO���駟�s7   ��I�   ��R�����ԩSq���X^^�R��"}}}177���  p��pzkkktvv^W�z
�>|8z{{   �Vp   ��޽{��{����w��G���Z���H�����155   �JCCC^D\[[{�ϭ���Gy$��    ���  ����:>�`���1<<� }ߩ���9FFFbii)   n����<'I���*5��ڵ+�Ů��   `�	�   E���%~�ӟ�g�}����cnn.JAjIܶm[LOO���Xɴ�  �+͟���r��Z�����Ç���)    ���;   P�v�ޝ�ɓ'�رc���� Ls�}vv6   6Z]]]twwG}}�5?7�>��OD___    w   ���۷/��ݛC���_��B!�]jOLm�)�>::Z2�|  ��UVVF[[[tttDEE�5=7�:�����w�    �J�   (	)ı�����������Ν����(v�Mq۶m199�G)|�  @qJ��]]]Q]}m�y��{�7y�    (v�   @II���=�\LOO���K��>4�Z���se||<fgg  �j���Ewww^@{�v���ʋ�   J��;   P�ZZZ⥗^��/Ƒ#Gr�إ�Ş����������R   |�Լ���mmm������8|�p466   @)p   J���@���?��?�8���?���B�Ժ�m۶����A�B�   W�]�������r���=��S9   P��  ��p�w�q������+++Q욛�s����d   ����������������k׮    (e�   @Yٷo_�{���[o�G}kkkQ�*++s�b
��6����   ������؞دEMMM<��Cy   P�  ����!�����Ĺs�>�B)}}}177����@  ܸ�赭�-/|�������ٳ'��|   �\�   e���>�{��#G���x�kll������������  �/����Օ�^��ߵkW����   @�p   �^www��?�c�����b�+�����ԔC����  �����<OI�r�Eoooޭ*�    ʕ�;   �e�0��~������㭷��-�Ŭ��*zzzr�=�򗖖  (]�?5����\���\��'�̍�    �N�   �rv��?�����O?�w�y����q۶m��}||<VVV  (���y�jGGG�}5��N���9؞�   �U�   [�m�ݖ��ӧ��ѣ���Ŭ��)s bb"
�B   �-��wvvFu��_�M��'�x"?   `�p   ��{�'��'O����cii)�UjqL͏���199SSS���  @qI�S�����������Ӣ��<   `�p   �Ҿ}��HA�cǎ���r������� ���cvv6  �[���.7�����J�ݿ�a
   `�p   ��r߻wo������j�������ɭ�)辰�  �͗�������ժ���Ğ={   ���   ��Ԑ�~�����������������n� �r��)����W�����x����{�    �N�   �;\	����[o��q
�(V�}����������� @�kii���Ψ���������~���c    ��;   �U����C�Ł�w��]�;w����)h���SSS9辶�  ��hjj���X��q<�@    |7w   �kP__�>�l,//��o�]ԍ���֖�����133  ��K󁮮���������������   ��p   ���15�?��cq�ر8}�t���F1�������vOm�  \�T������W����_�   �:�   ܀\9x�`�߿?�=~�a���D1J��������sss  |�t���y�������#�ĝw�    \w   �P]]���>�hnt?u�T��S(���7s�}~~>  �������ۣ�������?�p�q�   ��p   �@�����=�[�}��8y�d,--E1�������t����  ��,�ӎG)�^QQ�M�ohhȍ��~{    �1�   6A
�?���y����'�:���ߟ��SнX�O  �,��=5��p��ۛ�����;v    K�   `��۷/�ӧOǱc�r�����4���bbbB� �����)ԞF����f�G}4�o�    lw   ���{��#�S����l����<����WVV  �IjaO���������---q���    6��;   �M��A��Ǐ���b����U�=5�� P�RX=���`{UU��}lWWW<������    ��    �ȕ����~��crr2�M
�477����t�WWW  Jɵ�SS{jlO��    �\�    ��m�ݖ���x���;q�X[[�br%�>� (W�c��ڢ���/�VVVƮ]�������    ��p   (��/���\��f�B���/�� (V���^SSw�qG8p ��   ���   �Lccc<��ӱ��ǎ�?���B�W��i\	�///  �J)�~%�����������   ��!�   P�jkk�����裏ƩS���ɓ9L^lR�{�y>�S0  n�fokk�㻂�i�fKKK�߿?v��    w   �"�:������ٳ��}rr2�Mj�LC� �����*7�_M����3~���#    �K�   ���ٳ'�������������(&W�����9辸�  ��R��Jc{
�������lO�   P��   JP����?cjj*�y�8�|
�(&y,,,�{: �����Ρ����]����;�3y�|   ����   ���=�=�\����ٳgcuu5�I}}}�� p�jjj���=����3؞X����o߾    �4	�   ��"?|�p<��q�ԩ<�����\	�/--���d���  |����������;���?�p�ر#    (m�    e���2�U�q���8~�x\�t)��֢X���FOOO!�~�B!  �����hkkˍ��&��n߾=8�w�    �w   �2500/��b���űc��̙3���Ţ��:��Spiff&�����  [SEEE455E{{{^�m�����x衇r�   ��"�   P�R��O>?���ԩSq��ɘ���b�BI����u3}_)込�  l�|0����i�I�#S�}�Ν   @�p   �"Rph߾}y\�x1�?�.]����(�����9��:��� @y����S��ۚ���۷o��<    �O�   `�_|1ɏ;gΜ����(�u>�p���*��y  nLmmm����i��=���΍��~   �<	�   la)D��O���8u�T�<y����uuu���9�>==]4��  \����hoo���&���P�Ν;   ��I�   �܊�o߾<.^�Ǐ�K�.M����::;;s�畠{�P  �[jhojj��������s��۷ǁ���%    ���   �����x��cnn.�;gϞ����(UUU��3�R�|
�/--  �%����zkkk^����F�;�37���;    $� �����X]]��}��t��jjj�   nLccc<��y�9s&�}���b��@����H�tO�w  n����lO#��}S
�www�������'    ����TW�&i����Z Ә����15B.,,��z�/��7"rR>]TI�ߦ�{���O����k��I�Bi�0��,  [��ߞG1���s��������<�(
 �͑�������jz��o��   �Ւ�ຬ�����dno�����������P����-�>S�&I!��q�L
���LGGGy;�� `�(�V������=���r�{1�I  �Y:�J�P�VY��v    ���; �*5������p}uL#��WVV��]i���Ǥ�tq&����<��N�  (W���D�B�4��*��  l���N
���ν�I[;    7B��dO��.�ŋ�1���b�Q�����Mi;ށ��ضm[>^�  �E1����UZ������N)��@  \���ޝ@g]������$d���"��	�E�E�}��V��ڱ�e��z�̙qڞZ���.ETv
HQED�N�	KH H��^�FDH����ޯs�yB�&3��w���ύ��wm��y.��     �-� �TVV���ڵk����ݰ`�W_}%x߉'\��FU�d��֭[�ѪU+5mڔ6#   �@mu���t7,%%%�6w�3  �8{���v�ׯ�ݭE��  ��a�V�gE���io[�r	gΜ9��<�_�=�۳{UVb���_��3tt�  �7� �lc-�(��u^^�kg����l��}�v7<l�زeK�i����  �`U��ݞ{7l���JHHp��ɓ.�na��@   ���Â���n�PUY8�
<z�꥔�   �O	Gii��=�n��[���x^-�^Wl}��U_=�JDl�`���� �[�@�ӹ۶ms�O��އ�`�sC�6�ݭ)33�I!   �N�v�ܰ֠��׻g^���7;dڸqcw�>�<��  �3�[���%���h�;u��m�   ��ٍ�TQQ�>|vX����׆'`_\\\�����d`mX����4�k!x  ���; 1�[;{nn������$5c'�?��37�m*edd���m"�kTT�   �``ϳ�{�v�6w֭[��{��kt���Y��!;xj�I6hu  ���y������۶�تU+��?Pll�    ȕf�����ڰP��9r$,���ކeW������.��ym֬��6m�� ���; ;�kA�/��҅����#���$=-�,P���]��ݳ���Fӹ�   ��Q�F>|�{�n�ڸq���{�c�.�,D�;  ejk�߳�^�z�I�&   �WZp�����s�v������q׮]n�+99مݛ7o�^[�hᆭ� �w p�w�>h�p����0o޼ٍY�f�)�gee�K�..�   ��mۺa����tZ�ܟhu  ��Bm����;�5F{   ��[��ؖ��f÷��ކec<lNbn�{V�g���  �>� `<-�6lp��C�	�.�Y��c'��u��6�lc�M)   ���(���ۍ��b7/�$���  ��kk�P�=�dff���/Wll�   �pa�j���矽I�u��a<������ۼ�}����֭[��L���  �� ��#,���矻ӨL��-��ނ\�R׮]]����-<   ���4:Խm!w��M��  ��kk��Gzz�z��ƍ   u���w�^mٲE[�n�Ν;]����ѣ���O�0�}�vw�_v�e�5..N ��F� ��B�_|�{����J�d��V�X�M�սW�^43   �y�����6�({������ǏwAw�*  ����			.�~nɅ=�dee��  �Pf�vkf��D۶ms�x=v���������e˖.�ޡC�j7Z �w �Cv�w͚5.�n��i�����0m�&Wvv�ٰ��t   �@�ZFm��jݺuڳg�_o����٨��PYY����   u���4h��~��Ђ�ڵs�:��   �������{vhOv�a׮]n,^��͗����Z���`0  �� |�&L"�P�ƍ݃4H,�~�z7<�����S��ݙ�   `%''k�С�m۸������'O����d��IIInX���ݭٝ��  �W�fF�a;;xW������֭��   ������Kw룽8���Z��kx��?�[`׮]���. @�!� >`M}j_�z���܇`Q��ݚ�z�쩾}��}���T3   �5jt6�~���<�o�>���,Tf#55�|�Vw�  \*+��@{bb�ق
[���7o���vc�   �Pd!v������@M����ؘ>}�[_���6hw���wc �"P�Z�J+V�p� �Y������HIIQ�>}4x�`���	   TM�4�����ۻw�v�M���Wee�_>���Q��f��6_d�  Ԅ��[������ξ�B�-Z�p�1�   �v�ڥu����>s�����%K��a�Ν;�2�.]�(::Z  � � �Ȯ���v��ٳG@(:|����kѢE�ԩ�����/����   hn�[��5�ە��`��֦j�Z�,�ns�ӧO  �|,�nm�6<7,�3Ezz����>    Y���O?�'�|���`�qڿ9v����z�r󯪇� �G* j)??�5[[c��S���X�;�l�aÆ�Y�f   �'�nϴ[�n��͛]3����111nXӪ�m�8qB   �hM�j���t��ڻv��Z   BV^^�>��cl?r� �,���ذ9Yvv�~���2@[� �w ����rwJ�>��a�N.�!�?�PYYY4h���y6�   �@T�^=u���O���/�t��#�nM��VV�|�9��;  �ǚ=�����;סC��   ����b�Y�F}�M�Xg��f�~���fw� ��� P���ג%K�z�jr���溑���������L   ��j�����r��URR◰�}>�`[ee�������ɓ  ��B���n��ƺ�YyD�F�\��]�v   Bѱc�\S�e0�������6��V�+��Bmڴ �{��l۶M,���k�`b�Ľ�3g���>\-[�   袣��3�O���͛UTT������Шk�4�v  ���x;�V5�nA���t�o�^m۶   �l�mӦM����׻5/ �ٚ�e��hڴ�������6 ��p�sXkߪU�\c{AA� Ԝ-F�ב���,6L]�vUDD�   �@W�������e�wE�?6�,�f"6��ۦ�5�[S  |�lѠAl�W[#���7V�ΝբE   ����>��C��~��Q�j����9s�f͚�.]�h���֭�� j��; �����裏\c;�*�{��k�2d����JEEE	   ��`M��6�ݻw��[ۘ�G���ᒒ�ܰ���naw�  ,UC�qqq.�n7�4o�\ݻwWJJ�   �Pe�7ntł�����6lp��q�����+--M ��#� 암����/^�'N�oj���?��_}��ns   &n{���/��_��OZH�Frr��[�����J ��g�v[���n��Z�r����   eV&h�|��:t萀pg_V��p�BeeeiРA�ѣ�� P��-k۳���L�P��P��ٳ�t�R:TW]u�{   JvK�cϹv���w��u�J�Fjj��fw��:uJ  �w<M�e����H%&&�P�]I+    �mݺյ���g�����zqnn�M�4q9�+��­� Ώ�;��STT��}�+��,lcA�E�i�����԰aC   �ȞemC�Fii�>��s�޽[ǎ��ϥj�����ݭ�  \����0{�P{JJ�ڵk��h�  @8�u��������v��! �c��S�L�;Ｃ����ꫯVZZ�  �F�@� �&��i~��$�  �P���p6�n�Ok�ڶm�����Q�x�|m�6O�8���
  ��~�Z�݆��GEE�q��j߾�233	�   lX��|�e˖�[�Nyy��J����_��vp �5� B^aa���}}��'u~E<��t�븮��w�3   �,�ֱcG7����]�}�޽�U�.Y0/11��[��vg� �wY���Y�ݮ��ז-[�K�.��   @89t萻���s�)�[�]�v�p���kյkWEDD �w !ˮ�����ŋ]K��`�!����?��O:TÇw�X   @(hڴ�櫯�Җ-[�ζAXYYYg���-�g���r����r�  ��:Tզ���T0���hi  @X�R��K���[��om߾]/���Z�h�J{����H@8"� �؆��\t]_��{�ky����j;�6�5N   �"::�5��0�����w=m]��[�ݞd�>�}lO�;�� �Pg����8�s�B�v��y�����v�v    \���kΜ9ڰa��u�n ����{������O^@����aavkk�?�ۄ�6��3gj���=z�z���U\   IU��-dna���<>|�N���a,�naw�9 
,`av�/��m�ֵ��4    ��ٳGs���ڵk	�~V\\�I�&��I+���+% �=�P����EEE�<�q��)33S��r�ڷo/    T��ƺÝ6N�>�;vh۶m����������6t���v�܆�+++ @0�\����Ҟ����eee�q��   @�dV�2}�t-Z���;��A�@P۹s��~�mm߾] 5X���U�n�t�m��Q�F   BY�z��O�!OkR���]m>v�Y]�p���6--��=�w�� ��iٍ$�s�j�Ϯ֭[��   �Â����6l�  ��j�}Ĉ�߿�[?�PD�@P��3f��� -����jذa����#    Xm�.]�0��a�wی<r�k|��a-��1������  @UU[����բEu����   ��Y�b޼y�裏X����	���[�օ뮻Nt% J�*Z�l�;=|��Io�T9�|�Z�J7�t����ˤ   a'%%E�{�v��߿_[�nUAA�JKK��Jik	��`BB���5�{��� ��ii��Av�_��͕��ō   �;v̵?/^��e0 /;�2q�D-Y��5����K *���<m�4	 ���ʜ�}�ᇺ���ղeK   �iӦnk��������u��A<����5�ڰ�}r���}|� �ڲUh�a7��P�6mԶm[   �0[����\㳭� ����+���}�|����� ;� ^aa��N��/��B p!�R���k���5j���   -��	����m۔����}���ׁ��aDSYY���w��  ��n�S�3$99�m�[����.s?_    \����^�Z3g��ѣG tmڴ�e&z��1c�(--M ��X��m���}�]�� T��C.]�T�~�������O    �f!�.]��a�6$;(ZPP��>u��?���H��ǻa,��	�۰gz @����9hoѢ�Z�j�v��)::Z    j&77W3f�О={ <ء�K|���:t����z�. ���;��dmr�&MrW� @m���(''G�|���NN&   �a��޽{������6=:��V�~}%&&�a쐻���^}�0 �/�9РA%%%�u��n�iӆ@;   p	
5m�4mܸQ ��W_}��F��>}����  XpP�������]+V�`�Wآ���iĈ��꫹�   ��sޭM=//O���:x�JKK}>_��^t��o!wϰM�  �EEE��������왙���    ^�	�ڨ��� >����^Ӓ%Kt�w�98 � �]�3q�D�` �d�vx�N&�;�m�   �8�m��c��{�����\ི�ҧ�Z}m����݆}N ��e�v�>n�v�D�ܹ��4i"    ޵a�M�:U����sٚ���g���W7�|��5 Pp�wǏ�̙3�|�r�/�ٳ�Mج��G?���   @�Y�<##��4ݱc�{�>v�***|���
]k��a�ƚ�,�~��	x�e� pa�}:::�m�7j�ȵ�ggg�aÆ   ������ɓ�y�f��X�ȪU�\	�1cԿ7��@D��_}�駚2e�� ��`a���&l����[   ��IKKs�w���ׇ�Ν;����f�s_� �'Li,`�iw��u� �;v�)..�؛5k�:�P�D   �[�����C���O ����2���Z�b���_�E͛7 � ���&N���k�
 �a߾}��_��믿^7�p�ې   p�RSSݨ���z?x�JJJ\뺯�MM			n���w���c@�������n��ܹ��6m*    uk�֭�4i�


 ��m�6������o�Q111�@A�@��k�rrrt��a�?�>}Z�g��ƍ����L���   �}~������]������� �������<�B�6,�n��w �.+�&���$�fҩS'7(	    ���P�O��իW�̙3�Ke�A,Y���&��=++K ��3�@4w�\͙3���������\7�|�$    �e��mۺ�QZZ��{��ё#Gt��q��x�6<l��v�໵�[ �EDD�����a���4]v�e�޽����    0lذ���ۺ	 x[aa��~�i���W��v�4h  �'� �]E>a��� ��,'Nԗ_~����]�   ��X��s��n��z���<�cǎ� �/DFF����6�(o�O��^9� TDEE����n�Zݺuso   <�&2c��Z�J �K��i�krss]��~ !�����g���>ۄ oZ�v�v�ܩ�����С�    ��5�7o�܍�����{�n8p�5�Y�ؽ�Z�-to��控��z?u�  �U�gdd(;;[͚5   ���駟jʔ).� u��ѣz��իW/t� �?p�36�z뭷�~�z@09|���|�I:Tcƌq�    �������j�޽ڷo�:��Ǐ{=|���X7<�e�>�O�݆� �}����vs5j���Lw+FJJ�    [ۘ4i�֬Y# �;d�}�v�s�=��� �%�Z |®�y���]� #kg\�d�����g?S�&M    0Y��cǎnxTTT���@{�����]�B����-�2ㆧ���-��	�۫/Z��/��cn���\{۶mթS'p   �v�ء	&���H �o��z��)P��n��l������zs� �%??_�?��n��v���_    ��m�ddd��a��v߽{�{���N�8���}l4����4�[�݆�[�����(w��^a���0O�-\c;   ��aks���ܹs�@@�nڴI��{�[�  _#��klSx���ڼy�  �X��7�p����.��    �X���t�Mָn�h���w�G�uW����u��Ӷl��6�-�n�w{�: �k_�� ���q��.�ޡC�o�   �l=�Zۭ� վ}���?�I7�t����*��)� �b۶mz�W�0 ��U�V�	�����Z�    �k[oڴ��*..v����B��QZZ���`����7��P�'�n!{O �^�1n��k�ݰ7�[�V�v��   a�� 'O��J�  ��:������_h�ر�> �w �l���:u��p�P�k�.������v�S�N   ��p��Ν;��t߻w��>|�l��W�[ ֚�m��j��3��qx�� ���SRRԼys�m�V�Z��f8    ��%���Z�~�  �X������]Ƚk׮ o#���l�N�X�B Nl���g�Ս7ިk���k�   �0�����;�Q��,�n�����Ǐ�u�_j����8�߫��W}���O�=>>޵��a���teff�fv�}    8�M�6)''GG� �cǎ�^���u뭷��� j��;�Z���q��iϞ=�pd���3gj����{'    ��kj>�5�:tȅ���ą����]�R������&6����s#pa���ns֚���m�7m��5�[3��>    T���g͚��r @H��e˗/�Ν;����� o ���6nܨ	&�X wve����'����q    �>��`��s����UTT����~d��'O����e���>��B��f;B�}}DEE��!��n�u��l����ccc    �`��W_}U����Pc%��?��~򓟨G��KE�@�ن��"~�w�܄۔oԨ���PPP  �8p@��_4v�X���S    PS��P�����n��eeeg��{���ǵ9��]�	�WVV������ EDD��u;�a�boذ�[�JMMu-��j    |i׮]z��ݼ B��T9n�8]s�5�����# �w �b����nM�-��g-U6�m��ܳ�mo{ެ�*>>�]�nv%�m�m޼YS�L�l���+��nЈ#�   �Uj��E���O��B!x��m6���]Y˺�m��q��JKKs�����   ���Z�J'Nt��@��u�(//O��w��@mppQ�!����+??_��gmT�a|���m���_l��:��k6Q�={���ۧ{��+_c    P]�	�;v̅�m?~܍'N� �'o�tS�P�5d۸�oYӻ��=�j;����~|�Oh݊<ֺ�Y�JIIQzz������	�   d6ǝ:u��/_. 7V��������Wff� ���� iZ��k����/��2eeei���:x�ڴi�m���&�m,�ƣM�|m�ڵ:|��~�_�w    ֘d�u�����F��G�����-o���	�_,ok�	�{T�����@`��ok��a�vd��ຕ/Xh݆�-Y�zrr�{��j    ���
Ǎ��;w
 }/|�'t�wh���� ��{mڴ�M�l���6 -�n�m۶n��t���/��m:������P �a�Uv��P�V�    ��:�����._ZZ�֒��6,_�ޮc�\7���$_��{� �������'$�ayO(�^=o��<A���m�ʚ��՚���ڍ���+    [�l����URR" w���o�����Z�j���Z�b�&N�ȕ��6-�ޭ[7l���/5jԈ�;pG�����7����:w�,    U���n4iҤ��[�����`��Z(�jS���m#�jx�s���V�Wf_���ws����x�/��<�s�����ϳn����������{�����������R���Ն5�[P    pq6�[�d�f̘!n?�y���z�ܹs�T �-_�\�v������. �b���p͞=���m@�o�^]�vUǎ]V���;�����^w�y�$    ��Y�ښ�mx���[���������m��y���sٟ;7�na�s� �6�{�/�n!����?�	�WekD>��������~�8�W�D�߳p:    ��ٜ��W�^-��ۺ��=��ږӰ���ڼ�s���y{�� ���IOO'�����|����/~�eff
 .��;���p���4j�ѣ��7v}�>g ���&Mr��#G�    ��<��6     �b�_z�%mٲE<�g�ԩ�Z�h�iӦ��zFF�Z�n��V藒����Di ���G��'�Џ�c���G �}�p�p��M����ճgO�j�J��q��pa�2:�������         EEEz���~!p4i�ą�m����k��^5k�̧a��!�|۩S���k����1b�yoD � \��g�a�����.�ޫW��^Y�l2f��^��V�X���2�w�}罢         @�۹s�^x�;vL𿤤$h�޽����2-[��?X�<�o�Z�}�ر�' |w ���'�t��Q7l�ԦMj��U(�8[}bb�JJJ��֯_�g�}V<��bcc          x�[�ε��W��X�`�Νխ[7eddl��)��O>q��_�򗊏� xp5�?��S:r��{vҰG��ׯ�kn5��N���-[����>� �4          H,^�Xo��6ae?����٭�݂����l��6�ѣG�v�ء����.?��* �C�S�w��3�<�UYu����{�V�>}ԠA�*��'�������O?�_��WJHH         ��t��iM�6M|��P��Vy����3(��� �|������ֿ�ۿ�C, @�C�|��gUVV&�NJJ��&X�pb�R�d@��ڵKO<�z�!%''         @`9y�^}�UmذA�[�Z�R߾}թS'իWO��2۷o��g�@,?���\�����af�֭z���U^^.����=z�䪦��g'���~��%          �Xy�3�<���|�nԯ__�;wV���դI����4�8˴������{]�
@�"����7��_֩S���`��\���o������         �����p��={�kذ�kk�ի�bccJ�T �WQQ�W^yEw�}�;� <p������~{ �w%''k�С�ڵkX�=�fP;�rM�=��Z�h!          �a{wO=��
߲v�>}��`����"�@͜>}Zo����!Y.@�	�' ����+''�����4h����ׯ_�N�j"""�M����+ �g-O<�|�A�i�F          �ݾl�v{��n�ZT���]� �Q�ܙ3g4m�4W�:|�p/$2��z�jn����pX���+�Ptt���w?~�]u����E          uc���.�~���7Z�j��:tP�� �5��۷O ��2o3f�бc�4z�h܁��g����_'��%6��֭�;��� |�M� xǉ'��s��7����5k&          ��{�nWDeAJx�ۇ��m�*Yi w�v,X�2pr� |��;�rss5~�x�>}Z�t������kմiS���d������O?����w|}         >����g�}Veee�wY�}ذaa{5{���Y�p����u�wr� w m߾]/���***�K����k��F�:u.�q���]v�����7�����         ��nݪ��'�=�!�����l¨���^�����t߫��իWO Bw ��ܹӝ(>y�P{����ݻ����*EGGՓ����9 �C��mroذ�          x�ƍ���/�ԩS�w$%%��+�T�=�VA�;����&���?u/ ���;B��٣�{�ŗ(33S7�pm�`��z_\\, �UXX�B���o/          �fӦM�۽�
��﯁�~}bi�wJ�X�f��Z���8H�(�$�q��=��3*++j'11Q�^{�:w�,Ԟ�8&���޽{��SO�׿��4h           ��c���⋄۽ ""Bݺu���Õ�� ����������p�֮]�7�|Scǎu߇ ��@8x�|�I����c�vkm'0z�,�y�f��ݻw���ׯ~�+���         @�؞�s�=��'O
��u�֮L�Y�f��Y���;�=+W�Tll�n��v-܁ g�O?���9"�\rr�F��v��	�a�1 ��}�v���Kz��%          ճo�>wk���ǅڳ�aÆ�gϞ4'�@ZZ��n�* ޳t�REFF�[n��A�b����DqQQ�P36��ӧ��lEGG�C���������}��ǂ         P����D���L�ۛ�֭�~����;j�L����?����뮻N Bw HUVV��_�޽{��IJJҍ7ި6m��׸qc��~�������4          �����.�~��Q�vZ�h�n�A͛7j��;�;�f�rM��\s� ?�@:s��z�-�ދ��ܹ�F����8�7bcc݉���R�y��)99YC�         ��*))�SO=���b�梢�4x�`���_���j��;�[3g�t٥+��R �w ͞=[+W���\���zwM|�&d܁�3m�4����=         8��]?��:p��Ps�Z�ҏ~�#��^b���a)// ���ɓ'���>}�@�"��O>�Ds���/33S�G�VÆ��aۼ�<��O�ք	����N-[�          ����z��UPP �LLL���^�z)""B��T�ٳG |�B�999��X��� 8p��֭[��믻¸8�ˮ���Yu+--M ꖝ�����#�(%%E         @8����+���ݻw5�����n���"�Lw���(p���z��ծ];>܁ a��_|�EUTTgW:�d���j2�?�9�g�}V�������8         �Ȋ�z�-���
��A�Q$�cd*��q��)��������t.܁ PZZ�~���Y�����k���jР���7 �طo�^}�U=��,:         ,͞=[+W���V$جY3���u�rwVh!���D܁ g'�^x�
�誫�"��gIII���r�~Խ�7jҤI���         ��O>�Ds���ǲ}����W_�������@�:x�ƍ��z��s@�`veք	�c���bbbt�7�S�N���8--M��� ����]��-D         �`�֭z���]���#G�s��B�IMMuō�O���a?rrrt���\��G�`���Ӻu�kڴ�n��V7@�����1c��٥K         ����@/���***��kѢ�n��f���u+22R���:t� ԝ5k�(==]�F���G�P�6m���/\X�4f�����Z��yny��G�$         E���.�~��q�¬�x���:t�k�X���;P��Ν��\y������X�Ǐ�*��	׀4l�0��	P܁�`�x����#��+        �Pr��)���*,,.����8;;[�/�TlٲE ��ԩSոqcu��I w ���kܸq�t1ί~��9r��w�..�@��srrt���s(         !�s��;��=��n�ͅ:�d* ������/�����wjٲ� &�@��<y�����KHH�wܡ-Z�---�imA��}��g�?����:         ���w�Ѻu��ڵ�+����e* �Oyy�^|�E=��JLL��C� ˖-ӊ+��KMM�]w��^��������Ç@`x��w����5[         zV�p�B��Y)����5d�!����_qq�^z�%��׿V��Di�@�W% 캬�ӧ痑���4h ��p���?��� 
         �8���n� kk=z�������20Ǐ �پ}�f̘��o�] w  ����W^QEE��]��ٺ馛\#8��ܷn�* ��رc7n�~���*22R         @09y�k�-//�/))Ʌ5�5k&���4�@ X�t�Z�l��
@� ����ӧ5~�xZ��G߾}u�׺k�|�RLvkȻ��         �`a����


��kժ��[;8�e*v��- �7y�d5m�T�۷��@��Y�fi˖-�w٩����Z^v�@`Z�p���u��M         @0X�`�֮]+�_vv�n��&EEE	��L8*++]I���G%&&
��p�h�֭Z�h��m��~�5��+���@�v���=��cJMM         �6m��n)�����O?��]���LX�9�B�=���ի' �E���Ǐ��^��ӧ�o���ȑ#գG!�%$$�k���;��c_�r�ᇙ�         `:tH���*��}�k��V}���w �l޼Ys��q�5 �E��I�&�	���o�Y�:uB�]�E�\[�l����u���         4�N�Ҹq�t��1���ׯ�1cƐ�R))).+SYY) ���mڴQ�.]��~��Gi͚5�7���[nQVV�Z����ݻ p�����ر�ڵk'          �L�2Eyyy·EGG��nc�/�YV�B�EEE8Μ9��^{M��\�' � �Ա��BM�6M��=��z�.\��ÕZ@೫'L���{Lqqq         ��U�\� ������Nedd��2܁�SVV�r���oU�^=�{܁:d��<yR��]�e��:���;��������'         ��B��ގoKHH��w߭&M���L��o߮��_�F���G��C�oǎ��<���C�1 x�\�R]�t�~�         �b�������˅o$''k�رJIIB�
 �͛7O;vTVV� �-�@�]����fW��=�p{���5�WTT@���.�LIII         �aΜ9.g�onMiii�Μ9�	&��SÆ��p���'�:;a����7�t�:w�,�>��NMMUaa� ���R����z��!         �.����\|�p{��|%%%z�7��_��P��u`�ԩ*..�~ȏ1B]�vM�����/�ԇ~�A�	         �+���?~�*++��Y÷��iMqqq���WYY� ��7jٲe2d� �mذA�V��v�uשgϞBx��1|f̘�nڰ         ��0e�	_������'JLLB�e*���r:tP������>t��	M�<Y�����էO!�؉r ���1슭�z�+�         �sk׮�@����$���?&�,����/ ��ԩS����#�<���H�-�M�6M��^�zi�СBx��N�6m�ʕ+տ         �bي�'
_KHH��w߭��d!�Q�]�vi�ܹ9r� �w�Grss9Y��u��Q7�p��,�n�gΜ��2}�tu��I)))         ��������L����5v�X����@p��{�.]ԦM������7� ��Z�j�[n�E����WLL��6���D �ˉ'4e����         �m�-��͛)66�5�7n�X܁�r��iw0��STT� �w�f͚��
w��{�m��~}����	w 8�_�^�֭S�=         xˁ��{�	Rdd�+lڴ�^���]����B ����z���5z�h�R������kٲe
wqqq�뮻��Y�����; 8Y�{VV���         \�3g���7�ԩS���ի�1cƨ]�vB������T
@�X�p��w���n�G�^d׏L�8ѽ�3;U|뭷*--M�Wj���ѣ�=�n�          .��ŋ�m�6A�����l!|YƆ�;\��[o��?����� �"�x�M�v�ڥp�Q�F�M�6�"���K��w��j۶�         ��***r�J����}�
�L�


4o�<��G? �"�xɡC�����+�0@ݺup.&c@��Ǔ&M�����:         ���=�7�xC'O�T��ҥ�,�L��ϟ��={�e˖�=�/�>}z�O�ڷo����J��$&&*&&F,R �mϞ=��?���C�
         ��+Vh˖-
w�[�֍7ި��܁�UYY���zK����U�^=�����jݺu
g��}��7�C��&���d�޽�f͚�^�z�aÆ         ����L���]jj�n��VկOt_#����<W8d�����Kd'��N��p�;�C���.��;���]���?��         ��>}��;�p֠A�u�]�������İ�� �����˕��, ���;p�/^����+\Y+��Q����&�b�w��:rРAjӦ�         ��ٲe�V�^�pV�^=�r�-��8�e*�����~�m�w�}p������Ds��U8�pcVV����J- t�9sFS�Lѣ�>�;         ߧ��B'Nt{L���k��@
��2yyy�֬Y�+��B]�t�KC�����u��	�+�t2D@upBK~~�V�\����         �>.ԁ�.��r���G��!S���S��?��?% �G���ݻw���Y			3f��>�.�N��͜>}Z B�;Ｃ�={*66V         ��>����+�eddhĈ.��;<�E������#��Ҍ3���,(�z�.��Ddd�RRRT\\, �����M�F�)         �\o���N�<�peي�n�M���pB�ܹsշo_W
�vxrj��>ӦM����V�Z	���pB˂4p�@w�         �غu�֮]�pe��G��@Ւ�����(�:uJ ��}Ϝ9S��w� �w��N�>�Y�f)\effj��j��7o��a���{Ocǎ         `,_1e��9sF�jذaj۶��ꈈ�Pjj�8  �o͚5.g���- 5G���e˖���@�A�3f�;a�Wj�i�ʕ�ꪫ���!         ��{��U��С����/�&,SA�o���{�1�v@-pj��ɓ�;w��5j�\
�@h��w�yG>��         ގ?�ٳg+\���h���.k��
 ��۷O}��$ 5C���E����D�w���ر��K�d]_|�6o���        �0g健��
G��k����X5���& ���w�u�;~. 5C��&�xY�=����ꫯ�qqq���WYY� ���3g�G��         Li�ҥ
WC�UFF��ڠ4=ǎӂ4j�(�>�@5͛7O���
7��������&d܁Д����?�\ݺu         "UTT(eff���w��Y�w��_W� 	�@���D�S9��֎�t���m����{g���1{k���tvg����*�(g-�H�� B!�����QAr�|>���gƙ�`5\��}]������~7��J=E&���@q����?�|6hx8wxW�^�w�y'�(��>��Ciƌq��� ��W^�e˖��     P2ǎ�ݻwGM�0!~��_e���J(�ڵkǝ;w�w��]��?�c G���C�&S6�gώ���C͕ZPlgϞ���?֬Y      ��o���N����~����RS!p��ٹsg���K1gΜ ������˗c���Q6�Dq�|UWW���� ���W_�U�V�P     P���q���(����X�hQ�PH�{�(�t ����}�˿�K �L�����_����(��>����w(�.Į]�b���     @��h/Mo/�����я~0T��ڻwo=z4�~�� ����ƕ+WJ9�=��)p��2eʔ����;w�P\���Z6ŽR�      ŕ�:u*�&}����,�������Pl���J���k _O�_����6_55^>��,�8��O(�s��ef��     �b���W_}5�h͚51����$p�b;|�ptvv�ҥK�j
V�
iz��mۢl֮]O>�d�pK2�;����x��gMq     (��۷���ts��/�0�cܸqq��� ��w��],Y�DK_C�_�7�(������x�F��Pi��|+W�      �%Mo�ӟ�e��ğ���Y�C-�|555eߵ�t���طo_,[�,���|��g������8Ə0�P�И�     �xv��.\��Y�bE<����%5w(�W_}5���Lq�� p�ظqc���D�̟??/^0R�P'N��ĢE�     �b(�������������&�Ŗ��wvvf�;�ew�O
�7m�eR[[?��OFRڌ�����_�pS�     P;w����G����?������dh �����X�t�)�� w���͛��>�2����S�NI�`Ŕ)S�ʕ+����>�;wn      �oiz�믿e�`��X�xq�p�C9��b���Y�|���{�nlذ!ʤ��1�{ѐ��ܡ<�|������       ����?ǅ�L��4�FB�)�D���� �����@���X�bۗ^z)ۄ�h�1cF9r$�rؽ{wtuu�6      �si�Q�|��ߏ�S�����L�<9�^�@�>|8�=O?�t ��� o��V���ٳcٲe�%�8�#]U��;�į~��       �����O��2I�m�;�	Iip����7ވ���sw��)�'ND�����mv��S��|�}����O~�Ǐ      �'Exe��ߪ��Y1�RSq�ȑ �o�޽q���hii	�+/�6n�e�dɒ�;wn�h�C�tww�����?�a      �/ip�C��L/^���#-� �C�������#p��_��gϞ=Q�����/��I�&E}}}ܺu+��x뭷�^p�     @���O�2I}�K/�0�ry����?�yL�:5 �;dRhw���(��k�:�ɘ�6d�O��<.\�}�Q���      �p�ҥ����L�{�9}�F���ŷ�~;~��_ p����m۶EY�i��?�|�X!p�rz�w�      9�q����닲H7��{�-QWW===���͛�'?�I�g�N�N��ڵ+�_�e��/d�;�NC9uvvFWW��      ����.�����_2������_(��7o���۳��N�N�	�e1mڴX�jU�X"n�r���-[��/~�      `lۺukܺu+ʢ��9�/_0ښ���P2�Ɣ��Q�T�L�N��9s&�=e���?�����;�W
�_~�娩�$     ���2L^z饨��
m�
(�.Dggg�������R{��w�,��������f�ԩY����@�\�~=����v     �1l߾}q���(��s��3�<0ܡ��z�-�;�'p��zzzb�ΝQiz��ŌE��2E�/^�|Ҵ�;     �صiӦ(�4��
�;������I����e%p��v�����Q)6���,m��PN����Ϙ1#      [._��Eve�hѢ�3gN�X1mڴlp`___ ����[�l�_��e%p���m�eaz;c]
[?��� �'mʶo�?���     ��%��[���R��/�0������ɓ�ʕ+��֭[�?�i�������R���#G�DL�2��vƼ��� �+:{���     Cz{{K5<pɒ%1k֬��f���w(�7n�|k֬	(#�;��N7���e���WWW�ei3�W�0�����x��      `lHQݵkע����W�X���ÇP>�������S:)l߱cG�A��h���c]ڌ��r���t�L�     0v���,���b�̙c���P^�p˹s�b���e#p�t8�/_�20����������Ҝ��lϞ=q��͘0aB      0����J31���*~���Uw(�m۶ů~�����S:;w�2H��;::�"m��P^w���"��{.      ]��ݲ���n3�555P^;v�_���R:wJe �+�u��yS#W�ǎ���{�=�;     �(Ka{������n�X6iҤ����[�nP>i`�}�b���e"p�T���[��޸q�bŊy�D<p����z�jL�2%      �;�˗/G̟??ZZZƺ4��̙3�Ӷm���RI�aˠ��#Ə�'w MٵkW���     ��غuk����?����Cy���i�{ccc@Y�)��7ofWu]�R�5k���H��}�;     �(���={�D<��1w�܀<�T@�����)(�;���Dooo]�>ˢ�<jhh�������	���?/^�3f      #k���q�Ν(��}�{y���@����{wJE�Ni�ڵ+�`ݺuy�nH��g�Pn����G     ��J�\L�<9�y晀�0�8q�D�?>fΜPwJ�֭[q���(�����Uڐ	��;     �Ȼ~�z)ڊd͚5QUU�ӦM����{�n �������/�PwJa�޽���E���|'��y��1��<y2.]��=     �������E����Ɗ+�$��S�LɾG�K�N��)�4	����룽�= ��@���{��_|1      )p/�e˖ń	�&5w(�O>�$N�:O>�d@�	�)�۷o������V�\�ƍ�3�;0 N�     �������2X�fM@�������۟��g�;� p����ۗE�E�����S�N�555EUUU)����ѣG�ڵk���      �4|(ݲ[tO=�T̚5+ �RS�k׮��/Ptw
��?�2x��c۶m����W��!#����c�ԩ���P?����w�      �>� ���v�,MpH���>}:�̙Pdw
-�q���Q===�	�����ĳ�>���Q[[�iC&p�;     ��z�j?~<�.��p�����+w�N�N�;v,�_�et����Y�~},]�4֮]���c]ڐ<x0 ���w��qP     `���i�`ѭ^�:�U�j	�s��� �-����Pdw
-M~-����/LuO�{[[�Mc����t3ɡC���Z      �4��*�J,^�8 �RSq�ԩ �����q�ܹ�={v@Q	�)��{��K�_y�l�{GGG<��1u�Ԁ�D���	�     �Ǎ7�ȑ#QtiB���ۿ��V���5 ����t���"�SX�/_����/����-[b�֭1o޼l�N*WUU�6�;0X
�����>      z��틾��(�������̞3f���˳^���> /��� I=ŏ�〢�SX����^:�|�ر�ihh�6o�W��ɓ'�����ĉ��>�����p�B477      Ck�޽QF/^�6��͛���-k%f͚0�8~�x\�v-�H�Na}����û~�z6�}۶m��SOźu�b��Q�TFZڐ	܁�=]�     0��޽[�����'v�ڕ=---�D�����������4�6����s����BJ/�]�zl`���i�b�ʕ�bŊl�6���!;y�d $����     ��9|�pܼy3���ٳٳ~��X�ti6pƌc�ԩS���:;���G	�),�;�t�ԩl"9�����ٕ\�6m��f'��͛g�;�Ήc`���h�5      ��{�_��ݝMt߽{w�H�VbѢE��bL����V^�x1 ������QS#�x�TSH酛���;;;�'������>`8܁�҇��V����      `h�۷/�j���q�ر�ihh��˗��իc����)5w I=ő#G��XP4w
����������T��k�ƓO>0������5�;     �иt�R�?>x8ׯ_�-[��֭[����֭�D�R	iMMM0��?�SHw
'M?z�h0�Ouoii�&�/[�,ƍ�L����q�Ν H</��r      ���p!���ӦM��+Wfτ	F����`�=������F�N�?~\;�Ξ=�=o��f���Ś5kb�̙�V:�N��'�����/      <�4��s���ذaClڴ).\�t#1#A�v���즑����"�S8�FGOOO�ڵ+{�������V҆L�Hq�ɓ'c���     �������s�����ٙ=3f̈�˗g�D}}}�p�������ի�D�N��ǆ����ׯ��K�ƺu벍<,2�~��     <�S�Nō7��w���l���͛���-�g͚0�Ə�&M����t3�����S(}}}q�ر`�����&��޽;�͛��R^�hQTWW|�;p?��      _��^===Y+�������hoo���ڀ����$p�j���E#p�PN�<�Ռ=�*�t� =�iGGG�Z�*�L�� w�~G���w�:$     �ҭ����g�f����c�ҥ�nݺ�1cF��HME� �+W�DWW�ފB�S()|c�K'H�l�[�n��T�ŋGUUU��tڸR�d�# �4��̙31w��      �����i+FIؘ&��޽���ĢE�w�[��Kؼ6P$w
%M'?Ouoll̮�Z�fM�א�f�<yr\�z5 ���;     ��s�ԩ,�f�n%b���z����qxX"V�~���{.�(���=��]��Mu߾}{vB9�TN'��o�+m���`Ǐ����     ��K�];�_���[�n��u��ł�|���� �{<E#p�0>��Ӹr�J�ow�ލ����I��+V�ʕ+c	A����ȑ#0 �      |;i�+c���ӦM�:��KL�81�A�N�555��� IWWW�O��(�;�az{�\�t)6l��6m��fS�[[[��p�p��/f�,�u�      <�Q06�]�|Y+�7JS��a�.��t�m͚5E p�0Lt-�t�t`�{
�;::�\}}}Plw�~�������      <�s���͛7�|�J�M�υ���ѣw
C�Na�8q"(�t���I�K�ƺu�b���A1	܁I��w     �Gcp`~��7o����X�zu̚5+(7Mp?�����BH�\O�>�G:���fOKKKvJyٲe1nܸ�8&M���>�u�V �     ��Do�����v�ʞ�V"����ʧ��) ;s�Lܾ}[CG!�)�K�.�F��Ξ=�=�ׯϦ��kVfΜC:q,f;u�T      �h�;���ĺu�bƌAy�����ݻYS1�����SB7���n'�H����իq�ڵhll      �Y�>�ܹsA���w�y��e�ĢE����:(��ST*������@���"�S�W�7pRyÆ�|��X�vmL�:5�Wj���Z�dI      ��N�<}}}Aq��9E��ihh�Z�U�VŔ)S�b����I�&����`�����@�N!���W�u�V�ر#v���rN�Bx�t�M�     �pR�Ny��y˖-�u�ֿ��/�����X�w�;0؉'�@�N!���7qR9��f�~��     �����ӦM��+WƊ+b�ĉA1��´f`�˗/Ǎ7� ����g�}�~�i��rR9_�N�555��� ��      �� R�aÆشiS,\�0k%Z[[�|kjj
���9s&-Z�gwr��ٳ����ʍ���I�իW;�<Ƥ�)r�x�b �p�B���9�     �zzz��V I��:;;�'M�����b���� �C���:uJ�N�	�ɽs��<�k׮e��7oޜ����[��^�T�ї6dw`���[� v֬Y     �WK��� 8�_WWW6�=�mmm�P@߿��x7�Pwr�w��ݻw�zR9]�bŊl���	��cC<HZ��     ����&i���]�����%
��������6y���ӝ;w`��~�@�N���p�t�RvR9Mv_�pa��kmmF��xk      �o&r�Q�!S�Y�~},]�4֭[3f�ƦJ��p��O`���糃/*�gwrO��p�����T��i[�jU6�}ܸq���b      ��R�����;��{��7o^6pѢEQ]]�-�������e�s��	�+�;�v�֭���OF�ŋ��c���[����W��Y�f�+m�ҩ����  p     �z�;V�+�#�;v,{b����`�)S�c������nw�L�N�]�p!`4���d'����Ғ�Tnoow��0����6�׮]���Q�@-�     �ˮ\����p���زeKlݺ��S�/^UUU��ijj
��H�	�ɵ��hK��ҳaÆ����6pN��t]N�s��<�A�a��!Zccc      �e�6����ӦM��+WƊ+b�ĉ��Ө ��"���	�%������cǎ��SOeWr-Z�(�����w�������ȑ#�f8� _%��      &pg�]�|9�iӦX�pa6���59i�{��:< `@�	��5��҆�����3iҤ�r��M�2%x����СC�k׮8z�hܽ{7 F
��ϟ      |�魌�������̞4Q���#k%����5nܸl(ا�~ ����Ν;Q[[�GwrM��Xw�ƍؼyslٲ%0�T�DUUUY���Ķm۲S� ��Z      ૝?>`���2MuO�D[[[�^�:f͚�t�@���ח5---y$p'�Dm�E�P~����<yr�\�2{�����7n�+W���e-      ���m�0Zzzz����3gΜl(�ҥK��F�6�nݺ�Mq�_Z��+�r+]m��!y�~n�~��x��wc�ٕ\���Q�T�Ҥ��^{-�= ��ҥK     ��������c��ӧ��7ވ���,v�6mZ��]�G��cǎe�N�S�WqЍ<��[W�^ͦbC^ݽ{7��ߟ=iӖ&��X�"&N�E��fq��۷`(�     ���M��
ƚ�7oƶm�b����0����UUU�WK��޽{㣏>�S�N��<������[i
4E�yްaClڴ)�,Y�Mu�;wnE�q��C�ٳ' �R�F�UWW      �3���,�����466fCӓ���ݸq#;�{������G!p'��䖉�Q
�Ӊ��477g'����c���W�������Z,����חE�/     �"Qyq�ڵl �ﾛMsO�D��^�T��zzzb˖-�s��lz;���y&p'�Lp������_�7�|3�����i�'ׯ_����������pIk�;     �	�ɛ4���?Ξ��_��bŊ�8qb�ɡC���^�}<�4D��ݻQ]]�7wr�w�"Mu���̞����r[[[�7.Ʋ������?����:     �e�g��wÆ�d��|Tw�܉�7Ǝ;`(��C���>}z@��ɭ�W���ٳg����}6ս��=�ݛ��c��y�f�����^k      �L�N
8s�̬�H�D]]]ɥK��׿�utuu�P��Wwr�ڵke�����^�����r����֎�?Z����o~�p�B ��tc      _dHEs���x�ײ��˖-�b�Y�fEޝ8q"����;nݺ Ć7�J�Nn	��4�==�ׯ��K��ڵkGu���o�G�	��bM      �E)�M�Ӡ�zzz���s�����������?��?q�Ν w�J�Nn��
_�>�صkW�<��Y�hѢ�����C���͛`$Y      |�����P��7FGGG�755E<x0���޽ �Ś����K)�}�v v�ԩ�ihh�+Vd�ɓ'���駟�+�����0�Lp     �"�Z)��7oƶm۲g��>�3g�������ہa'p'���I��pҟ�w�}7��>o޼,t_�xqTUU����?�1��`�Y      |QPe50���1V�\�=�Ǌ����Wܹs' ��իW�H�N.	��Ѥ��ǎ˞4�}���z��!��~�ȑ8p�@ ���.H�s�J%      p.$����M��w����+Ml��o~c� 0b�	�+�;�t�ƍ ���nٲ%��k��ٵ\i#�m�����lz;�hIuwwG}}}      `p 6x(�iӲ��+V���'��?��������0R$����͛7x<}}}q����ijj�U�Ve��'L��H��֭[�ҥK0���@�     p�i��`�/_�6d��.\�Mu�����СC�s�� Iih`j*F�P<�;��Z)P�7b�ƍ�������۷�h�6      ����^�����3{fΜ�loo����a��������o�)� #-Mq��7wr�w�7pӧO����,v������~tww�h�6      �\
ـ�s���x�ײ��mmm�z��5k֐�o����4�Q����7�;�dJ+�����^˵t��X�n]̞=���{���������A      ��ãK���ڵ+{ZZZ���i�{mm�c��.\�~M��b]@	��%��4���?̞�ܲe�b߾}���k     �����ٳg�g����P��k�Fss���^�������b]@	��%�at����x�k     �{��t#7��������w����X�jU,\�0���������ĉ0���:�\�}�v �'m� �k     �{Dl0������ѣ�3iҤ����b�)S�|�߷u�� m��GwrI� v�Ν      @���ƍ�e˖,^�7o^<�쳱x��/Mu?y�d�9s& F�g�}�7wrI� fm      p��FF��~�ر�6mZ�\�2V�X'N���m۶�X`�;y$p'�Dl �`�      ���`�]�|96l��6m�%K�Ă�СC08�F	�ɥ;w� � k     �{�������w���+��#�;�dJ+ 0��     �=�7 �6 ���R:� 0�w     �{Dl �`����\��� ��      ��� ����#�;�$b �6      ��ͷ �`w�H�N.�� ���      �� �Y�GwrI� fm      p�� ���7����R����\� �Y      �s���  ����UTWW���\J/�  �      ��� �������K��; 0�5Z      ����Y�7wrI� VUU      � �/�{�n@��ɥ�ِ �      ��) ��(L���% 0��     �=w �~&��7wrI� fm      p�	� ���#o�䒈 ��      ��J�  ��*��;�T]]  �      �� ��> o��RM�] �s���     �� �2��F%L.�7.  X      �S�T `0�;y#p'�Dl �`�      �TWW �`����\� �Y      �cB+ p?7��7wrI� V[[      ��
 |Q�ۭ��;�$p �6      ��`  `������;�TWW  �      �1 �ڀ<��K&L ��      ��� &p'��䒈 ��      � 0��y$p'���� `��     � 0��y$p'�� �`w     �{Dl �`���y#p'�&N�  ~     �g��� 0@SA	��%/� �`&�     ��{ `0k�H�N.544 @�����X�     $"6 `0��#%����  �u     ��� �`����\�4iRT*���� ���      �3� L�N	�ɥ���,r�~�z  ����      �SWW�u}}} ��y$p'�R�&p Lp     �\�R�&�޸q#  Lp'���V��Ξ= @���     �E���; �H	��-/� @bM      �E)p?w�\  H	�ɭ�S� ��i�     �� �. ��䖘 H�	      �H� $UUU1a����[&� �5     �544 @:�V�T�F�Nn��
 ���9i     p��ġ7�J�Nn��
 8�     �e�'O  k�J�NnM�81jkk�Ν; ���     �� ]y%p'�*�JL�>=Ν; @9��       _$f ���+�;�6c��; �XZ      �E&L�������	 ��z#���Zsss  �e-      �`ib�'�| @y	��+�;�fj+ ���      ��	� �;y%p'�Dm P^�J�Z      �+� ��RW1eʔ�<��k��� �Sڄ���      _6}��  �+u552a��O.���Ԕ� ��� P.��     |5C�ܬ�3�;�VUU���={6 �riii	      ̰  (7�;y&p'�R�&p��={v      �`3g� ��v#��䞸 ��w     ��6~��hhh��ׯ P>w�L�N�	����      �^
�� PNw�L�N��
 �3iҤl�      _m֬Yq�ر  ʥR�Dsss@^	�ɽ�"\SS��� ��n      �,� @�455E]]]@^	�ɽ���lCv�̙  �aΜ9     �כ={v  �c@�	�)�'�|R� %��O      _ϭ� PN� ���B0� �%n     ��555E]]]��� P&��ww
A� �QSS�f�
      �^�RɾW9y�d  �!p'��B���6e��� [�F+E�      |��	��<RK)p'�AB�Nkƌq�  �-l     ���Vv�� @9477gM%���;w�� J��'�      ��V �\��Ƽy����� ��Z[[     ����J���� ���"�Sb7 (�q���O<      <����GSSStuu P|w�@�Na�嚚���� ���ΝUUU     ��KS�� Pw�@�Na��=mȎ; @1��     �ѥ�b��� ��ɓ���1 ��ʼy�� P`�     �G�n� �逸�
(�;�"z�b�^     ���w,�J%��� (.]E!p�P�y�  ����9�L�      <�����5kV�;w. ��jmm(�;�2y��,~�p�B  Ų`��      ��I]� P\UUU��SO����I�� ��M-      �^
ܷm� @1���D]]]@�)��oݺ5 �b1�     ��kmm ����S$w
�tW (��S�FSSS      ����Ǐ����  �'��E!p�pR�6mڴ�|�r  ��      �㩪����~::;; (mE"p��-Z۶m �/^      <�����N�ӧO(
�;��d��; H:�     ��1� ��{<E#p��Ҕ�J���� �[KKKv�     ��3w��7n\ܾ}; ��H��@��)�I�&�O<�O�  ���,      <����hmm� P&�S4w
+Mq�@���t      �F��*p��hll����"�SXi��o� @~�)"��     :i�Ы�� @1���J�P$w
+�p�Ǐ����  �)�����      Cc޼yQ__�n�
  ��0`(�;��&���I|�A  ��lٲ      `�TUU�cϞ= �[�ܞ:I(�;���8�; ��     `�N� �����'O(�;���ޞ�P���  _fϞ���     ��Z�dI  �gz;E%p��b�ܹq�ĉ  ���v     �ᑆ555ťK� �/��(*�;���8�; ��     `���b6m� @>�7.�y晀"�Sx�ꫯ �'N����      ã��]� 9�x�⨭�("�;���O�̙3���� �C:�VUU      �����㣻�; ��I��@Q	�)�ɽ�� ��ʕ+     ��SSS�-�={� �/�JE�N�	�)��	� &L��}�
     ��Ja�� �gΜ91eʔ���S
s�΍����t�R  c[{{{61     ���4���? ��0���SQ
i3���7n `lK7�      0�&O���͋cǎ �+V�(2�;����
�`�?~|,Y�$      i��� �c���1gΜ�"�S����{WWW  cS� ���6      �����������;���?��a���c AD���QA0"���hS��[�&�$�MbV�ny$�dc��^+I���w<QO0FQ��>_�嚣g���z����-���3���TUU ��Ұ_h��䍂��2dH�q� 䦡C�      ��u�����_= �ܗ6�AC'p'�TTT� G�h�">�O�  n�IDAT��      �v�PN� ����,�t���	��+:t�N�:Ŋ+ �-餕���      �v80n��  r[ڔVPP��	��;C��@J�;      ��}��@=p衇��;y'�i��m� ��ڵ�8       �@nkݺ����!p'�EϞ=c��� ��Ç;B     �����o����  rOEE����!p'/��N� �!]|6,      �;i`��K�.  �2$ _��K�f͚���� �[�{��~`
     @�JS�� �{:u�;v�w�RqqqvQv�=� P���*      Խ�����Ɩ-[ ����o���	��n���f'�      P���n���O>�d  ���� ***����եK��ܹs,_�< ��1lذ(*�      W���w ��{������|�&"�~��q�u� P7F�      �C9$��g�x�� �{i���;y-�q�7Ć �]tPt��1      ����YO�hѢ  �Viii���? ���k%%%1lذ��{ �]GqD      �{�)�w �{C�����|#p'�5J� ��E�1`��       ��������J  ug����H�N��СCx���lٲ  jǈ#���GQ     �\UYY)p�:Թs������בG)p�ZRXX��@     ��5t�����~�ׯ ���5* _	��4(��w�x�w �Y�}�M�6     @�*..�aÆ�]w� @�jڴi2$ _	�!>�$�v;���� �f�3&      �}GqD�}��QUU @�I��JJJ���Oeee�v�m�q��  jF�.]�[�n     @�k߾}���#�,Y @�9������O�f͢��"���  j�رc     ��#Mq�@�I��:v�����	�G������Z P���bРA     @��~��~ϳf͚  j^�!�	��:t��rH<��� T���:*5j      ����1jԨ��� �Y�[���;�;��c�9F� լY�f1r��      ��9������o��7 Ps�<��ls�;�;��8 z��K�. �z��&M�      �OfTQQ��{o  5���$F���vh���w �&���ٱ�      �_GuT�w�}QUU @�>|x�������7:w�˗/ `�92Z�l      �_���ѻw�x�� �^1z�� >"p�Hocǎ�+��2 �=רQ�l�      �߸q�� P�ڵ�#w�C���n�-�z�  �̰aâM�6     @�׳g��֭[���� T�����ww����q�1��UW] ��K�G}t      �p�;6.��  �G�^��K�.�����СC���o7� �@����,     ��e���ѡC�x��7 �{���g	���ɳ&L����: �]gz;     @�TPP�Mq��/~ ���ܹs���3�O��NTTT�w�a�; �4����<      hxRKq�-�Ě5k �s�sL�y�4�;�D�@��D���  v�Q�F�{'      SQQQv����  �Lǎc���|��vA�y��?�!V�X �9rd�m�6      h��������w �C�&M2�>��vAz�<yr\r�% |����0aB      а�)��Ǐ����7 �:��_@�����ѽ{�x饗 رѣGGYYY      ��UVVƝw�i�; �c�=��v�w�S�N���� |VӦM�)      �S�`�u��1����n�ѣG���;/^ ���7.JKK     ��������U�V �s�'O6�vB����㏏^x!�m� �GZ�jGuT      �_���'�5�\ ��ҥK0 �/&p��ԩS�8��� �#S�N�ƍ      �gذa�hѢx��7 �|��0�vN�{�㎋�<6l� ��:w�     @~*,,�ɓ'�e�] �����#z����	�a�l�2Ǝ��rK @��>}���      yn���q��+�� �gM�6-�]#p�=4~������c͚5 �*���gϞ     @~K��L�?�� ���Wt��-�]#p�=T\\�w\\u�U ������b      >֫W��۷o<�� |�Q�F1u�� v���BEEE6�}�ҥ �f�رѮ]�      ��N8�X�xql۶- ��Q�FEyyy �N�{!�5s�̸袋\��W���b	      �Ծ}�9rd�{� ��Y�f1q�� v���R�Ν]��w�O�%%%      �h����裏Ƈ~ ��R�^ZZ���C58���'��>�  ��;��c���      ;ҢE�?~|�t�M ��m۶1jԨ v���A�a5eʔ��� �F���'�      �g�ر����ʕ+ ��	'�EE2]��s��TVV�C=/��R @Cu�QG�~��      �ER�7}����K �M�^������;T�4�v֬Y�����u�� ���u��1q��      �]�¾�}�Ƴ�> �/�&��N:)�='p�j�&ڎ3&-Z �Мx�QRR      ��fΜ/��Blٲ%  �����<�='p�j6iҤx�'bժU š����      ��ڵ�B�;�3 ��kٲes�1��;T�ƍgǋ\|�� AӦMcƌ      {b�ĉ��#�Ě5k ��W4i�$��#p�зoߨ����~8 ���>}z��>      {���$fϞmX  Z�>}bȐ!�=�;Ԑ�3g���?k׮ ��z��#F�      �iX`���㩧�
 hh���㤓N
�zܡ����f��/�� ��h�$����      ���¿_|16l� АL�81ڶm@��CJ;��?�x @}3u�T_      T�����4iR\�� EǎcܸqT�;԰�O>9�,Y��~ @}ѭ[�5jT      @u=zt<��#��k� �w1{��hԨQ �G�5�y��Y�~�e� �%%%1w���"      �Saaa�r�)���~7�l� P���[ݻw�z	ܡ4(F�<�@ @�;��]�v      5�S�Nq��Gǭ�� P_�n�:�L�@��C-�9sf,[�,�z� �\էO�9rd      @M�8qb<������ �71gΜ())	��	ܡ��7�y�������غuk @�i޼y�z��E      Ԥ���8�S������z���2z��@��C-�ҥK{�q��7 �Y�fE˖-      jC�Νcܸqq�w �eee1mڴ j��j��G�/��K� �#FĠA�      jӤI���矏W_}5  ���ٳ�iӦ��;Բt�ּy��_��_b��� u�]�v1cƌ      ��֨Q�8��S㢋.�M�6 �ѣGG߾}�Yw�鈒�����/ �KEEE1��hҤI      @]�СC����_�:  W����S�P��PG��� ԕ�ӧG�Ν      �ҨQ�b�����SO �����đ��� j����I'�˖-�իW ԶtdV�A!      �9s�ī����^ @.�4iRt��5��!p�:Դi�8����G?�Qlٲ% ����q�i�EAAA      @.hѢE6��?�iTUU �=z��G@��C�֭[�p�	��_�: �64j�(�`UZZ      �Kz��Gyd�u�] u�Y�f1w��(,,���!�5*^{�x�� jZ�Xս{�      �\t���ǒ%KbŊ u�K_�R�n�:��%p�q��'�o���� PS=��l�      䪢���7o^\t�E�y�� ����0 ��'p�Q\\g�yfvq�� T����3gN      @��رcL�:5~��� Զ�>4}�� ��rH:���N��/�8��� �K�&Mb���-      ��G��%K�ēO> P[JJJb�����Z�n�!����'&O�7�|s @u(((�SN9%�]      �E�=�ܹs�{��^��� ���O�:Pw&L����z��/	 �['N���      �7���:+.��ذaC @M:��#cذa�-�;䠴��SO����ov �W����{l      @}U^^�Mr���UUU 5�k׮1}�� ��rTځ�`����w�k2 {$����N�6N     @}6`��;vl,Z�( ��5k�,�8�(*��B.�9�}���$��.��d vKiii�}��Ѵi�      ��`�ԩ�bŊX�xq @uI��͛mڴ	 7�!�80�L�7�tS ��hԨQ̟??��      Eaaa�~�������z�� ��0mڴ�۷o �C����	����/ `gN<���ٳg      @C�N2NÞ~��Ė-[ ��СCcܸq��;�'�tR�\�2^|�� ��3~��8���      ��]�fC����� �=թS��3gN �G��D�F���3ό�}�{Y� �h���1u��      �����2^y�x�� vW�-b�Ѹq� r���t��W������k׮ �.M��;wn      �Y�f��o�K�,	 �Ui��g��[� 7	ܡ�iӦM�s�9��(6n� жm�콡��$       _�@q����}/V�\ �3ip�)��|p �K��P�.]�d�\rIl۶- �_�Ȭ/���-      ����8������~�_�> ��L�0!�@n�C=u�!�dGm�� �S�ƍc�Ѯ]�      �|վ}�8묳�'?�Ilٲ% `G�'O �	ܡ9rd�Y�&n���  �řg�ݺu      �wtP̜93��� �t��i���>�;�s�&M�M�6ŢE���PXX��zj���7      ��~����;��w� �]۶mc�Q\\@� p�`ڴi�aÆ���{��-�$�5kV2$      �O�2eJ���{��� 4o�<�=��hٲe ����;�|�ɱq��x����k���1r��       >+5�g��"��{. �_ib��g�����/wh �ک��[�n��{, hx�N�GuT       ��Q�F1����˗/ �Oaaa�~��ѭ[� ��;4 �My�ܹ�$�g�y& h8�=��8��      ع&M�Ĺ瞛E�+W� ����<@�$p����(�<����OK�,	 �ѣGǤI�      �u��O|��_����z��  ?��1bĈ �/�;4@���q�9�d���e���k���1cƌ       v_YYY�w�y�$���{/ h؎;�;vl �������,r�����믿 �?��9s�dGg      {�]�vG��֭ ���:*&L�@�'p��iӦ��/9~��śo� �)n?�3���0      ��ӱc�8���A��ׯ �#�<2N8� �;4p-Z��o|���$^}��  �2$N;�4q;      T�Ν;ǹ�?��c�ƍ@�p�a��̙3h8��5k��u���K/� ���ʘ5kV      P��u�.����g�y�� �~4hP�r�):h`��}۶mU4hM�6��|�+q饗���? �Q�Fŉ'��      jPϞ=�3Έ�.�,�n� �O}��y��Eaaa ���}[ ^III�s�9q�WēO> ����Ǵi�      �y�����O?=k(�S �Oڬt�YgEQQQ O��]����=�B���+��� �V�֞��q��      P{_�җ�k���#|p,\�0���h���>�AI�{څ�&�?���@�Hq��3b���      ԾaÆEӦM���/�-[� ��o߾�`�q;4pY�m�6�!��)���]���O
 jWz�3gN><      ��ӿ�8묳��?�yl޼9 �M��z���ـW�a����yh���&M��m�� Ԏt�5o޼��C      ��_�������cÆ@n:th̝;7(4|Y�y�f��@�<yr���č7�UUt �IiSQ�MܧO�       r�A�~���?�u�� ������O>9�
�,pߴi�������m۶q�W:n���l�2�9��ҥK       ��k׮Y�����$��� �n��m�ԩ�v�3Y�q�F5+��V�Z�%�\�"���k�.�=���      �]�;w�����o��o��� u#��ӦM �l��.p2ݺu�/�0.������� ��ںp��hѢE       ��}��q�d���U��ړ����1v�� �S�oذaK ��6m��7��l���e��=7x���;wn      P�~�k_�Z��\�2 �y)n�5kVTVV����}�ƍ&��RZZ�~�����~8 �}�G��3fd_      @����ƅ^�^zi,]�4 �9EEE��C=4�������� ��?0�m�6n��� `פ��ٳg�a�      @����w�yq��Wǣ�> T�f͚��G��=p� ;��O�4)Z�n�^{mlݺ5 �|�[,��:(      ��!��7o^���P�R�v��F� ��w�}wc |��ÇGYYY\q��nݺ �:v��&N'_       ��!����կ~eH @5�o����=��l�}����Q�F�yz����ַ��K/�7�x# ��~���i��M�6      ��9rd�j�*.���ظ�\Q�=շo�8�3�I�&�IE��|��Ѽy� �"i*�7��͸���'��|��4�7.�N���      �e�~��/�5k� ����2N>��(,,��q�~�z�;�KJJJb����hѢ������* �Q�A<w��0`@       �e����/�0~���������KA��3��#����q�nݺ �UiJ���㳋�+���k�w:v�,����       �S�V��.�+��"�y� ��A���~zr�!�E>�׮] �+����|'.���x�� TTTĬY��-      ���~o�p�¸���㮻�
 >+<묳�C��3w`�����׾����\�ZQQQL�6-ƌ       ��̙3��_���y�� �#i��y�Y�f�+>���� �S)��~�v���ƍ�!�w�}c�����      ��:4�N|饗��ի �ĸq�b�ԩ�}�]e�;P�҅Z�.]�+���˗@C0p��8�S�$      v�s���o}+.���X�dI 䣒��8��ScРA���@�+//�/�0n�ᆸ���* ����l�1c      `W�h�"�?���馛bѢE�	 ��~��3ό���/ ��ǁ�{� ե��(fΜ�rH\u�U6� �N:6��3�p�      ���6mZt��-���X�~} 4t�/}�KѴi� �S�k֬	��ֻw��������+��_�\WPP�F���?>��      �7�غ���cŊ��M=�w\�?> �ƺu�����m۶�E�:�j�*;v���������iӦ �E-[��9s�D�~�      ������7��͸��⡇
���u��1���ڵk �w�y���֭[c�ڵY�
P��D����8���i�z �A�ŬY��y��      P�7ns���n�򗿌?�0 껁f�KKK�:|*p�����I�ȭ/�0n���l��# �R�&Mb����&      ��6x��l������/� �QqqqL�:5ƌ �i͚5��� 5�Q�F1iҤ�ݻw\s�5��[o@]H�Ci���       ��u��q��m�ݖ���� �/Ґ��O?=:u� ��3�W�^ ��{����|'n�����`�;Pk�6m�|�92


      ��f8��l@�ڵk ����#���ӧg�j�g�U�V@mJt�M�C��.֖/_ 5�o߾1{��(++      ���~������q�u��_�� �E-[��9s�D�~��&���۟�W�\ u�s��q�f�n�y睱u�� �N͛7��3g�СC       ��h�",X�?�x\{�~�� ��ʆ	���@MK=���EEE1eʔ6lX��W��^x! �V:���";+�P       W<8�v�W_}u,Y�$ �R�&M�ޢ��2 júu벍~�
��y�زeK�ԕ���8�����믿>>��� ��ڵ��O>9z��       �A�֭�_�j�u�]q�M7ŦM������7��^VV �����n?U�WUUŪU��}��P����4ɽw��q�7d�{z���5���:*&O�l�      P�nb̘1ѿ���//��B Ԇf͚Ŵi�Lm��ʕ+�ۢ}A�䊖-[�ܹscĈ���&�x� �"iZ�̙3�C�      P��i�&�;Ｘ����w��]lذ! jJ�~�b֬YѪU� ������ً@.9蠃����v�}��q�-�ć~ �Զmۘ:uj<8       �4�=MR�ӧO\w�u���@uJCH�0�C=4 �R�ؓ����_ f�o6,n���,v���
 �5n�8ƍG}t      @C���ƹ�O?�t��W��5k���Hh***bƌQZZ um{Ǿ�	� �,}�J;��_}������Y�w\���      @>�ׯ_���#���+��ضm[ ����/f͚ݻw�\�>Ӭ\�2����=MDN�@.�֭[|���v&�������~;������O��"      �KM�6�x8�u�]+V��]Ѹq�8qb�;65j �⭷ފ-[�d�?�oڴ)V�^mڴ	�� �L�ӧO�+��[o�����0�k�.��>h� ��      �����}��ߎ�~8������������O�֭[@�ICڷ+����׿
܁z%�&3fLTTT�����{ol޼9���e˖q�1�Deee       I����rH60ܶm[ lW^^�������ԯo��B���_�v� �7͛7�3fdG��v�m���h�z���$F����M�4	       v���4X;���o~/��R �-u���0a���@�[�|����v������,fϞ�}@K��Q\UUU��*��eʔ)ѢE�       `����q��O<����cժU�t�CEEE��Ѳe� �Ҁ���@���י;wn�3&;��駟�C+..����?~|�j�*       �})n<xp���/��l8��h�z��ӧO�N�:@}�~��X�f���a�z������y������.�7�x#n��l���r�����{��      ���!ci�؈#�^�{�m۶��t��!��~�!�@}�����,��'�)�i'@C��~������}ѢE���ݡ	�      j^t:s��8�����o�'�|R/D�֭cҤIQQQ���P����>7pOO�U
��Ν��R���;��G��[�P;�4iÇϾ��       �#Mx^�`A����D���~:��)m\7n\�=:;��>K��?�s�W^y% ��;f���ɓ��c<���q�� jF˖-�� cƌ�f͚       ��k׮q��gǲe�⦛n��K�P?���ĨQ��c��4/����,p����IGqM�81����{�>�z�o�>ƎÆ����       ��x�����=���,tO�݁ܔb�#�8"�>�hC����ߏU�V}��-��}��X�fM���@�HG�L�4)&L��=�X,Z�(�x� �L��ݳi�����        ����+[)t���G�"l��ޞ|��� �&M�N���J�q�u�]��%�m��K�?�zh�7.��o�       �~��?��q�m��08jGiii�=:,شi� h�v������@�K�q���[o�����ğ���X�~} �ֶmۨ���#Fd�!       P?���7[i(��w��<�LTUUP�Z�l�~xu�Q�v /��w >R^^3f̈iӦ�SO=��w_v4䳂���ٳg�80
      ��a�P�+V����x�Gb۶mT�4X��#������� ��s�k����ǿ0pOaӦMѸq� �#EEE��i-_�<���裏Ɔ�ž��Mj9rd�j�*       h�:u�s�΍I�&e������ظqc {�G�ٴ����g���믿�����-[�dS��dV >�s��1{��9sf<����T�^x��\4HisG��6lXv�i�       ��M�6q�I'�ԩS��?��O�z�� v��#��ݺu�|�dɒ>���{�t�R�;�N�c��Ou_�jU�S9-q4]�v��Çǐ!C�Y�f      @~kҤI�3&F��<�L�u�]�����Ś6m�vX�7.��� ߥN}Gv�^������H��^{�x衇����k���[��C=4F����       ���� ��뗭7�|3���l��ƍ��.]�DeeeTTTD�ƍ�����x饗v����Jl޼9�N��IN�:���_�b�'�|26l��kZ�j��N"�޽{��       �:t��3gƔ)S��G�{�'V�X���IC��#�8":w� |�o��֭���v���=E�tP �g
�W�^�J���X��<�z�����J:�o߾�n�t���      ��JQo�T�ֲe�����'�x�Tw�F�n�b���1t��())	 v,�<;ܓb
��G:c��\۶m��_~9��{�X�vm@Mkݺu���ߤv       jԁ��Y�f��O?��w_���QUUА���ƠA�bԨQѩS� `�}�����.�/Ύ��z�i��/�N8�X�|yvA��3��k��Pҿ�t��!��m����E�       Ԛ40aK뭷ފ?�������;�P_e-�a��ݦ>�]�y��X�t��~}���_=֭[��2�f��]�t�֤I�����B���#��:���ݻw���o߾��      �	���q�q�e+�{衇��G���? ץ��ݺu�6kTTTD�������/~a�K���m۲�aҋ2 ��m۶1z��l���?�����q�x�.>i����={F�^�⠃�F�       �� �O��/�Gy$�aÆ�\����]�Ɛ!C��C�}��' �;�>��~}��$E�w�����J�rZ�ڵk?��S��r�� �l�{��E�)h/))	       �o� �tByZi`j"R���O��N�HQ������L��۵k T��{���ˁ{*�Ӵ���@�jٲe��9�$�K�.�b��^zɄ�h{�޽{�8����͚5       hH��~��e��O�_|1�x�,xO}Ԕ��"8p`�Lj�i��Ά��r�f͚X�bE��[R�N��~�F:��W^ɂ����}ݺuA��.��1li7p
�S�޸q�       �|QTT}���V�׿�5�y�xꩧ��_6���VZZ={��xS�a� 5/]ߙ]ܓ��@����4i�M�N+It��߲�=�˗/�6-����6(��״R�~�DYYY        ױc�l�?>�}�ݬgK�\�����LAAA6l�w��YО�� �����sv+pOǼs�1@��>�w��![Ç�K���o����)zO���Z�z��5$�,o׮]v�ݩS���vGZ      ��iժUTVVfk۶mY���/���?K�.�-[�$i�`�=�A�)j�i ԝ͛7ǒ%Kv���
�_}��X�vm��@����[�5x���ߴiS����J�{���B��қ;���j۶m��v�Ƃ��?       P}���Ӊ�i����D�ϥ��˖-������6?t�AY�~��Gyyy ���sjwf��4�7�}�/ O�ƍ?��������J��ʕ+���;�|��{ｼ�,..�����w�}��6m�|����͛       P7�4i�M�N+I��K/��MvOa]
��k8R�ѽ{�����n ���{�]z�n��O<!p�Ci�{���J�(��)rO���5k�����V:�#���׭[~�a��ߗ&��h��㕎�J�z:�$�O;|SԞ�       �)x�ӧO���8��S��&����kٟ��?r[IIIt��)�x��f����xꩧv�y��/^�8�KKK �K�}m�w&]��}����Ziwt:~d�ƍ�u���9�o?i��?)MUOk��7m�4������4�>�O�����o_�b       h�R�бc�lUVVf�}��Y�|��W:�^�^wRϱ���G�Ν���o�>kB ����U�v鹻�����'��#F ���޽YU����c} �����$jlJM|%F�ֶ��M��δ��&M�S'�tҙ���bZQ�5���@�"��G��օ]XvY��.��۞�BMb"�}�{��3�s��=砻�}��ږ�       �PK>���[��\.�x�hjj����ؾ}{zL>Ş��,,L�����~�A��z�@�X�r����������         �����'N��Λ%�ޓ�}ǎ���;w�L��'[i�O�筍;6N?��ÓD�g�}v�v�i�V} J[]]�������ק�B;餓         �E����.H��
�Bttt��{[[[�޽��$�'�8p JQ��|�����$dOfܸq�ׇ���Ç �)�4��MaG��|>�V�W]uU         @����8w�&]]]��ٙ.�ݳgOz<�8�������><�\.�BUUU�=���5*��IB�d���'3lذ ���r�ʣz�1��˗�        �UWW�3~��#z}��P���חｽ��$��e��^��%�9�~��d���M�#G�L��$^O��#F��O��m���t�G������]c��rJ          �+�
h�: ����hii9�s�9pO��UWW�\sM           ��-[���9��=����          �f�B�+V�y��oڴ)v���ƍ           H�_�>:::����
ܓ�>��~���           $�.]zL�W��X�xq|������           ���߿?V�\yL�w����7n�.�            (o���ӹ��'�-�w           �,Yr���K�����ԧ>���          @yjll�m۶��������k�?���           �i����u~��E�	�          �TOOO����u�~ܷo�1a           ��$q{.�;�k�[��H���          �Oғ�~ܓ���o�ѣG           ��7ވ����N��i�~��W           �?��'�5pO���+q�UWEEEE           P�zzz����_���{SSS�[�.���           �m�������/����=1o�<�;          @����`��~�ހ�?���c۶mq��           �iŊ�k׮~�ހ�_|1n���           �4͟?�_�7`�����S�L��c�           ����>^��~���}}}��K/�'?��           ��̛7�߯9`�{b��O|"F�           �����X�zu�_w@�\.K�,�뮻.           (s�΍B������=��/Ƶ�^Æ           ��޽{���v@�=��{{{{�X�">��           �m�����; ���=��/�����FEEE           P����.��J���Ԕnq����          ����/FWW׀]P��̙3��.����           ��twwǂ������Ĳe�b���          @q�;wn��A����/�<����           �}���K/�4���Ҽ��-�.]��G          ����s�E.����*�9s���ɓmq          ({��W^yeP�5���ݻc���q�5�           ٖlo?p����kH֨?��q�W�	'�           dS��|ѢE�v�!	������          �lJ��<xp��7$�{��矏�|�#1r��            [v��?��O��C��ݻ7�ܧL�           dˏ~������{Y���7o^\q�q�g           ٰaÆ�����i�~��������o�=           z�|>�z�!����_�n]L�4)           Z�-����!����������          ����3g��3�777��ŋ㪫�
           ���ٳc߾}Cv�L�g�y&>��Fuuu           0�v��/����2�wuuų�>7�|s           0����+�����ߐ��=�`�����?g�uV           08֬Y��P�T�����G?�Q����m           0�����,�T��H��������K          ��5w��رcGdA����?^xa�=:           ���1gΜȊL�QSS����          ��W(������ȊL�ŋ��_]tQ           п�f{����%��������c���          @���쌚��Ț����֘={v�t�M          @�x��ǣ��;�&Ӂ{b�ܹq�e����           �U�VE]]]dQ��|>������O�Æ           �M.���{,�*�{���)�ϟ�_}           pl�~����般*��=1k֬��K�3�           �N}}},^�8��h��������aÆ           G���'}��(
�eE�'�瞋o�1           82�=�X���F�U���3gNL�4)&N�           �v+V�����(E��������_��c�ȑ          �[koo�3fD�(��=�k׮x�'��[o           ~]�PH��wwwG�(��=�t��x�{��Ї          �_6gΜ����bR��{�����'Ʃ��           �-[��g��bSԁ����ӕ�������          P�zzzb������Ŧ��ĦM���矏?��?          �r��ODKKK����gώ/�0&N�           ���W_������bU�{�:ڴiq�=�Ę1c          ���ر#f̘Ŭ$�Dggg<����/|!��J�?          �m�r�tixr,f%U�o޼9jjj�[n	          �rP(�?�Al߾=�]I�����y��'O          �R��s�E]]]����3f̈��>;�=��           (U�֭�Y�fE�(�����7���o�=�����          Pj����{��^���(%�'��~����������          �R�,��w����RR��{bժU1gΜ���          �T<���e˖(5%�'fϞ�x�;��/          �b�p��X�dI�����B|��ߍ��+�=��           (V6l���z*JU��\.=�P��?�c�;6           �MsssL�6-<��,�DGGG<���q��wǨQ�          �X�ٳ'�N����Q��&pO$�X��w�w�ygTVV          @�����q��ݻ�ԕU��X�vm̘1#����<           �,������c۶mQ�.pO,Y�$�<�̸�           ��|�����~�,�ď��3fL����^           d�/�/��r�����B<��q�i��ĉ           +V�\�.�.7e�'z{{�[��V�}��q�g          �Pۼys|���O�z���������/��t�;          �Pijj��z(]�]��>pO������ߟF�cƌ	          �����<�@twwG�����;wƽ�ޛF�'�|r           �C=sggg�3���z��������          �������tttD��������:uj|�󟏑#G          �@ٻwo��{׮]���-���������>��1bD           �����4n߾}{���`���1mڴ��;����&          ���r�4n߶m[���ۿ�������������          p�8���7���1�e��QWWӧO������aÆ          �����I�������	܏�����_�������Ç          ����S�FCCC���Gh�������w�#G�          �#�w��x��b۶m�o&p?
�� �w�}�w�wQ]]           o���3퐛����N�~������}�sq�'          �o��֖�ǭ�������[��׿�����?cƌ	          �_��Ғnnooo����m߾=����������i��           �$�q�����#8r��k׮��7��F�g�qF           lٲ%x�����
����8�޽;��~�w���          @�Z�vm<��Ñ�傣'p�����&��n�->��          P~�,Y�=�X����F��Ozzzbڴiq�-�ĵ�^          @y(
1gΜ�5kVp|��(�����عsg�|��QQQ          @�:x�`���G,[�,8~�0��hkk��n�-N8�           JOWWW|��ߎ�7�C�>@^{���7�w�qG�|��          ��]�v�ԩScǎA��������W�w�yg�?>          �������ַb�޽A����_��W�����.          �x�X�"y�������}tww�}��S�L�n�!          ��R(b�ܹ���8}����|>555�������cĈ          d_WWWL�>=֮],�� [�lY477�����~z           ٵm۶�6mZ�ڵ+x�!�lq�������[�K.	           {jkkcƌq���`p܇H.�K��q����M7�          �|>�<�L�������B���ҿ��q�m���ѣ          :��|'��'pπ5k�Ŀ������g�}v           �o�ƍ���Gggg04����_��W��o�+��2          �������矏Y�f��:����3f�ڵk�3��LTWW          0pv���<�H���CO��Auuu�y����g?_|q           �o�ʕ�ꮮ� ����=�P|���O~�QU�G          �!����O?�-
�E5�a�B!�ϟ�֭��n�-�9�           �]cccL�>=Z[[��������򗿜nr���k���"          �#���c޼y��$����l�����x��'c͚5���~6N9�           �^[[[<��#�q�� ��Ef�ڵ����q�M7ŕW^          �[+
�x��x��#���'p/B]]]1cƌx�������bܸq          �����x��G���>(�"�f͚����������xTVV          �����x��c�̙q�����܋܁���&~����g>�?~|          @9jhhH��777�I�^"6o�_�җ�뮋?��?��*?Z          �C�4z���1o޼���A�RA����^x�X�zu��}	          �l͚5���G[[[P��%(�H��~��q��W��ܫ��          JI{{{<��ӱ|��t�KT�P��_~9�-[���Ǣ�ʏ         �����,�9s�DOOOPZ�%���;jjjbɒ%q�-���_          P�V�Z?�����-(M�2���S�N�I�&ŧ>��?~|          @1غuk<��S�q�Ơ�	��̺u��K_�R\s�5����1jԨ          �,ڷo_<����K/E>�J����������c�ҥq�7��{eee          @$���'?�I�r��|��XWWW<���ӟ�4�L�_|q          �P)
�lٲ�5kV�ܹ3(?wb۶m1u�Ԙ0aB|�������          �%	�W�^�nlojj
ʗ������fL�81��O�4.���          ���nݺ�����[���5�7o�{�7���wŔ)S���~w          @J��g�y&��mڴ)����ǤI�⦛n���??          �x$˘�����>�W	�y[ɻc֯_�^zi���Q�s�9          Gc�ƍ1k֬ذaC�o"p�
�X�re:�z׻�n����}QQQ          �V�u�����s�ECCC���s�6mڔN����k��ɓ'����          ===�lٲ�7o^���)�;Ǭ��)f̘3gΌ���:>�я��ѣ         ��w��X�pa,X� ������������f�J�a��8���7n\          PZ[[��_�W^y%z{{����~���b������/�<����x�;�          ��B��ׯO��5k֤_�����������6��������率�O<��          ���ٳ'�.]�nkߵkW@�3��o�5551s����>W^ye\t�EQQQ          �C��-Z���Z����Aq���X�bE:g�yf����+���N:)          Ȧ��������F[[[�@�3�ZZZlu         Ȩ|>6lH����ե_�`�3d޼�}�رq�e��?���0a��         `
�hhhH��W_}5:;;����Lhoo����3nܸ���K��}�ĉ         @���Ew2g��݇c�SO=5.���;         @?ٲeK��֦a{GGG@��ɴ���ñ�Yg����Ɍ?>          x{ɦ����X�|y����d������ܜάY�����y�{bҤI����7F�          �BWWW�_�>֭[�W�����!p�(%��-Z�NeeeL�0!�����E]�w^TTT         @�H��oݺ�pԾaÆ����F�N�K��nڴ)���'��nwO���8jԨ          (5���KC�$h_�jU�ٳ'��	�)9����t��t�����|g\p���w�;��>bĈ          (6]]]�q�ƨ��O�۶mK7�C)�S�<��O&1lذx�;ޑ��'NL���N:)          ����-bӦMiԾ}�vA;%O�NY���͛7�s�駟�nvOb�d�9�t�;         �`��r�u��4hO���_���΀r����ܹ3��������������8�����Ϗ��ǧ����         �xuww��طlْN���� p�_��磹�9��K�~~̘1i�~�Yg>&��G�          �*	ٓ%�I��t����v�
�	��utt��nݺ��UTT���g���駟�N����N��#G         P�:;;�`=	ٓimm=|ܷo_ GG��!�(����t6l��k�5jT�;6N=���8nܸ�x�'�)��'�tR:Æ          ;8�����ݻ7=&�r������w���� �ϡ�����_VQ���QOOO�ر#�ߦ��:�ޓc��}��ч'��G��F���UUUq�	'�����Ǉ$߷1        �r�,������璖/���������/r�\�'����$�O���+ړ��4;��笇.���{�ox�{��}����* (&�w�u��        8F_��ϫ���@Q�,�l�뮻FE�*            �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��       �v�X    `���4vG   � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �  Ԯ�6 �h ���T���,Sĕu�@�'pg���8        �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��~�y�_˲� �<ϗ       ��^��x <�i�~O��~Ǿ��[>         /c۶�[> ���           $��k����    IEND�B`�PK
     �)K[��n  n  /   images/98e53ca1-f8df-492e-a5f5-3061f52364da.png�PNG

   IHDR   d   �   +n/�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��io[U��Wl'q�fh�6miZ(P(C�2�|x��
�*\^!U�B|������ $�2�I@�g(3�<�i�$�<��ݿm/�4��Nb;��U�:�9�׸�^۷v�Z	����as�J|*0���o��Y�FNt
��[�1m_��?(}Q>P y�2�I�2��d��0��a�$�(H�Q��< Fy@2��d��0��a�$����SOɓO>)Ӧ�1���/((���By�g�D���!x������<�hKKK�u����TWWK �/�A�_��|�/F#�x�
JKK�D�U�V�=z���s���/���<���E�Ge}��O���.�����r�9�șg�)ӧO�_�F��2�O�W��ϟ�ɕ��Ef@���� '������o�m۶�P�%<���򴵵Y ���3g��2(�P]��G���zc�� ����<>묳���[��w�{�C���t�M�b�
��@;O�!� GU=����7�xþf��E]$w�u��D�y��C��}��7KGG�lذA|xW��8��8r�<��#5��z����_����eƌqՔ�� :88h?��,..��<����ò<`䫗
�U܈�***�ꫯ����� ���#�������r��!�wsB<1<�e˖Y`���O(�Q#�{�n��?d������ky?/^,K�,��<s#@����R,@ ��_��_]�9b_}e:�mٲE>��+v�^{�}�D�xs��ak�qaǒqi�o������n��.���%ڀ�u�A��5��������k�9��ڱc������}�Q�n�:9x�\��8�r����s�=g�ǢE��s���)���q�mmm%��}��ɽ�������NXTT$?������L��>Y�`���w#F�����+	ut��y��g���ώ�/�Ђ�:��h6���>��o=Z7�D����nG<����=�!?L�%}��6�d��ZL�qګ��j���[��K/����!��������vl�駟�7Q�~����|�r����~���	I���g>��SH���x��N;�4��#�@%�p�裏�w��~�Ao
�{@
���ᤵ��V7�L����%����#�i�&�=JJJ����'*͍0�dxq�4���@PI���f����I֯_oG<��t�RkS���c^4�sҪ���u�jµ�`��/�l@E�}��V:b����Μ93> �'F���h�y<b�J�g#�l��Ih
��~+555�����7�6�-k	����u��D�H4¦&��� �JB��ro�n3�%�C��`?�s�o"��ƛ��pR� ����ܹs�n�AG{�z�68�(()�� �� ��_|1a��#%�\�*� �u�1�\`A��W�w�6���'�������/�8���� F�HU�@�͛'W]u���/�]����\S'|�y�g�ډj���ґ�(#��P1�P)�}T���'Su�o�ݺ��[���<`y4��	�0��裏�+��"�y_7"2_�j�̚5+)ҡ �t�v��dp8t^�kU�G�hpL��<���L��c�=&/���͆�#�{T�Xj<f�#�?��CV��k�ڵ블	7���f`w��ɂSQ90~�޽6�RCc#��jj�#Xm���=��q4��xnj#⻤����P�H�XUI��95̡ǳ�q+u4�{�6e���q��o�H�����Ǎm޼�zy���n���M��&���ß�)�g϶G�~s���d2��kll��L��ʄ/'�tR��Od�&\J�?� 8/�c2�����n�߄Yc��t:�q�Pka�atõ��7��T�s�ZhH���x�sq�\+��)��r�{\�x4Ƹk{�m a8*f�ƍ�@j�NrdN�<���eV���5Sf�AQkF^yY��N�F���_::�䰑��C����Ez��#��B�0#Q�ؙ�J�+L�2���E#����Q�,np��`�a���e�YK�43�j���Q������2��2��a^
T�6��J�4̑�b����a���l���wȠyn%J�͇�3~��6͚�L�I�(3��O?ّ�TM#L#�/�@�_|�̬��ζViڹU6:(�248��Q���{
�WX$e�RS7S�<�t�	�ɮ��rd`� � �R���[���Λ�)��7Jf�:$5�j��������/)/.��[7��쐞��F�cm�S��Q� ��~T:����l_(�J�>���A9�;$�<��ະae
 *ݩ���`|��W֋rf����"�,�V"��e���d���� �����{b�|pN{d�%2��H�t�38q a���V���⊈�.J �����TQH��r�,�.�B�G�6J��	�`T'���3�,/�ș�e��{P{�1��T3�H��S}�F�/��b� c4�߂�2i�*������_Zp4@C�_J|���/((OXRv��i#~���	"�Ci��۳g�5�c��)5e2Ϩ��y5*-�J��k������V�l$L�QA�r@{�׿��kk #	?É��K�'a�f��k)���Ԑ�*	��Rm�S7�\<�AUU��܊i�V�`(q]uFR��h��5�H
e�����ȓ�kQ0 �ʸ���L,5���I�p@Z��#���@�I��J H�C�y)��3#nQm�}�fn�/��{( ��p^��r$$u�A*(e�  �z���o��3��@����{^E����鳪�()q+M�����cS�"�>�̭,�h�P
��|s߰t�=AJ�:<��#�}�)%� �='f��C�7#/��@�Po�I�P([���$e���$%�0��t� =�bVyqVH��y��'e&��ZՅ=dS�P�MI�Y��Ө-��ߨ�l"X�nTW����s�X�46�0�V[)��w��|��7����H��_u�O��Bb�O�d������P�2��}�4��h�I�%��*1*�g$h]`@���E2)%6�Y��+/�I��@�K����t��H�V�$���ǩ��d�9<fl$;�VJ<�{�'����${�$��p�\$ӡ�쇉?
�Y
E�Bj�+#��v��{c�j��2ɤ�K�h-ģ��l&��A5B���2��:�P,����<����hVˈ���pd��{LE�$��۲�l�e��6��7�#���&��$���H�>���[2�QH*԰�������@ h�

}٫�
B�;��үS��kcG�gP�;lt��X��
̠
�0ނ!  #�Z�.!�w8���%������did��S�:l���= F��TBXA�n�5����������30hT�h�����(���2�c��r���=��/���2�B� �%T�3�2>�9׏P}���/��[����0e���c۱:d�ɤ�KEJ�]Qe]Ds}C#���'��*�M�.Hl��!i�鋬[�5�1+�� BA˸��eDy�>���!��+%��&�utK�qL�U��V�H�SQ4���2�|;�������]�i���,��=-!�HS������J$�h��ֶV9`�dѬ�22��6H����FB���*��XYU� =
�c*4Q:+v78,3��O��փGl�)��d؏TUç�r�~��!�k���=��"�����9u6��d"_u��K��f �,{H��[��dPJ�(�� &aޠ���o{�dn�4)-.��
�Y��Ws�d|���6�r�HJ��ѷt1`1����
i;�.w7ʕ�J���Ǿ&i��^``?h�Ò��p�x$g�q�]9 ���<�*3*�dɼY��|��E���;o�� ׍!�+C�WR�|}��H	�-R�4m��(�b�o�|���d�v��w���VK(�`���A)Dq,��=9��Lp���|�u�\m���)0:���-�lv��o�����0J�C��nA,��(~`xX>۴S�0�d���)5�j�/��ξ�H��8�A�tu�N�*\n7�!Z�
�����7�e'ϓ�s�lf%]ޗ��3�^�o�97�/'���Ő��y@Zpc,1V#���������+�Ε2��.M%,0~hĸ�����f;l!����%�\bU�xvJ��1mt��� �
3o��P�4wt��sda]�-
��J���1��O�V��0�ל.J{��A�#Q[�π�=0h��n���"g̝)sk�I����:�x���oj�-�Hc[�Mr��$H-�ߍ7�hw����@S�Hk��O�%�۠kK�FCk��������D̨��T��m�����F����#�����t��fm[���Æ["��_$��Q�>�[lLi�,n���l��Ma�.��X�f0�����(] �+ʤ��T*K�RRTh��Z'��a�g$�hO���xN8����x"�PQl9���=���N���ʋ�ԛ�h#)���lS��vx`�g[�zCK���C�CxG�0@�ZC"F�Փ�v�M�z}�c-c��'���������Pg�Ήxg	���H}�Z(4�pɄN�ŝ~�u�u�YF
�x�W�Ą��Q58 �1��nq���g+8H�o�ħ��I��������9���DS.q�޹tc���/m_D�Fps������W^iG��<�E��k��L#}�9YhI�E�m�H[h0f�Z��m�)=�^��d	o��}j��U�!�(���&��`L@`8K��>�7C� �Z0�xK�n�ak�׉�2
�#�d#F+��1H+��Vm�1p`�Y
���&� ��-a����=2o����ZF��O�g�F��Uu�7Dʈ����J���6c��p� I���РF��n2�;+��E�u���
��DM(s��%��*����o�۳U�4J��1jv얂��޲�wi5�!ZL@�L0�w�y�e
���F{��=�$������.���s�F�����B���-�!�n�Arcm)F@ ��5����21ʈ(I9Fs*����v�`����R��ڦ�-qZܺ
E�T�Am���]�=����v�A5 &�-�@訊M��@�F�RC���嶥`�]�Hc`� l���q�}N�H��%�梨 y����d��5G����s�v�7��q�]�
ށn���xQ��-���X'�8!���d&ݤˡu�F\\T���`g�`�"���m�Ǩ*�7��0��܉�Ts�TB�d�(6�$��r�U	IB�%�m�G��������%�7�R��%7U�.�x���7ri�6�|9l?ՐO��3n��� D��b 0Q"e��sIm�ц7ZH>b�>a@���B6Q@k���b̝I�k≐��O2���S;�m���?�1��⫉n)HP�vn�k�/�X�º�L%J�i���p�	�'��۫1I"D��ʕ+cnH�3��f�5u��#��X�tH,�o I6ܹ\2�c�{�~W�^-�֭�Y�x�d i'7�<�8ad�1[{���(� �(��G�D�p$�	$#��P�_�B�ސ!Fs���e�5�{2F#���c3.MiG#��a���q��y��)��6#iJ��	��0��&��0��i�h�g.}�z��bef�=�R��^�6�D&����Lx��0���A�|$ ��z������]ɗM4�I0-a��^���K/ى�B.{H�D�ԟ�4�}�v�iY�p��b+��P^�KZ����y���T�x46�L�9�ׯ��)�ݱ[�:~�Ɉ�_���m���d;��}�����=�*��۶m�h^f!��[���r���������:��ۺ�/��w�o��<���:;;�� �f�V�}�RM��K�����gÆ?c�!�K�e�He�s3y72�an@wL>�)\��͹!&������ O?���/d͚5r��ڵk��q�NJ����[�韔$�(H�Q��< Fy@2��d��0��a�$�(H�Q�#' �M��S��iR|q�g���c<*I�s'1I��;��w\e���7㳑Y��    IEND�B`�PK 
     �)K[3��C� C�                  cirkitFile.jsonPK 
     �)K[                        p� jsons/PK 
     �)K[Ȣ                 �� jsons/user_defined.jsonPK 
     �)K[                        H images/PK 
     �)K[tM�G.  G.  /             m images/cac5f02b-fb1b-403b-a5d1-1baa7913483a.pngPK 
     �)K[]�I��  �  /             L images/898fbbe1-f190-4098-9ff7-64122b8b80b8.pngPK 
     �)K[�wp�&
  &
  /             '[ images/1cdb40d8-22d5-4761-8204-85ee5f97d036.pngPK 
     �)K[!��Ů  �  /             �e images/9ee875d8-7c7b-435c-a3d9-92ac29f03ab9.pngPK 
     �)K[�c��f  �f  /             �h images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.pngPK 
     �)K[��EM  M  /             �� images/d3694a2e-5bba-40c3-8069-8db85c4c9209.pngPK 
     �)K[	��} } /             ]� images/bbfae99c-8036-4c5e-89fd-a87441410720.pngPK 
     �)K[d��   �   /             �` images/a262aa33-74c4-460b-b0ad-c746896f6744.pngPK 
     �)K[:\�iE E /             �� images/7be072cc-a725-4446-be13-eff8a797d760.pngPK 
     �)K[��R�(  �(  /             &� images/d39a4f5b-af2c-4f90-bee3-bb82593c1b3b.pngPK 
     �)K["1^FHo Ho /             C� images/6b6fcb51-98f7-4a52-b90f-3140c0078893.pngPK 
     �)K[��n  n  /             �* images/98e53ca1-f8df-492e-a5f5-3061f52364da.pngPK      G  �C   