PK
     ��d[M8�  8�     cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_0":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_1":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_2":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3":["pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1"],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_4":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_5":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_6":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_7":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_8":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_9":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_10":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_11":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_12":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_13":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14":["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1"],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_15":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_16":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_17":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_18":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_19":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_20":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_21":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_22":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_23":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_24":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_25":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_26":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_27":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28":["pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0"],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_29":[],"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_30":[],"pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0":["pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1"],"pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1":["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14"],"pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0":["pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0"],"pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0":["pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0"],"pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1":["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3"],"pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0":["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28"]},"pin_to_color":{"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_0":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_1":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_2":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_4":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_5":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_6":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_7":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_8":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_9":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_10":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_11":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_12":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_13":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14":"#ff0000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_15":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_16":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_17":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_18":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_19":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_20":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_21":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_22":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_23":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_24":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_25":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_26":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_27":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_29":"#000000","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_30":"#000000","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0":"#000000","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1":"#ff0000","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0":"#000000","pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0":"#000000","pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1":"#000000","pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0":"#000000"},"pin_to_state":{"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_0":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_1":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_2":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_4":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_5":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_6":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_7":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_8":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_9":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_10":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_11":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_12":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_13":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_15":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_16":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_17":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_18":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_19":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_20":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_21":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_22":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_23":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_24":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_25":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_26":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_27":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_29":"neutral","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_30":"neutral","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0":"neutral","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1":"neutral","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0":"neutral","pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0":"neutral","pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1":"neutral","pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0":"neutral"},"next_color_idx":27,"wires_placed_in_order":[["pin-type-component_a3ae65d4-c858-4cbe-bb67-1538767c17f8_5","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_7"],["pin-type-component_a3ae65d4-c858-4cbe-bb67-1538767c17f8_7","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_8"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_29_polarity-pos"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_13","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_28_polarity-neg"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_29","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_29_polarity-pos"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_28_polarity-neg"],["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_1","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"],["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_0","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16"],["pin-type-fake_0","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16"],["pin-type-fake_1","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"],["pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_17","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16"],["pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_12","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"],["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_0","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_1"],["pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_0","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_1"],["pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_0","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_1"],["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_1"],["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_1","pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_1"],["pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_1","pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_1"],["pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_1","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1"],["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0"],["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_1"],["pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_1","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_1"],["pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_1","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_1"],["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_1","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_1"],["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0"],["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0","pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0"],["pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0","pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0"],["pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0"],["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_7","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_0"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_8","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_0"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_9","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_0"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_10","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_0"],["pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0"],["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3"],["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0","pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0"],["pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28"],["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0"],["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_5"],["pin-type-component_b00b0f46-5dcc-4451-a676-221697210905_0","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_4"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_19","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_6"],["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_16","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_7"],["pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0","pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0"],["pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3"]],"wires_removed_and_placed_in_order":[[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_a3ae65d4-c858-4cbe-bb67-1538767c17f8_5","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_7"]]],[[],[["pin-type-component_a3ae65d4-c858-4cbe-bb67-1538767c17f8_7","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_8"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[["pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_7","pin-type-component_a3ae65d4-c858-4cbe-bb67-1538767c17f8_5"]],[]],[[["pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_8","pin-type-component_a3ae65d4-c858-4cbe-bb67-1538767c17f8_7"]],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_29_polarity-pos"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_13","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_28_polarity-neg"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_29","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_29_polarity-pos"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_28_polarity-neg"]]],[[],[["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_1","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"]]],[[],[["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_0","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16"]]],[[["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_0","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16"]],[]],[[],[["pin-type-fake_0","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16"]]],[[],[]],[[["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_1","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"]],[]],[[],[["pin-type-fake_1","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"]]],[[],[]],[[["pin-type-fake_0","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16"]],[]],[[],[["pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_17","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16"]]],[[],[]],[[["pin-type-fake_1","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"]],[]],[[],[["pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_12","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"]]],[[],[]],[[["pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_12","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_15_polarity-neg"]],[]],[[["pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_16","pin-type-breadboard_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_17"]],[]],[[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_13","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_28_polarity-neg"]],[]],[[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_28_polarity-neg"]],[]],[[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_0_29_polarity-pos"]],[]],[[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_29","pin-type-power-rail_295e808d-80c9-46a1-9a2f-f0256ea548ee_1_29_polarity-pos"]],[]],[[],[["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_0","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_1"]]],[[],[["pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_0","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_1"]]],[[],[["pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_0","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_1"]]],[[],[["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_1"]]],[[],[["pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_1","pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_1"]]],[[],[["pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_1","pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_1"]]],[[],[["pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_1","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1"]]],[[],[["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0"]]],[[["pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_1","pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_0"]],[]],[[["pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_1","pin-type-component_58c69d60-1524-404c-a65b-4620d583a77a_1"]],[]],[[["pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_0","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_1"]],[]],[[["pin-type-component_22d00f1f-0745-486c-8cd6-bfd25d6b5e47_1","pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_1"]],[]],[[["pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_0","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_1"]],[]],[[["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1","pin-type-component_dc601ec5-59fc-466a-95c6-ea5efbf86d55_1"]],[]],[[["pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_1","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0"]],[]],[[["pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1"]],[]],[[],[["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_1"]]],[[],[["pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_1","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_1"]]],[[],[["pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_1","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_1"]]],[[],[["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_1","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_1"]]],[[],[["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0"]]],[[["pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0","pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0"]],[]],[[],[["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0","pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0"]]],[[],[["pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0","pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0"]]],[[],[["pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0"]]],[[],[["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_7","pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_0"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_8","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_0"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_9","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_0"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_10","pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_0"]]],[[],[["pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0"]]],[[],[["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3"]]],[[],[["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0","pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0"]]],[[],[["pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28"]]],[[],[["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0"]]],[[["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3"]],[]],[[["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1"]],[]],[[],[["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_5"]]],[[],[["pin-type-component_b00b0f46-5dcc-4451-a676-221697210905_0","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_4"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_19","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_6"]]],[[],[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_16","pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_7"]]],[[["pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_10"]],[]],[[["pin-type-component_07201ce6-242e-4070-beb1-6b1ecc8e9a32_1","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_1"]],[]],[[["pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_9","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_0"]],[]],[[["pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_1","pin-type-component_f7b311cb-2dd2-4362-af91-c7568e208d66_1"]],[]],[[["pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_8"]],[]],[[["pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_1","pin-type-component_c059b081-dcbb-437e-bb8b-813da336182d_1"]],[]],[[["pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_7"]],[]],[[["pin-type-component_4d0af7ef-6915-4a65-b658-362c305c51f1_1","pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_1"]],[]],[[["pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0","pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0"],["pin-type-component_8bc6f0d9-3ee0-4f84-84b0-8d65a769c427_0","pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0"]],[["pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0","pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0"]]],[[["pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0","pin-type-component_9d6a5121-9e9a-495e-ba64-f8cf5049df87_0"]],[]],[[["pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0","pin-type-component_68792fb0-2eb6-44eb-88c3-d5bd97335509_0"]],[]],[[["pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0","pin-type-component_5bff362d-8f79-4a23-b1e8-04253d472f65_0"]],[]],[[["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3"]],[]],[[],[["pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3"]]],[[["pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_4","pin-type-component_b00b0f46-5dcc-4451-a676-221697210905_0"]],[]],[[["pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_5","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14"]],[]],[[["pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_6","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_19"]],[]],[[["pin-type-component_0232f75e-f080-4dd3-8137-8958c98da454_7","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_16"]],[]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_0":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_1":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_2":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3":"0000000000000009","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_4":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_5":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_6":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_7":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_8":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_9":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_10":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_11":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_12":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_13":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14":"0000000000000010","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_15":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_16":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_17":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_18":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_19":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_20":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_21":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_22":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_23":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_24":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_25":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_26":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_27":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28":"0000000000000011","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_29":"_","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_30":"_","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0":"0000000000000009","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1":"0000000000000010","pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0":"0000000000000004","pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0":"0000000000000004","pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1":"0000000000000009","pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0":"0000000000000011"},"component_id_to_pins":{"f0fd6315-2925-41b3-9764-248681cdce0c":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30"],"636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35":["0","1"],"2829c8e4-4312-47ed-a029-8eab57667ef2":["0"],"28debeb4-25ba-40b7-880d-a84ab194857a":["0","1"],"a21c1a89-038d-4d33-9463-f2151579a9e0":["0"],"e87dc4da-e2d8-41cc-bc12-69ed72c01d9e":[],"d710e40b-242b-4d55-aff1-d25d4416cf71":[],"b1be3c37-6458-4463-9c21-0cddf8035423":[]},"uid_to_net":{"_":[],"0000000000000004":["pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0","pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0"],"0000000000000009":["pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1","pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3"],"0000000000000011":["pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28"],"0000000000000010":["pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1","pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14"]},"uid_to_text_label":{"0000000000000004":"Net 4","0000000000000009":"Net 9","0000000000000011":"Net 11","0000000000000010":"Net 10"},"all_breadboard_info_list":["bf214f1e-c792-43f5-846b-d34128e4e83a_30_2_True_955_100_up","bc941250-d2ab-4f36-99ca-60371a583e71_63_2_True_835_10_up","295e808d-80c9-46a1-9a2f-f0256ea548ee_30_2_True_940.5_145.49999999999955_right"],"breadboard_info_list":[],"componentsData":[{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"161","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"Adafruit Industries","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[625.654174,295.80002],"typeId":"84ae97c1-8e69-5e6b-4fa6-dfe46d477633","componentVersion":1,"instanceId":"636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35","orientation":"up","circleData":[[602.5,305],[648.8083479999996,305]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[453.1307005000001,383.442893],"typeId":"98d6e125-552a-4063-90e5-58c04872effd","componentVersion":1,"instanceId":"2829c8e4-4312-47ed-a029-8eab57667ef2","orientation":"up","circleData":[[452.5,365]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"10000","displayFormat":"input","showOnComp":true,"isVisibleToUser":true,"name":"Resistance","unit":"Ω","required":true,"validRange":[0,70000]},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.25%","value":"0.25%"},{"label":"0.1%","value":"0.1%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false,"isVisibleToUser":true,"name":"Tolerance","required":true},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"string","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false,"isVisibleToUser":true,"name":"Number Of Bands","required":true}},"position":[502.22504875383447,305.69373781154127],"typeId":"72c75556-baa3-04e7-55a5-e13f447c8c5a","componentVersion":1,"instanceId":"28debeb4-25ba-40b7-880d-a84ab194857a","orientation":"up","circleData":[[467.5,305],[542.5,305]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1008.1307005000001,383.4428929999999],"typeId":"98d6e125-552a-4063-90e5-58c04872effd","componentVersion":1,"instanceId":"a21c1a89-038d-4d33-9463-f2151579a9e0","orientation":"up","circleData":[[1007.5000000000001,365]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"5v dc","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[688.5146147612892,322.037732766394],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"e87dc4da-e2d8-41cc-bc12-69ed72c01d9e","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"5v dc","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[891.2520860259777,419.8110375396785],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"d710e40b-242b-4d55-aff1-d25d4416cf71","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"GPIO34","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[693.7762858314251,242.75732919044282],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"b1be3c37-6458-4463-9c21-0cddf8035423","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[803.2100499999999,309.8848895],"typeId":"5dd9522a-ac85-4cae-b2c3-8ba3fec8b601","componentVersion":2,"instanceId":"f0fd6315-2925-41b3-9764-248681cdce0c","orientation":"left","circleData":[[752.5,230],[751.6624749999999,240.99967700000002],[752.7453145,250.29215899999986],[752.1075655,261.7580989999999],[752.3877774999999,271.7645255],[752.5665445,281.7735544999998],[752.5665445,291.86251249999987],[752.1075655,301.8715924999999],[753.0255249999998,311.49889699999983],[753.5859504999999,321.96691999999985],[752.5665445,332.78988649999985],[751.9287969999998,342.6227749999998],[752.8467579999997,353.5204279999999],[753.4845054999998,362.90210149999996],[753.4845054999998,373.2634804999999],[854.4709314999998,230.39584999999988],[854.4709314999998,240.90942199999995],[855.060628,251.10101299999997],[854.5456779999997,261.6919805],[855.135376,272.437451],[854.7284064999999,281.4854839999998],[854.3214354999998,292.41885049999996],[854.063962,302.0928889999999],[854.7284064999999,312.6888079999999],[854.8819884999998,322.9092259999999],[853.6610784999998,333.63743599999987],[854.4445854999999,343.0979329999999],[854.8819884999998,353.7271684999997],[854.0680494999999,364.2397129999998],[854.851555,374.5201729999998],[804.8739519999999,408.6976309999999]],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"196.37686","left":"425.30875","width":"610.64390","height":"251.93417","x":"425.30875","y":"196.37686"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0\",\"endPinId\":\"pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0\",\"rawStartPinId\":\"pin-type-component_2829c8e4-4312-47ed-a029-8eab57667ef2_0\",\"rawEndPinId\":\"pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"452.5000000000_365.0000000000\\\",\\\"452.5000000000_305.0000000000\\\",\\\"467.5000000000_305.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1\",\"endPinId\":\"pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0\",\"rawStartPinId\":\"pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1\",\"rawEndPinId\":\"pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"542.5000000000_305.0000000000\\\",\\\"602.5000000000_305.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1\",\"endPinId\":\"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3\",\"rawStartPinId\":\"pin-type-component_28debeb4-25ba-40b7-880d-a84ab194857a_1\",\"rawEndPinId\":\"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"542.5000000000_305.0000000000\\\",\\\"542.5000000000_261.7580990000\\\",\\\"752.1075655000_261.7580990000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0\",\"endPinId\":\"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28\",\"rawStartPinId\":\"pin-type-component_a21c1a89-038d-4d33-9463-f2151579a9e0_0\",\"rawEndPinId\":\"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_28\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1007.5000000000_365.0000000000\\\",\\\"870.7840247500_365.0000000000\\\",\\\"870.7840247500_364.2397130000\\\",\\\"854.0680495000_364.2397130000\\\"]}\"}","{\"color\":\"#ff0000\",\"startPinId\":\"pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1\",\"endPinId\":\"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14\",\"rawStartPinId\":\"pin-type-component_636bd1e9-d2a6-4f1b-9edb-25dbdd21dc35_1\",\"rawEndPinId\":\"pin-type-component_f0fd6315-2925-41b3-9764-248681cdce0c_14\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"648.8083480000_305.0000000000\\\",\\\"730.0000000000_305.0000000000\\\",\\\"730.0000000000_372.5000000000\\\",\\\"753.4845055000_372.5000000000\\\",\\\"753.4845055000_373.2634805000\\\"]}\"}"],"projectDescription":""}PK
     ��d[               jsons/PK
     ��d[��+��,  �,     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"Photocell (LDR)","category":["Input"],"id":"84ae97c1-8e69-5e6b-4fa6-dfe46d477633","subtypeDescription":"","subtypePic":"b63deb06-c33f-4ae3-8f73-25229955b1c1.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.58334,76.55539","endPositionMil":"14.58334,14.58330","isAnchorPin":true,"label":"pin 0"},{"uniquePinIdString":"1","startPositionMil":"323.30566,76.55539","endPositionMil":"323.30566,14.58330","isAnchorPin":false,"label":"pin 1"}],"numDisplayCols":"3.37889","numDisplayRows":"1.51833","pinType":"movable"},"userDefined":false,"properties":[{"type":"string","name":"mpn","value":"161","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Adafruit Industries","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"a5640015-ff5c-4848-bb8b-6d4b42e5489b.png","componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"GND","category":["User Defined"],"id":"98d6e125-552a-4063-90e5-58c04872effd","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1cdb40d8-22d5-4761-8204-85ee5f97d036.png","iconPic":"9ee875d8-7c7b-435c-a3d9-92ac29f03ab9.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"2.37626","numDisplayRows":"3.61380","pins":[{"uniquePinIdString":"0","positionMil":"114.60833,303.64262","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Resistor","category":["Basic"],"id":"72c75556-baa3-04e7-55a5-e13f447c8c5a","subtypeDescription":"","subtypePic":"bbfae99c-8036-4c5e-89fd-a87441410720.png","userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[{"type":"double","name":"Resistance","value":200,"unit":"Ω","showOnComp":true,"required":true,"validRange":[0,70000]},{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}],"iconPic":"a262aa33-74c4-460b-b0ad-c746896f6744.png","componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"GND","category":["User Defined"],"id":"98d6e125-552a-4063-90e5-58c04872effd","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1cdb40d8-22d5-4761-8204-85ee5f97d036.png","iconPic":"9ee875d8-7c7b-435c-a3d9-92ac29f03ab9.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"2.37626","numDisplayRows":"3.61380","pins":[{"uniquePinIdString":"0","positionMil":"114.60833,303.64262","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"ESP32 (30 pin)","category":["User Defined"],"userDefined":true,"id":"5dd9522a-ac85-4cae-b2c3-8ba3fec8b601","subtypeDescription":"","subtypePic":"f51f6ed9-d8f0-454d-af8a-e11415a94f15.png","iconPic":"53dea2ad-2eb7-451c-84a6-1b4fef66a2aa.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"13.80107","numDisplayRows":"7.59928","pins":[{"uniquePinIdString":"0","positionMil":"1222.61943,718.03100","isAnchorPin":true,"label":"EN"},{"uniquePinIdString":"1","positionMil":"1149.28825,723.61450","isAnchorPin":false,"label":"VP"},{"uniquePinIdString":"2","positionMil":"1087.33837,716.39557","isAnchorPin":false,"label":"VN"},{"uniquePinIdString":"3","positionMil":"1010.89877,720.64723","isAnchorPin":false,"label":"D34"},{"uniquePinIdString":"4","positionMil":"944.18926,718.77915","isAnchorPin":false,"label":"D35"},{"uniquePinIdString":"5","positionMil":"877.46240,717.58737","isAnchorPin":false,"label":"D32"},{"uniquePinIdString":"6","positionMil":"810.20268,717.58737","isAnchorPin":false,"label":"D33"},{"uniquePinIdString":"7","positionMil":"743.47548,720.64723","isAnchorPin":false,"label":"D25"},{"uniquePinIdString":"8","positionMil":"679.29345,714.52750","isAnchorPin":false,"label":"D26"},{"uniquePinIdString":"9","positionMil":"609.50663,710.79133","isAnchorPin":false,"label":"D27"},{"uniquePinIdString":"10","positionMil":"537.35352,717.58737","isAnchorPin":false,"label":"D14"},{"uniquePinIdString":"11","positionMil":"471.80093,721.83902","isAnchorPin":false,"label":"D12"},{"uniquePinIdString":"12","positionMil":"399.14991,715.71928","isAnchorPin":false,"label":"D13"},{"uniquePinIdString":"13","positionMil":"336.60542,711.46763","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"14","positionMil":"267.52956,711.46763","isAnchorPin":false,"label":"Vin"},{"uniquePinIdString":"15","positionMil":"1219.98043,38.22479","isAnchorPin":false,"label":"D23"},{"uniquePinIdString":"16","positionMil":"1149.88995,38.22479","isAnchorPin":false,"label":"D22"},{"uniquePinIdString":"17","positionMil":"1081.94601,34.29348","isAnchorPin":false,"label":"TX0"},{"uniquePinIdString":"18","positionMil":"1011.33956,37.72648","isAnchorPin":false,"label":"RX0"},{"uniquePinIdString":"19","positionMil":"939.70309,33.79516","isAnchorPin":false,"label":"D21"},{"uniquePinIdString":"20","positionMil":"879.38287,36.50829","isAnchorPin":false,"label":"D19"},{"uniquePinIdString":"21","positionMil":"806.49376,39.22143","isAnchorPin":false,"label":"D18"},{"uniquePinIdString":"22","positionMil":"742.00017,40.93792","isAnchorPin":false,"label":"D5"},{"uniquePinIdString":"23","positionMil":"671.36071,36.50829","isAnchorPin":false,"label":"TX2"},{"uniquePinIdString":"24","positionMil":"603.22459,35.48441","isAnchorPin":false,"label":"RX2"},{"uniquePinIdString":"25","positionMil":"531.70319,43.62381","isAnchorPin":false,"label":"D4"},{"uniquePinIdString":"26","positionMil":"468.63321,38.40043","isAnchorPin":false,"label":"D2"},{"uniquePinIdString":"27","positionMil":"397.77164,35.48441","isAnchorPin":false,"label":"D15"},{"uniquePinIdString":"28","positionMil":"327.68801,40.91067","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"29","positionMil":"259.15161,35.68730","isAnchorPin":false,"label":"3V3"},{"uniquePinIdString":"30","positionMil":"31.30189,368.87132","isAnchorPin":false,"label":"USB POWER"}],"pinType":"wired"},"properties":[],"componentVersion":2,"hasComponentImageSvg":false,"componentImageSvgUrl":""}]}PK
     ��d[               images/PK
     ��d[��F�} �} /   images/b63deb06-c33f-4ae3-8f73-25229955b1c1.png�PNG

   IHDR  �  D   CzWF   sBIT|d�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<    IDATx���{��y^�'�U�Y�s�����xYD�F@P��;�Ჱ�ll쮷]5aa�V$��uB�n�0ܼ��������,������Ow�S��2뒷�#+�T�S��\��WY��Dd����'�'N�y�����   @�	I~>�J   `!���3�<S:   eUK   ��OK��(�   P�S��zs�    ���  ��ޒ�g�|b�     ,�7$��$�[:   �(�  ,�?��ǒ\-    �'y_��(  �2j�   P�W%yg�V�     p�F�/O�����  �9Sp  X<_���'��    �QM�G29�����   p��  G%��M��    p�U�|v�ߐ䇒���  �<(4   ,�z��L򕥃    �#xO��%9(  ����  p��d2�ꭅs    ����$_�d�t   Ύ�;  ��v=ɏ'�=��    �)��$_����A   8
�   ��'&��I>�t    8E�$��I>\:   ��Z:    g�w'��Qn   ����$?��3J  ��)�  \>oM�I^W8    ���I�M�/(  ��U+   �S��$ߟd�t    8cK�{6�*�  �S��  py��I�i�f�     pNjI�x�^��+�  �S��  p9��Ç�   �h*I�p�V�S8   �I�  `�}K���ɉ<    XD�$oI�II�[6
   �C�  `~U���$�t    �@~ �ےJ  ��)�  ̧z�wfr�    8�}I�<�A�    <w  ��SO�I��t    ���]�/N�+�  ����  0_���7��    s�?fr,m�t   ��;  ��XI�I�R:    ̑&��$/�  �kSp  �kI~<��/    �Ї3)��z�    �:w  ���$�6��(    �سI>7�ӥ�   p��   xUoJ�3Qn   ���	I~.ɛK  ���  .�OL�I~K�     pI<��'��g��   p2w  ���S��?�o.    .�k����@�    �K�  ����I~&�[&    �o-ɏ&���A   8N�  �b�=I�M��J   �Kn5ɏ$����   p��;  ���Ln�|�t    X�$?�䏗  �D�t    �$_��2�    ��z�/O�t�_*�  `�)�  ���I�?�iQ    ���e2�]�  �0w  ���d��I�T:    ,�Z&��>��g  XX
�   �L����A    �$I5�I�J�   �(�  ���    ��;  @A
�   ��OdRn_*    8��;  @!
�   �K�    �C5ɗ$�p��  ΍�;  ��Qn   ��R�d���;  �9Qp  8_����,�    <%w  �s��  p��0�&i�    <�i���$�T8  ����  p�� �r{�t    �LK���;  ��Qp  8;��    p�Ԓ��(�  �w  ��񇓼'��    p�(�  �!w  �ӧ�    �۴��kI>X8  ����  p���   `1(�  �w  �������;��     �B�  ��)�  ��v    XLJ�   �H�  ��)�   �bSr  8%��   ���&��$��A  NK��H�ٜ���jY^^>�O�s�ھ���T���륥����{�ܥ�����Z���۫�jZ��}�W*��ۧ���~��888H��?�?ooo/���^����� {{{�֍F����[���������h4�o��`������\ �9t��O%yo�    �J�  ����$�:�z�  @9��˩�j���G�V+�J�XI��l޳=9�P}R��V�ssΓ��GK��j����џ��\F����=%��_���e0�^��^��ce�����*�O�?Z���ߟ�����?��E�n�a>6 p��%��$?Z:  �<Rp  x4�=ɿKr�p ������=e񥥥Y�{Z����l?Z@����I�z�~��>��ۛ�f�ƙv`��P�����p��x<+�-�O�G�G�?-����������t���?}�i�=  ��n�/N�S��   �w  �����L�7� �mZ�>߽<�>�P~�>�{��<�}&���~�?+�O�f������|������y�t���� � v���$?[:  �<Qp  x8o���'� �"x�ݞM,�N+�N:�N_^^N�Z��?�����d�ݯ�qMK��i�w�~��$���I�t�����i����f8foo��G��[I>/�J  �
�   �Z��'���A ��f3�Ng6�|�|t��t���������3�|� xu���t�|�׻gB}�۽g:�t�`0����=S鷷�3J< ��+I�P�_,  `(�  <�+I~*��(�ӳ���f�����,//�^���j���N'�z=KKK���v{V@o�Z���'m .�i�}ww7��`6I~0�����g?{{{������z�{�3-����Ϧ�pi��䳓|�t  ��N�  �u��D��(`ѝ4��t�N�s�4����v�=������Z�V�# �׫M��N��n�{J����l�t���݌F��`�}4�<|  �>�  ^�R���t% ´H�l6�n�ge󥥥c��ѧ�ޯ� �㙖ޏ��f��"�����b���M_�P>�I����A   .*w  ���'yO�/.༴��,//��j��jeyy9�v{�z���j���dyy9��˳������ ���������������eoo/�����z��ݝ=�ۺ��׻���}M�ȯdRr�t  ��H�  �d�$�J򕥃 <���v�=�����2��~����������Z���(  ,��t�����S�N�?i����́$��$ۥ�   \4
�   '�'I��t�r�V��I�G��O�����cէ�wOTo6��?
  \�~6!~gg�ش�����z��z�ٺ�������f8��(����I>?�^�    ��;  ���A�?_:p�M'�7��٤����O���G�]__O���  \D��(����&������l�۷og4������I�8��j   9�
  p��&��J� �G�ٜ�ϧ��z�>[wA���z��(�  �lZx?� �<t�ty{{;����G ���%y[�q�    ��;  �-�7�<������GK��v;�v;�V+�N'�Vk�  �"������nz�މ��'�O���g`��#�W�  p(�  L�wI�a�j� �hN��~wY�u  ���j��.�����F���a��I��t  ���  �?��;��J�y��%���������  �ˣ�㷶�2KǇy5��.��\:  @I
�  ����I�/I�t(�R��J����-]�n�S�8�   ���������3{L_O��G�����$_�䟕  P���  �"{K�K�)N��&�oll�ʕ+'NS_[[K�Z-  �� S�oݺ�����>������i$�ϓ�`�    %(�  ��%��$�J�W����������euuu65����N'����t\�  ��x������������v������[:6���$_��'K  8o
�  �"��$�w�7����t:���x���W�\I��.   .�n�����{��O��O�O��ߺu�td�f��N򋥃   �'w  `�\M�I>�t�_�����F666f���$��֯���R�Oq   �G�~?�nwVx������f677O\�֭���ұ�/&��$)  �8�  ,�N������j6��	�G'�}LK���   ����?�?]w�������ұ�x�N�I^.  �<8  ,�z��%���A8{G���b�݅��E�����j�ұ   f��i���+�-��z�ܾ};�Ѩtl��J�$;��   �5w  `T��;��J��4����fcc#kkkY[[��^]]=�����F�Q:2   ���F������N����������lmmekk+�oߞ��}�v���JG���D&<��   �%w  `|k���t�k6�������FVVVf��	�G_����R�OX   ��5���v���9�����N677s�������&��$��A   Ίv   p���$�t�E�l6��t�n�����+W�̊�W�\I�ݞٯ^��Z�V:2    ����+��z�ܺukV��.�z�ܾ};�Ѩt�E������!   Ί�;  p��Iޙ�Z:ȼZ^^���F���f����r�ʕ���fuu5���Y__O��,   ���A�������۷oϞ777�������ܾ};�o����N���o$���!   ΂�;  pY�5ɏ&Y.��»r�J��ַfuu5W�\��766��   8�2�t:���Vnݺ�_��_ȇ?������(�W%���A   N[�t   �3𻒼'���>��e_�e�c    �@��z�\��+W�[�h4�L5�?K�B�[8  ����   p�>1�'Y/d^����
   ��acc�t�y�L��I~G�    �I�  �L6��X�7�2O���JG    �$�U=��$�:�'�  pj� �ˢ��I~k� ��T,    .
Ǫ�SI~<ɕ�A   NC�t   �SPI�]I�`� �h}}�t ���V��T*��\�TR���y�I�ﻟ�h��x|���px��x��x<{߫= p~�zd���G��5�~�(   �G�  ��^��(b^��3 pT�VK�ZM�Z�-�j��.O���'��_��>��%��`��h��h��p��p8[�ߺ�2  fuu5�jՅ����g2�O%���O  �9��  ̻�1�_(b���3 \~���G�ZM�ј-���4�T*��q/�ii��l>������>2^u��I�  ��R�duu5�o�.e^}y�oJ��J  xT
�  �<�#I�n���m�`~-�O��G�^O�V�MV��J�2�o������-�������������� �e������x�J������A   �3  ��zs��I�hc4I�4��Z��1 �����~R����A����I��� `^mll��h���[�|4ɏ�  ��� �y�T��&Y+d�mll��  �R�+�7���s��L�Z-��V��V�eyy������X���� ���988H���x<>��  �OE#ɻ���$�_�,   E�  �7KI�e��P:�e��� 8k����>}LK�J�tD.�J�2���ݦ�����Y�}�|ppP - �q
�f#���|F��g  x`
�  �<�d2u���rY8Y ���4����,--��lfyy�$v.��*�O��O'�O�M} ΋cV�ꓓ�H��N�W8  �Qp  ��7'���!.'����>-�O���̻J�2���Q�� �yr�����$ߙ�O�  � � �y�g����!.����� �B�V�Y^^���R���g˕J�t48W�+��F�Y�}oo/{{{����h4*� ��:_���I�f�    �E�  ����%�$;eN��Z�X�}yy9�fS�^E�ZM��J�՚��{����^vww3& �cVg�o$y&�;J  x5
�  �E�[�|O�f� ���� ,�Z��V�u���h4JǂK�~��fޕ��W���^:�eUI��|8�O�  p_
�  �Ev%�%�Z:�e���"�T*i6�i�Zi��Y^^��x��f��f��u��� �^/������x<.� �(VWWS�V3�JG���I~ �g%���Y   N��  \T�$?��SJ��VWWKG �SW�׳���v�=��^�VK�NP�׳��6��r<g?�^/{{{��� �b�T*YYY���V�(��F��%��$��  pw  ���I>�t�����w�j�X���j�V���<�J�����,//������fwwwV|7� .���U���30�9I\Q  \(
�  �E��$�t�ˮZ�fee�t x(�B{��J��I��2�.�z������݇F�Q�������n����݌F��)�Ӷ����{�t����%��$_Y:  �Q
�  �E�UI�z�����(p�U���d�v��v��J�R:PP�Z��}p�ڵ����������eww7��tL �1������(ޖ�W�|C�   3
�  �E�$ߖD��8I�ET��f��v����%�v�UU*�,//gyyyVx���K��Sx�9��չ��$O'yg�    ��;  pq��$�I�*dQ8I�EP�T����N��N�cB;��*����wOx�Ny�ǥc �auu�t�ERM�$�&���Y   � �a#ɏ$�V:�"q��R�.�W�n����'��F�Yٽ�����tD ����#,��$ߗ��%y�p  `�)�  �U�|W�O)d�8I�y��j�B{��I��(	X`�j5����>�A��nvvv��v3' �
y"�'��I���   L�  (��%���!��� ��J��V�����t:�,//��gj��g���$�u:��j��0��z��׳����x����Y�}��+ p�g(�&yg�/-  X\
�  @I_��ϗ�����JG �9:�}ee%��C���x4�pg���8�����3�vg�L�g4���������~F������f��[7��I��#a�lo�?f��=��lo�3�Y�^O��~�}�'\�X?���I��VVR�V���tR=,��z_����v{V�-/��lN�7��^�R���|�J���u�\k�S��OL/�i�Z�~�z���쾳�c�; �#����I��$__:  ��.��c  `Q|f���R:ȢRp�q5�ͬ��dee%�v;��_�gaZ���L
�;;���{{�z����������x8����ϊ���-�O�ݣ�݌����2:8(���x0�`k��=q��;�DgoV��TR_YI2)ԧZMmy9�F�X�q���n'�ZjKK�.-M�?,��:�T��Z�T��&?��J�јl�VO��$�Z-kkkY[[�x<�����ׅ ��2����M�KI��t  `�(�  %�)�$Y.d����ÚN6^YY���j�����`{;����`k+���;��~���w
��nF�A�;;�"s�7{���x8�`kk6u|t�$s�lF��)�o���V'����;e����Z�T��YѾ��6+�ז�S]ZJke%K�zvG�����'���r}�ٜL�w� <�V��F���]w���T��#�/gRt  87
�  �yk&��$�+dљ�����j�t:Y]]���J��j�H�dtp�a��a����V��ެ|>�ޞ�lOZ���po/Ý���&��#�v`��F�I��[�%�=|��N��aٽ�nO��G
����Ia�p�}��J��Jm���N��N��u�p X$����y�f��l-�{�|z�!  �s��  ��o�������� �5-�O'��,��4������v�������ome��u|����d����J5I��1Τ��K���g��g����:�_m6Si4R�t&����T��f��k�v�N*'�wX��	� \p���
��}r��M�I���   B�  8O_��+K� �V�i�ۥc p��j����dmm-�N'��(=�4-}����wv2��ɠ�ͨכl�ٙ���s�0o*I�Ӳ�t��i4�F�~F�����Tj��d�Ng2M�՚=���;������]Z��M����������%��$�t  `1(�  ��O&�_J�`bmm�� \�z=���Y[[K�՚�n�zw��oo�ylme��3������t�ay}���a���`P��\G��9�����t��=]�R�Φ�W'�O���_��k�S;�0_�tN�� pY������1�J�/
�   ��;  p>5�?OR-������ 8c�~2�p���ͨ��xw7��0����z������E���n�Ψ�/�ҹ��~����Qv��hrW���Gz�ѸS~��_?,�O��G��WWS�;�p�9�u�T���$L�g  .9G�  ���I�t8� ������e��;+�����^F��d�����p�����po�؟UM�J�N����*� ��J&/��d�i�}T0W	�~?����77���VkR~o�'e�Ng��#    IDAT��p�zd�|�p����� s�1����=I>=��   ���;  p�*I�'�o+������L'�vv2<|�,�6{�v3>�<�j&��i��r
���wt��8��{7����`�y0���pw���W�VS;,��WWg����kw���Zg�	 x-&�_HoH�%��$n�  �	w  �,��$_\:�rr��L���^/���nݚMP��ܙ�~8i}���v2>���R&�OieRr`~-��2)����ڛxh��(������}�N'���cS�k�Τ ����]�I�%f �Ð��3���$�M�   ���  ��/I�5�Cp2�w�Ѣ���>������[���[[�F�����I����V8 ������$��)��������J��+W���H��Q�x�a]h.�/%�{��   ���;  p>%�w����w�2�log�����v��Y������_��dԟ����3)�w� �eWK�r��'�fRv��y�R|��L}uu2~m-���IA~u5���ɺ����j*���%g����MI>��J  .�  ���I�$��p
��Evt�zs3�[�f��;;�u���������NV?m�$˙�[��X,�L�����4�n&���%CqjF9x�����_m4�8�_�t�,����_��Z�u��N����<��tT3��'��$�^8  p�(�  ���I~[��:�w�Ӹ�Os3�â��p��tݰ��p����wwKG�p�\A։ۣ 01��i9�I�Iv2������ٿq#�7n���F�%�z�����������h��j��땎��]O�/���${��   ���;  p��!ɗ��ks{g�Q�����3���`k+�۷3��N�����������GS�dR{'��; �O-���� ���$�qԨ��hs3����ܷ�h������z�kki��M�76R��Hcc#���4�^Mui���lmmM�����I�E��,�  �$� ����I�f�<܁�����������͌��ܺ�a��a�wg��V�#u��2���N�:| �y��Ȥ�ދQ�<�Q���͛�߼����=~6���<\6xTkkky�J�ൽ-�H�-��   �O�  8�����o��0��3py����LW���`{;��������o�����x8,y��2�Ծr� �����N�A&SݻI���=�d�j�1��ʝ絵4�^�L��r%�É���Qkkk�#��)�/$���A  ���|  <�f�Hr�t���0߆������ܺ���f�_z)���72�vK��-eRj7���TO��d-�n&EwS�9o�~?�/����_~�}��l�ѩ�Ǟ�\I��T',ǲ�J=�w%��I��  ��>  ����$�^:�IA����q���߼��[�ҿys�����+�L�o�ʨ�/��TM�Τ��(���R��wP;���;���G%C�	�n�n��{�U���������k��{���I	���4�^M��`�9�5w^��@�?7�  ��;  �8�l���t���j��pƃA��ln��p����w����R^y%��Y3�R{;��P^=�F�Lu�N�2:��`k+����~���ݧ�h���ө��+W�|��;��]K�Z=����Pp�K����&�K��   �I�  xToN�J��᭯��� �ʸ�OssVV�>�߸1�Ⱦ����_NFf�.�j�V&��f�, p�j���� �����1����F�o�x�������a!~�p]���TM��"k�[!�L�]��   �G�  xk��f�S:��+xp�^/��7'�[���f7o��֭��J�ne�햎�T���j&�A ����z&E��$��������y�U��w:�_���իi\���k����ki\���k�./�SbX�5̭J����M򋅳   sF�  xX�$�N�J�јz�nw2q��i��	�/��A�W:&s��ɴ�v&�0`U3�Hk%�n&E�����bt�t������O�ј�ߟxb6���w&�_�����9���gX�\�$��$�'���   ��;  �>����Spg��ܼ���/g�p���+����sp�f�ne40���Qɤо�I� .���v&��${I�%C�7����F�o�8y�J%���;S߯^M����T�k�Ҹz5�����rI�r,k�}j��H�奃   �C�  x(�ה��qR�y7���OZ�q#�/�d�:箖�(���e �̖�LƯv��&�95��$���]��zj++�I����+W����.âX]]M�Z�h4*�G�eI��$�R:  0� ��d�w&i���YYY)�k<ep�V�_~9��i���7s��+��J^y%��;ZSV#�R{'�ɶ �H�I֓�%�e2ս_4\>�� ��|�gNܧ�j�y�z��x"���'S�_����_�����9���S�T�j��u<`��I~.�ϗ  \|
�  ���&��$o(��g�;%��ɤ������b^z)/����l\P�$��L��EW��b�N��L���E�b��f��g���'n�6w&�?�T�old��'���i^��T\���X]]Up��$ߛ�w&�U8  p�)�  ��|v���9K�~?����߸��728�:8-���r��Μie2��Y: \P���A��$�Pިߟ��l���g{�^O���c���a�}��'Ӹv-�j�@r8���j^x��1x|��I����g  .0w  �|Q���tNG�ZM��)�96�2x��%�χ���ۥ#©�$igRlw  L3��L~�>4��b��I*�ZW��y�z��xb�|X�o^��ƕ+眘E玄���'��$o/  ����  ^͛�|{#�.�N���[����~�ľ��s��g����d5I�p �W�$��>��d��{��|���_z);����l�N�o>�D��zjR�����SO��nH�e掄��7$��$��p  ��Rp  �{�\/��c�S�^/�/����<{�?��>��)�]-w�����Qˤ辖;E�a�D�i9:~���g{�әL{�����i���<Ǵ.�z�w&�]I^,�  ��9   ��[�|V��.Ӯ�x<)<���������ǳ��g��U:\�LJ�$�o g��d=��{7����h"����y&�g��g[�ZMcccRz��4�z*KO=��'�L�u�K��*����1�K�u�X�ܸ�  pw  �$_��ϗ��s2�r�����ǲ���MJ��?���</���@uN�Ȥd�. H%�J&���lE��x4��͛9�y3;��+�l���f���f���%��)���K�s���$_[:  p�(�  w��$ߞɐ=.'�_�֭���},�g��,?��";< �v (��IɽEw�^����lo'O?}϶j���Of��o����/=�dׯ�Rq_���1�K�'��$��t  ��Pp  ��&��$WJ�l88?��������{���~�����_Ϡ�-�R#�j&e: �b�ݏNt�M\t�~?{�=��瞻g[�ٜL|?�������
��������֥VK�Iޜ���Y  �B�  8��$���!8;+++�#p���t?��t���}����y&��z<.�v �����0�F�}���>��=۪�z�O<1)�?�T�^��,=�T�_�z��9�֥�d&�W>7ɸp  �Pp  ��0�_*��e���q��K���f�C�ί�j�>��d����F��L�r ��Pt��h0����g�����V��Ҽv-�'���ߘ�7�i2����1����$_���s   ��;  �$�O�I���p��<?�~?�8��>���O���2:8�pw7/��A�W:"\J�� p9(��e<f�ƍ�߸��~�ضz�=�����O��o|cZozSO<������t:�V��F��p��!�O'���9  ��� �J����6�\rn�|�F{{���Cn��ϥ�k��Q_�K#�z�V�  ���ݻ��e� f��e𑏤���[_m6��������4L|?3�J%+++���*��UO�]Iޜd�p  � w  ��|^����Fs37~����O�d������B����v5 ��:�3��v�a�8�����3�=�̱����,��i��MY:Z|�v�P��E�}a|B&Y��t  �w  Xl���o���1��t�����������/����q`�Ԓ�&Y�b; ,�J��w2��>*����^z�HzwM|��Z�I��G�W�J:�nX(,�_H�J  �Pp ��u5ɻ�4J�|T��t:��1.��G>�_��o���ϗ���I�}�p X<�L�t�lgRvWt.���nv�~:;O?}l}���շ�%o�3�P����p��$?���)  8� ����$o,����tR��s|n������߮�稚d-�듬�A- `�}`=���.�|t����_(cn(�/��$ߝ��[  �c�;  ,����J��|9	x
��<��w�Ə�X�$�0*�Lg]KR+� ��jI�d�}a+I7ɸh"����K��l��r�9���~s���*  8_�] ����I�^:�oee�t��6��w�C��Q;���W�� ��i���$˅� <��h���+c.8����*�Y:  p�Lp ���L�L��`�|t�?��|�]���/��a)���3 ��j$y"�^��$��q ^��sϥ�ɟ\:ƅ���B��$�O�L�   ��Pp �������t�p�7���3������_.B=�Z\� ���L��Mr;ɰl������r�t�9���B[K��I>+~� �B��   ��?��-�r�|8��<�_���Sn�sP��L��� ��N��'وc�Ŵ�쳥#���g$���!  ���8  ,��I�Y�`�9	����>O�7�����Q�R�$Yɤp�~� �,T��frA�J|� .���+a.�@��I�9�C   gO�  û39��s��wv�o��z��Q�R[N�T�+q�
 8?�L�<��������͌vwKǸ��"�_�ߙ�u�  �%��!  \~5��AyN>�����ٿq�t����ʞH�(� X\�L��\��$�0g�c+���k�Z���cP�'$yG�  ��Rp ���w'�[�Cp1�����p��~��y���/.���R�
g �j�]e��a��JG��*�J:�N�\_��K�   Ύcu  py-%yW�u�C&�����ތG��1���$y]��$��Y  �V��{��2��P	���-���$��t  �l(� ���-I>�t.�_�pw7�?���1�RYʤ(v5B _-��-O�g����@�9b%�wg�+  �d�[��g�΃$�����'�y��*+��2�>zfZ3�:G:-����&8���#K^H\���]�»f9�?�`�]9 ��� )4BB��cFs�Y��u��GfUWOWwWwg���|ޯ����|���ROW���<� `8}�����p]�-��b�ӟV�Z����rXQ�g�  �^�j�3.s ��	��C�/򤤟�   ��(�   �g\��qJ:���8�1Bm��_�� <G҈�S۹�  ���?׌��s �RmwW��=����8�?��F�    ���   0|�����[���3�XG ZBҤ��8�  �����7EI�q ï|�u������JJY   �=�7   ���$�w�!>L���V���ښu` �%MH*H�   �v�}\R�8��ut��u���n�I��:   ���   �I��u��wVY[�Z-��@q$�H���4�  �/i��a~0�^�0������;�!1�   q�     ����F�� �X����Ɔu`����:� p,�L��n���d�8�$ɉ�K�O^s�@���|�۞�⸮�.�s|_n�|O����>?9�LJ���%7���=V�ۻ��t��=��rLc���N�VS�\�$5�u5�/4����wj�x,�^*���8~��/5�w�+WRNRJҶ��m C�	�w�9.܁#�_I�I��   w   `8�G�߰��b����J\ n�U�J��ګ� ��tQ<���K����r;E��8��DB����}�	�q���r�qqۉ����S_�X������hk�U���<n��jV���f�r�q�z�h_��qt���N��V*I����j6jH���j��j�|�f���ڧ��_RQҁ�]I\��A�)���pE��|�u    ��;   0�^!�}�!n�SSPq����R ��R{R��g&�K��z^�>�A�X�+�J�L6������TJ�����N��ssy=����@��R����l�0I�`�)ͷ�uՏ�����4�ە���'���}��@�rY�rY��=����#)#)��4��m �����Ύ�\�:Jhq���~Hҿ�   ��Qp   ���D��:�VwV/��# ��4�viT�﷋��t�P�%�����y&Ӟ|����=�}|�T�fO��N1=��7��0 Lbɤ�L��h�j6���o��e5U��o?>U�ot
�����㣣%�r��9GG�׸�r��%�.�oK���0��׮Qp��q�>$��%=o   ����   �_��r�?��l�_�� ���4���c��b�����X:���ȍ�y2��Ȉ��t�q���dڟ�J���dK����{ @w9��x6��"�M��K��Ǎ���t�NI�V*����W�s�88P}�}�L�G�%$MJ*Iڗ�� �U���<�u��J$�<O�Z�:
�-#�$�E|;   w   `p�N�OY��``��۫�J:|�aN�i��S�=� 8��*�ɴ���l������d�v���L�]<�|K���u���� @��i�����������|�vR���;y��������;�����Zu��WRNRJҖ$*� �Eyy�:B荌�hkk�:��Mj�?��u    ���;   0��'��=Ĺ0���v?�9��M�@(���j�9cj{4�TP?u;�s�i� �p8���/��k4+��S��OO�otn��]���T��U�s߬T��'<�����%�� Χ��b!�2�w��/I����b   ����   �_���Lp����>g�@Ҹ8Y4b���\�d��I��%u
� ��� �R>_�߬VU?�����z~X.Bu$�HJHږ��?���~wr�=HJ�CI���0�   ��f	   �7I���!08\�U���Zͦ������:��N= |�x\��⣣'�Ǐ�\��s�l���y�zl� ���
��{����ލ�{��Z����[�TR��GG=��<8ORAҁ��܇������j��r	�(�E���5��#���    8?
�   �`II�=�<�A:���8�1B���gC[��������~{���T�ν_(ȟ����*62"��1^>/�u�� `�xw�`f�?�^*���q�����Ɔ*���"����}u}]����	n�H���4�r_���i�TY]Urq�:IhQp�}�YI�����   �|X�   ˇ%=b��E����җ�# &\I9I��p�XL��X�6>.|��8�k��s�vI���u'�� @d_Tv^��#�wwU��Vu{��xg�侶�ݾ�����Z����Ӎi�;b�;�[���)���p|I �U�j�Y    �w   `p�7�~�:O&���Z{�A	���S������(����������r
&&?.���+>:j  tQ,�T,�T05u�ϩ�﫶�uS齶���Ύ��B|}gG��Mն���9*���:Ls�b��e��ƹ.ܧ'$�_�{��    �;
�   �`��o�����֪�t��3�1���IUt����2�՟��?1�x6��P�?1��Ȉ�lV~��`rRN��d  ��♌♌��<�Y������ޞ�����V*������ummmimu�=A�TR��\w �*++�B�s]x ?-�O$}�:   �;c�   �4g��m�϶����YcGbDCRҘ�1���Mߤ������(   '\ߗ_( qF    IDAT�/�z�3��V�Z^^����j���Ƿ�ݓǵӏwvT����`Qp�3�u��%����K�(   b�  ���FI�o��E��~�k���s՞���v���~��)� ��������]W���>�Y.��ݏK���v1~{�=5~kK�R�2<0 ����B�s]x@�Iz���X   p{�  �p�H����(��m��v@�C.�4�h����S?%/���  �@��ǕN�u��u����&
��LM������j;;����ꥒ�����v������Gp�GG����B�����.�'��/I��   �lQZ�   �oJZ���Ƣ��(�cX9�F$e;��b�e/S�[��:  @WA���%mllhssS�V�+_7�N+�N+1;{��Z�Z������ޞj�%���wvT��QugG�RI�z�+� ܬ��L��68ׅ.�$���WHb{    �(�   ��vI��u>�nU]_W�T��t����v�:�����.ɉR�  ;�qT(��dt��uU������������w=������n������������R�Ύ�������h�!90<����c�Y�%���*��u��%�O��Z   p+
�   @8%$��$�:_&���:�<c躌���5��X�u�S����  ��dR.\���vvv���">2��Ȉssw<�qp�Zg�{}{�=��~}�dJ|���Sr �*kk�Bmdd��;��g$�����   �f�  �p�����C`80��V�>k蚸�S�� �~臬#   ��뺚����Ȉ���U�׭#ݳX:�X:����m�i�j'%�Zg
|mkK��]U77U��7�8��R^Y��j###��ذ����K�=I���V#   @�Pp   ��m���u&����k_�� tEJҘ���G��4��W[�   �L&�.hyyY����q���<����B��5������4��榪[[�u׶�T��}-U
�w�@t��%�O�~�:   �(�   ᒐ���vW]亮��u�Pi�j:�|�:�@\���)� !0��wZG   �x<���y���jeeE�f�:R�ŒI�fg�7~{[��U��T=~���~~wWj���8���Z���XG	%:���+�����     �(�   �����J��z��^P�^���7�u5��+5=���v��T�޶�e"�J��-�b  ���訒ɤ�^��J�b't�3�U��L�om�ڹն�T��Tu{[���>�nh�˪����嬣�wt�/����:Iѻr   !
�   @x<)�ǬC`���w��g��� ܞ���?>.o|\~>//��76&?����k��G��o����7~�a`[�o~�b)�� ���}_KKKZ__��֖u���x���)SS�=������*��nn����~~cC�j���%��
��9/��k$���>h    w    ,\I��Y�pI���B��k_�����ӊ�r�r9���r9�s9Ţ�\N�Ą� ���b��fffnY�///���ۯ����ۭ#   �s]W���J�RZ^^V�Ѱ�4T�S�o�����Ύ*kk��������Ύ���nl��d 0�]umMz�1����bg���K�cI/��    @�   ��Jz�u
�:|�y�R�TJ��q���	��S��ޯcJ�Ӛ��Q<~�i�����F�������&�   �122�D"��ׯ����:N���i��i%fg5����~2~kK��MU66T�ظ1	~cC�Z� 9®��j!����IK�7���   0F�   �����X��pb��f�rY��u�@���/䏏��?1!?��76�.���r�����8���*
�=��_��{��K_��   n�y��������8�8��z��.������~r_��Pu}�|D�WV�#���Co��j�   ��   ���$z�	�nV�rEj��c �\�k���

�Ţ�\��.��[��433s�-����>%
��+^a   ��Q�PP:�ֵk�T�׭#��٬�٬�.��z��@յ�v�}mM��m�vv�e���ըT���Pe��m�k!z�7$�GI\e   ��   ��Q��)z�����\�� #�+����{Xd�YMOO�uݻ�	��  �(�J顇ҵk�tpp`(�N+y�¹��uUVWOJ��j�ω�������}��zPp�=6&�%��    @TQp   �LI�%�nw��5e
�C+�N����-vrR��o�x�f>�?�����v�!�R/ZG   �X,���mnnj}}]-v�Z�[��������V����8�F��Z�$ot�:J�PpG�m��l   �"
�   ���MҸu7�nvt��u�'otTA� obB~>/ob�]^��;�o�x�����{�(���g{�(�\�Wbr�:  �����J&��v����u�S��h�������j������I����ݞ"��
�gH��r]WM.�@o}XҟI*Y   ���;   `��Hz�u�t:m!Tʗ/[G�m��מ�^,�/�����bQ��YG�t:���Y�b�{���K�z�(�33��Z�   (�TJ.\еk�txxh!��b�����j5U77O
��UU�������(���8Z*���<��u��qG�dR�Q0ܦ%����   Dw   ��2�>d�@����֖�8Lycc���z�s�
�r9�x&������}}�ѕ+]N3833�   R<����׵��i��<SS
���|�V*��)����T��kk����9�𩮮ZG�t:M����%�����:   %�  ���uIs�!�L�:Bh1���\߿i�_,*��8yn���߫X,�����%��c��  p��Q�XT2������u$8/����*}��-�5+����WN�߫j5��Kye�:Bhe2���Y���s%����I�g   "��;   �_OJ�!��
�7Dy�u7ųY��JLM�/N��^�(ot�:�@H&�����������V�7���   0�FFF��^��J�bC�%�畜���V�����M��ӏ�����;���%����X   ���;   �?Ǔ^�9}�8�M�6����f�wJ��Ԕ�bQ��I�SS�%���Z.���Ԕ�y�U��6�T�:  �P�}_KKKZ]]��ΎuD������5r��������U�~����'��1*�o��;�콒����Y   ��b   �?�T�+�C :��\׵��o�e�
:�`r��LMɥ��u�XLSSS�f�]�����m  ��u5==�d2���U5�M�H�$��7:��ŋ
ff"[po�˪��k��>K�=����A   �(��   �Ǽ�n���Z��*���1L���Mʾ�U���$%�>�}_sss
���_7�����u  �����H$t��U�j5�8�M��I���������/x�����9   ��Ǹ+   �?~G:s�e�g�buCyyY�F�:���7��^�z%��(��Q:�օ�^n��V�'kRp  �D"�.��$B'�N+ῗ��U���J��# �>$i�:   0�(�   ��NI�:��B��+W�#�r\W�������5??/����X"ѓ�;�  z&�i~~^�|�:
p?�S�+++�Bid�y"01!��!   �aG�   譌�߲�hb���ׯ[G0�OL���q��u]��̨X,�q������=��a�w  ��rG�bQ���=�`�WA��Lp?�`��Iz�u   `�qF
   �!i�:��E���t��㟡~�}_KKK��{E�����u  �H�f�ZXXP<��D�����ù/r%�+I|�   z��;   �;����C ���~Cey�:��$��H�RZZZRЧ�y,���ʊZ��u  �HH&��p႒ɤuD\P,ZG0���q����3�!   �aE�   ��\`�)Vm�V+��Lp�\.����b���g�'��&  �Q<���r��uDX05e�L�\V�T��:��4o   F�  ���QI���hc������f�j�Tbv�:��rG333�����8}}�(�%����   ��8����M~�$)����`*��%�N����%�/�!   �aD�   �1I�0��-�S��Ubz�:�P:�b9::j��n*e�aqt��u  �H�ؽ��x6�X"a�L��o��u]%�I��wH�N�   ����   t�oH*X� (��U���#�
���x�u������L҃�	���2w   3�TJKKK
"����/�#�a�����!�[���   tw   �������! ��c�O8K��ZG:�tZKKK�/��y���V�r�:  @������%.�F_SS��Pp?���~�:   0L(�   ��H�]I�эP�d��-�ss��J.�����\����7>n����O[G   �<�u5??���1�(����u3����/��OKz�:   0,�Wc  ���^i8�����uSLp��q455���i9�cG��OLXG0UYYQ�T��  y�?+OF�x��	"�����f!�8��	$}�:   0,(�   �Q��s�!�c����<��Z������1L%ff�#�X,�����M��y�����U�   �����b16�C��Ţu3��5�c�w���%}�u   `Pp   ��7%����Hcq����*5��1�8���ۻ��}---��)����~�:   N�d2ZXXP<���!LMYG0��[��i���}HR�:   0�(�   ��u�0�q-����#�������u���J����$?�����1�   |��.\��D"aC�����w�~���[G
��YI�   :
�   ��q$}X�l��aq����b�T0=ma`���jaaA�X�:�m�A���uSLp  �x<���E���XG��q�Ţu
3Lp�CR�H�c�!   �AF	   x0?&�5�!�cq������W>���̌Ǳ�rWɹ9���^�j�:   �ຮ����筣`�$&'�#��Pp�CR��i   d�  �����s�!�����v��l�T�	���qMMM�8@� ����L�����1   p�bQ�.$����}���[G�< ľY�wZ�    w   ���I��Y(��U">�����O���rO/�KR�_��   �����\��I<8�.J�*�oA�!�[��   � �,   p�����C �C�]j���g�T05ea �b1����x�'�K���h   ��f5??�X,f.ʿ�V66�j6�c�
��r��~�:   0�(�   ����[� ng�����f�����c����ZZZR*���r_�ss���~�s�   pN�TJ����<�:
X"��[��j���1B��;��%q   �G�  �{����j��d2i�\u}�:���ԔǱ�j�dRKKK����^)���֖�ׯ[�   �9A���%%	�(P�Ą�x�:��J��w�X,S�1�;IK��u   `�Pp   �MZүZ� ��UR%�܃�i���N�����X,f���㊳c�J_��u   ܃x<���E~w��q���u
3Q߱�,�[��%}�u   `�Pp   ���K���M��k�'�SS�B+��i~~^�;�E���Qp  <��j~~^�l�:
P09i�L�w�;w G҇%��   ���c%   菇$��u�<�ɤus��/�&��~���	MOO�q�(]�~����(�  $�q4;;�|>o&����Xw
�OH�1�   ����   �߇$%�C ��������399��nc������V}o�:   �S�XT�X����G��^������R)��y����u   `Pp   ��풾�:p^Q_�k�Z�nnZ�0�OMYG�q4==���q�(=�wIͦJ���u
   <�|>�)~��9%"\p���g�d2������   � ��   ܝ#郝{ ���b��uS��5k5�f�lV�d�:F(8����Y�r�;+}�u�P���g�#   ����ivvV��)ܙ����}5���c�J�=`����ǬC    aG�   ����j��y��'UVW�#�
"<��4�u5??����(=卍���c���  0�٬����,c����	9�;R]_��*�t�:p/<I�   �]t�   �'-�}�!�{���,�Fy�ݱX,�����,r3�]���W�88��  �.�d2������d�='W|�w꺛�_��bQ��C�[$�M�   @�Qp   ������C ��	�R%���Op���Z\\T2����7ܥV����?o   ]�J�����x<n!
��T�֬#�
��0�>$�or   �mPp   noQ�?��+�X�MDx����Z\\T�Q�*��#�Ba�3���   �.
�@����}�:
B(���Q���Ř��uQҏY�    �;   p{�%):�142��usՈ/��]�r�%����Ba��;  �Љ�E��;/��#~���(�c�����u    �(�   g{��wX� �ܥJ�'�SS��.�JiiiI�x4wvN.-)Ƃ����%����c   �����H$�� D��	�f(�ߌ�;ظ�_�   �Q4W}  �;s$�f�8Q/��j5�vw�c��%����X��t:���9�nt��w\W�G��g?k�V����|F����:	�ЬV�,��8<T��P�VS��H��(�ժ�ڏ���j6�j6U�ߗ$��U5+IR��P�z�}l��V�����-��8u왙�e5;�{�׫�[���Rr���X2y��n<.�E?���i����ǎ���L5�%�r=O���M$��b'@�29��~�sL,��G��@�� @�b1-..����:�|_@��Q�ྱ!�Z���K��;�K������    aB�   ��Hz�u�~e:������y#*(�#���F�x��������X�ZU��@��C�K%5��ԬT�88h�v\N��T��W�V;)�7�u�K%�����u������s�<H���ˉ�o��;���i�(�����(�H�M$�d�&��ǩ�b�̍�FF��DB��_�	�������]�zU|ψ����{Z�VSmgG�ؘu�P���<_�Ŏ�   �M(�   7$��u�AD}Q/��t������r��F�x�:B(�|�S��Ъ�����q9��@�����>nt�;>��y���;M:�ph��j�˒��ϭ0�T�]v��>�&�%�e2�w^s��vi��Z|dD�tZ�ų���##r=�G)��뺚����������jF�g����������g����6I��   �w   �f�TҢu�AD��^Y[��`*��{&����,��S2/}�u�P8�tI��U�o�ӬTT/���RI�RI�����O�~r���t�J�s1E7
���+����ApR�?���Y�FFn�?~��g�4��!I�����U^]��b�����ŋ�1B#�NSpǠ�MI��ݭ)  �S8k   ܐ����!���d�#����B�:B�e2����q�(�����76����us۟��������f����j;;�mo��;���wvn*�����c�ԬVU�ظ�Ϗg27M����3�s9�cc�����˝�;\h�r]W���v���Y~�݂{���X*��6�c��J��H�#�    @Pp   n�%I��!��	�/�OMYG�l6�����y�K���[�0���S��_��-%�����Ǐwwo<��8:�N��������=����Tx����W��7:z��W,��Az �����,%���E޷S{����Q���"�%U��    �(�   m%��u�"_p�ܴ�`*Q,ZG���QMOOSn����^F�]��SOI����<�V������[[�nl����������������mȋF    IDATm���-5�֑���-����7⽱1���������	y������
�%�=L������U*���ςܙ�~���h��1/�]�~�:   `��;   ���|�@7D}A/�w��������'��WXG��֖��yF����:
B����.�������.�oo����PukK��U����2�z����9'�ƒɓһ��˛������

����z^����8��NO����q�G^��Lp�Y�>`��G��J��IN   @�   I����:���ɋp��U���m��Ba(�\N����1���}��x\�z�:���O~��{��vvT��T�S\������yRd?��Y�YG�si���]�r�c㣣���v�PhO������+>6��Xl���bH@j�܏o��Q��^��T���� �#�N[G �%+���~�:   `��;    }P+A
Q�VU�ܔZ-�f��I�]w<��K&�y�Q����j����?�����f���ꪪ�몬���'���4�f�j ��wwU����s���8���ML((������bQ~�(b���XǓ�%J�Q�G��ެ�T�ّ76f%(�c����ߒ��u   �
w   D��Hz�:�-Q_̫F|{�X���U���'��_�����.��/����x&cwЬVU]_o�66T�vM�S����mm��lZG��ЬVU�~]����x\<�mO�?�
J��ʟ�PP(�<�����Z��J��u�X|dD�DB�r�:�������}���$����e   �B�   Q���!�n�|�}s�:�)�
��l����)��W����us�z];O=��o��(�լ�T]]UyeE����_WumM��$������  �ꥒ��'�ǒISS�{��`jJ��)�[bfFn�15p��I�܇�_(����&���J_�h#�~NC���,�/��    (�   �~\�#�!�n�����֖uS�2EsddD333r�:�@}ի$ǑZ-�(�?�I
�=ԬTN&�]�z2q�������u Z��#>�����ǜ����Sbv�d�_((����}L�(9.��Z-���Y�AQ.�G|'��(�c9�~]���    (�   �R���u�ۢ��W����	�lddD��������)����^��bn����0�껻:�vM�k�T�~�=��3��������uD @ȝ����S����337��OM)��>�8(��Y���sG����z�������G��b��Q]_��Q?'������]��c   �7�
   ��-i�:�mQ_̋��`����4��.ɾ��%UVWu��J=��u�PjV�����:�zU���U>��N	 �c�J��S�]WA���쬒�����̍I��|c 9����9J�C,��
�Q?'���k�>*�-�   )�  EyI��:��T�:��(Op�g2r	��-�Nknn�r{�����Z����:F(l}��.��K%�;S؏oGW��//KM�� !�l�����ʊv?�[^v}_~��.��͝���J.,(F��'���Љr����O��91��%}���3�   �w   D��%�Z� z!�ӪZ-U���S����r���Q���OZG��O|Bs��}�1z�qp�.�w��/��ެV�# �3�j��������u|������Y��J-,�/Ò뺚��ӕ+Wtxxh]4ȿ?���Z��K�d2��^���'�b   �
�   ��I�:�+Q.��J%5k5�fuA?�JQnXTrqQG�.YG1W����8<TlP���Z������e]�rRb?.��ww� Zխ��E�_��-��A�����J��+ٹ%��P~Z��j~~^�/_��ёutI0��wC�^W}gG�ؘus����<�"|nCmN�?��A�    @�Pp  @�����u�W�ɤu3Qߖ{��ɤ���)��H��.�Y�i���J�o}�u�;��J'h�{N�=�.�_��F �f���g���3������%fg�z�!�zHɹ��4��i9��:�\���.]��r�l]�&�g2���[G1Q]_��ޑJ���E�^��I%�    @?Pp  @�|����:�KQގ���e����[G�'APn��k_��?�c����񏇢�^��R��^���ի:�|YG�/�|�*%v  B�Y��\x���S7�K&oL|_\TjiIɥ%����Z��tɽR�X�A��b��闼�:F(��i
�f����w[   ���;   ���$ŬC ���p���	�Ţu�s�}_���'��rO>)�u�j6�����˿��{���~|;x�Y>�ld7  ��ё�~ZO?}�k�lV��~�a%fgO&�'����B�XL���t�j��u< bB��=g�De}�:BhD��"��%���U�    @�Qp  @T�I�7[� z-�LZG0S��wb�:¹��q���+�D��GG�~��Q������^��������.]��K::�]���+WT/�S8  QU/�T���U���oz������pAɅ�.\�Fi!I��Lr����q� ��n�Rp?A����~I?b   �5V�  �"ɱ�Z&���`&�����Ŵ�� ����D��ORp����'��^/�t��s:xi��=��^���  ΩY��v�?1��C���=����*዗��x��K�.��hX��}��f����B��;"��ޭ�Y�    @/Qp  @|���X� z�u]%	�f����fC?��u]���)y�a�{�ku���[�����k�{�����)�.���N���I @�T76T����SO�x�u���U�ᇕ�p����r�X�'� ����._��&2� �w&��H�R��~�$����   �w   D�/Z �!�L�q��QA��a_�wGsss,4}�k�z����us���k�|�S:�z�]f�����++jQb  a�l���]��͏}����ܜ�/�o�<��ŋJ��H�]�[�ɤ���t���Z-�8�G����j���H���~Yҗ��    �B�   �^g�(��[���{{�1̄y!�q��̰�l$�Ji��/��g>c�\�Z��ǭc   ܿfSG�/���em����<K��\\T��e\�V��Eycc�aS:���̌�]�f�����n$/^m5�mo���b.���9�ڃ}�i   �
�   f�����K���ie�OLXG����)e�Y��6��7Pp  b��C�������я�<���Q��G�y�1�{L�����&�lV�FC+++�Qp�S<�Smk�:����&w1���^-��A   �^��  �a�}�^n�H�77�#�
�E�g���T.���ycox�^��߶�  �>+_�������O���9�PP�Sv�<��2�?��',�����hh}}�:
�AP(D�ྱ��ŋ�1�%�I�@?��~E�7[   z��;   �U\���C ��E�Z��a�����5���Pȼ�%�'&�;    Ҫ���Z_��_���s�Ą2�?���W���T��/��H����	5mE�0=���	�_��a"��E�Ey�"뿕�fIi   �6
�   V?,�a�@?Ey�J�a+��������p�^�:�}���I   BՍm��_��ޝx\#O<��7�Qcox�ҏ=&�u�Sژ��T�����u�C09i�L�w�;F��+��b   �6
�   F���X� �-���Q.�;N�
��tZ����1�"c_���  p.�z]��^��^/������{��5��7j��oV|t�:b_MOO�^�����:
�"L���6
7�=��Ϭ�    �D�   ��'$�[� �-ʋx�ܽ\N��Yǐ$%	����q�(x����z9��V�i   �����?�S�����<���*~۷i�-o�����z�q����^P�R���;��f(��E��"�E�   C&��	  `�����u�B������!�P�y����亜j#o|\����  �׬մ�������w�S��-z��Veu�:VϹ����y!��g�E�fj�B!ʻ"�^#�ۭC    �Ī3   ��OJ��X��"^�'������({��[�j   C�^*�����>��w�+�}����%�H=��5??�X,f�ፍɍGs���GG�1���q��Y��_�Ķ�   �  0LI�XI���L4+��c����jnn��0���XG   �j5Z��?��~�����i>��u��	�@sssr����8�#[�2�]R�w8D�}��wX�    ���;   ��?��aQ��^�޶�`�z����4��"}񢂩)�   V��6?�1}���[_}��T�~�:QO�R)��p�)���	�fj���B�s���)�   �  0,��@dEu����p�~rrR�l���q�G�o~�u
   �V����~T�]ߥ����ժu���f�*��1p� ��#~~�XTϏ_'�oY�    ���;   ��O��툸�.�ՙ�n��|^���&����[�#    "���.}�#��w�v>�)�8]��D��	�[[�B!��ǀS�/��  `Pp  �0HJz�u�ZT�/������Q���'�T,���  �9�|Y_����������q�jrrR###�1p��E�aP�ذ�
Q=?��2I�   <��u    ��%i�:`-��j�'��	�2���g"����T_�����r��6?�1�(x@�Ȉ⩔�x�����J��x\����f���ё$�~t�f�&I���~x�f�n�  DR��������O��_�Ee_�r�D]333�˗/��sl�Q.�onZG
�$�$����u   �~Qp  ��KI�I��5���y�u���=���<����u�n����V
�!�}�gg���VffF��I����y�cw}��Ͻ��j-�$�j��mc��`�mC�6�� `[� �2�0�$3����0���p29�$�2L�	�<,�L���q ����^��k_�>Twu�{�E�W���:G�dI%}�������/Q((����W��)��)��/�	+KKZ������ssZ����쬖''�t옖��ұcZ��k  @Z=vL��ַj��߬]oyKS��X�}_��㚘�P��	��XG0S��.�����,�U�>g   �.
�   �v����荒��̴s2],Ӯ]�J�v�;���j���Q��yʌ�������u�^s�F�=��2N�N+L��7>~��U���x�����¡C�}�1�>���T�\nSZ  �+��}�SZx�a��)h�T�����u��!�y�m**���S��V�^�Gv�	���#�/�w   t)V�  ����c�./ޭMMYG0�΂�����x�^�
��t�~�:J��b1�o�AśoV��땻�:�_w��.���R�_���_���Z�\���G5��i��I��E��  ��L�z�o�͟����w[�ٱD"���Q9r�:�Ӽ0T�ͪ�����z]ՙ�����i\<�Mb�;   �w   t�wI�tW�jU5���a�Ж�R��*��]wQpo� ���Ӟ�ҭ��p�*=�z���)�o�r��i�K^�q��ѣ:����C��Ci��A���8  p��Ç�Лޤ�~�w�{ֳ���X__�599i�iQ��d�]�ʧO;_pO����N�a1�   ]��;   �U$��!�N��t��쬓ێ�Վ	����*��H����u�&���ct�Xi��4���n�]�k����ֱ�e�Ɣ�5/{�$iejJ�����}�:��ojuz�8!  �$չ9=��w�)��J��ggǊŢ*��fff��8+���[�0Q>}Z�׻]=F\�͒���    �VQp  @��eIc�!�N��t���%�p`��ϟN�5<<��׀��S����V����u2cc~�s5|��ٿ_��;hlEr`@{^�)�s��7�����&��=իU�  �Z�\��տRuqQ#�|�u�R�\��Ғu'��d�NU����`��cd�|X�  Ѕ(�  ���g�$�N�*;^p�Z8Y=�k||\���5`�p�:���Y��
��>U��W�^�b���e�����Sn�>����Z�����{��Wt���V�\��  �4z��[^j�������yӡC����f�9Q�O�d�ӧ�#�s�pϔ�����    �VPp  @7z����!�N�rt�p��-�=�e�X,���q��ߒ�Gg(��Eܯ �o�v�s���w��{�X��Y�lV{_�R�}�KU^\�ѯ]���ou�[�R�R��  ڬQ��я~T�rY#�z�u�9��jbbB�Z�:�S\.�W(�3�����;   �w   t_���C ����T�'��٬�0l��z����qEQ���Fg��v��\Nչ9�(#=<�}�߯=/y��{�Z�qN��蚗�L׼�eZ��ב�~U��E�z�!�h  ��=�;�#?��+^a�fG�(����>�F�a�a�h���=F\��$�H��k   �,
�   �6o�t�u�Ӹ:���p��U醆���yr����?��_��uS��k����u<���H~,f	Z��~�����������:��/�����U�� ��F��G�R��[�ّT*���A�<y�:�3"��SS��%	���z�n�4�F�  �E�k   �ē�/�C ���Bruf�:��VL���r���M^t���w[G0��M>����E���_�﹇r{���ޭ[��n�����;?�q�~��yֱ  @�5�U=�h��ǭ��X�PP�ug��i���][YQme�:�)���\��\   ���w   t�_�t�u��Zpwy��x�'�'�I���4�9���o�]A6����u��z�st�/��F��GI����P��G��G����:����jkk��  @�Ԗ����ާg�ɟ(��q�����������
�=j�DyjJ�]��c�J�RZZZ��t��[ҽ�!   ��`�;   ���e �T.���*ss�1̄�BӞ+���S�u�*�u�u���|_c/x�^������4z���w���ݺ��]?��/��w�[�R�:  h��c���>�z�leG|��������c�5���nRqx�YLp.�nI϶   lw   t�WHz�u�S�Xp��ΪQ�Y�0�MyJ(�}�u��	3������/}I/��AO{�u$4Y��_7=�����t��>��޽֑  @�?��&�����c�\�>Q�>3w���)��\<Nl���)�   @ǣ�  �n�A� @'sq�:;k�T�I��CCCL6s\��X:m���Tj����/��y��CC֑�b�(�u<�������Wv��H  �Ɏ�ٟi�ߴ��c�dR###�1z��ܫ���̹x�؂���T�   ��Pp  @7x����!�N�bA����m3&�
���7!��E*�y�u��	������^���݊g�֑�f��k�=���������շ{�u$  �,�����Tun�:Ɏ�r9��y�=��{��i��(�W�K��   ��Pp  @7��Z�:�e��p�r��}};z�T*����&%B�+�}�u���P�=��^������_�B�:�m�?�Y=�#Qfl�:  h���I=���Y�h���!�{l'�N�t����%g�x�آ_���   �h�  ��n�t�u����q��{荒��̄���m���05>>.oρޒ߿_�n�	����/�+>�y���)�p�����y�����}N���*�D @כ�����/}�:Ǝy����Q�ah�'EM���[U(�Sp�.��A�   ���׀   @���x�
\���*�ܷ��}���+�51���H(��u�-)�t��������Uzh�::\,�t�ޠ���E����s��0  zɁO|�'�TA���1'OZo�0�������̌ԇ�zL    IDAThX�0E�ؔ7IbR    :GK   ���Hz�:���8u�	*33�̄�¶�wxxX�D��i�+��:¦$K%����?�c�n��:�L<��m�����g4��gY�  �T�������u��H&����{<O�N�f�JE����(�����~�   ��Pp  @'��$�i���E����m.����+��59zEᮻ��f�0�Ϳ�Kz�_���{�&pcG
7ܠ{>�)��ۿ�;   ЕN~�˚���c4E>��Z����nW�v��ce�6����u   �RX	  @���:�@7pu�{��{��E�x<�!J���X2��^`�����O�T���
�����}������K�����4 @�i4t����$M�n[���̸��D�؂~I�   \
�6   �T���t����KK�1�lu
],����|ʛ���}�YG�@�H��w�[�~�����g=����=�� �u~XS_��u���}_ccc��b�Qz�vN�k�O[G0��2`�+)�   <+�   �DiIo�t�*���L����?22�(b�
W���d��1$I#��������6�g<C/���U���݊�; ��q��_�z�:FSDQ���a�=��	�.�z'���!�MÒ�d   x2V  Љ�!ik�M�a..ڕ���#����b������A/��P/~�i�0���?����~O��,p����u�g>��7X�  ��|�N���e�i�٬
Oo&�'��~���a�}@�g   8_`    x_�;�C ���E��ܜu3��+��6��d2�R���D�5���Ӊ�����t=��U�����g�_{����?���G��?�鞙
�S<O���.��y
2�s_��"����l��<n��L�;F}}jl3j}uU�J��ժ��˗����Ը�k�����瞻\^�ZM��e��PuaA�T=���%5j�m���p���Hw�}���n688���U-_��	lN�p��B��:�m���
I_�   �E�   ��%�t�*o������q>�i||��"���ݦh`@婩�����io~�����\�\
��z��ަ�3��o��Z�������>�ɤbɤb����>�R��K"!?����ףH^ɏ��G�bg�K&��bɤ�)H�%�?�5���cv���r|�R9W�_ZR��X/�k�Xߨ�U]^V�ZU}mM�rY��5�VVT[ZRuiI���WWU]XPmy����T1 Zm��?���������Q���<��������q�ҶEŢu3�܃ PE*�wb ����(�  ��Pp  @�y�u ��Ppw�f'Ѝ��)�D���t�:�g֖�K��j�G?��-������~�s���~V��o�����i���(Z/����TJA*%�l9�LQ=�J)�ɜ�?�T��l|��:���V�����ᗗU]\T}ee��_[YQua��}g����������_0� ��؟�y��%)C�������jp�ж}}��P�K���ʎܥ�]�(�[�_��%}�:    Qp  @g�Wҭ�!�n�L&�#����(���c�N�ې��t�}m)���ɟ�s>�!��b��LFw��oi�����ߩցE?�d�뗾���K%E���)<�1���(���s�Hn�=�����6��g�W��U[X��ku~~��kezZ�z�	" �b������J��m�iR��t��)�(�����Zsp'�z���ҒbH�R�����t�J��   �D�   ��_Z �����Y�f�6�=�N���6�h���oVr�.�<�DK�ߋ�t�;ޡ�|�%���u<���7�����k���Q�0�W��)�f�f7
�a.w��~�%�f�..����Ri[�ۨV7J��'���T��UuvV�UgfT��Uev���@7k4t��7]��X'i���-//kii�:JW
'�������]<^4�+$]'�1�     w   t��Kz�u���`���+�c��FGGۘ=��Tz�Ku�S�j�S��y��i�9�i�s�P����g>�o��o����}��٬���KNS?{��D�h`@�6�)�����BA��ɁOvvR|uaA�)�O��������˧OK�F�� ��䗿���z��X�:JS�������V��Q�N��zIezZ�]��c�q�x���Hz�u   ��;   :ůk��)�-J$����	�����ollLA�G}4���_����4��W�����+��i�@'��@��A���O��|E���m���
��(��W��+*d��ql�٩�Q��Ծ}W}|�\ޘ�^��Y�?;����*�:����zI~zZ��5��6�) wU��5�侮�u��:{2��Ç��t��������LQp����>$�u   ��Uo   t�QIX� ��kv��U�VV�c����b����[���cc��z�����<��?�sz֯��baؔ������b��P^,&?��?֧��7a��o{����5:v��V'�Q���⃃Wp��^|?}z}���*gJ�k�N�r�}���ևzԩ���+�KR:�V�X�����"��#��Pp�� t����H���A   �6
�   ���t+��\��.]���L&Ub"6Z`��/�q���}���w�lR*`�/��-�_�����/����g�9rD�J�����ߘ5��e�MN�2=�^�?[�?{����ɓ�-/�!8�]����+�=xbe�T���V>�{����T)�[G ��/K�-Ik�A   �.
�   ����F�@�
�@a.�_Ief�:���I��|���証�&
�2p�=:�����wM�I������_��d��Xl��~��~������H$�w�^=��Ze�2�&��RJ��+��{��Ֆ��v��&'U>uJk'N�=S�/�:��	�pOuqQ���=9���<���jbbB�Z�:NW��.h.Xs���H$�# ݬ��u�?4�   �Qp  ���K�t+�\.����'�>22�(������_�r������&�E���P�Z�=�������"{��}��@{���ѣG���h�#b�R��)�o�eS_[[/�OM]X�?qBk�N�|fR|�^ocr��N��=Yp��(�4<<��G�ZG�
.�+�ܙ��دI����u   ���;   ���: ��\\�sy�{�������f�Fi���W�Z���/����3s��酟��2��-L���y��ϻ�Qj�ŬSn����ɓ'5��W :��+�{���w_�1�jUk�Ni��������Z=s}��q�?�z�������~�[�Z*��jqqQsss�Q:^��ȏ"'�Qpw��dO�t����   7Qp  �����AR ���b�����sQihh�0\�ڷO��P����M=~���O���������й<O~�+�?�k�ۇ$=����b������� ��xA��Ȉ##�}Lezz��~���z���W��ۘ����ǵz����QZfxxX���Z[[����<OQ���'���]muU���<v$�y�h�!
�   0�۫I   �t� t;�*����Dg&�{����1��o�����w��׿.��W|�ೞ�~�
S�6%�	�[/�G����*�J�}_����Q �)�BAa����o���������ǎi�����ǵz��V�U�I�h���~W#=\p�}_ccc���P�*��]:Zp��ON���Y�0��13��t���   ���   +O�t�u�۹�X����L�}ppP�D�8\���������_��e3��^𻿫X<��dh	��(�o�ϟ�N�}ӊŢ|��	GU �K����Z������W�v�V���ѣZ;vl���v����r������?j��c�T<W�T�ɓ'��t����\S��V��;���$�_�[��   �=�F  ��$1z�!K�.ܣbQ�LF��ag���N�����%�Q������W,��a[<O^�?;�=�֯����P�<�=#����}?~\�F�: �	2Oy��Oy�%���k���.e����`B5�h�ᇭ#�E�P��⢖����t����Е�i�f(�M�:I�R���P   `��;   ,Hz�u��R)�mW����`&Q,jdd�:d2���#�����>=�#��%��xA�1}��;S��.����}=z��; \F��*��*s��W_[��#Zy≍��#Z}�	��<I���z�*��
��������8�Z�f�#�Ţu3e
� v.!��~�:   ��J   ,�O+@�6�����z�l��ص�*��
C��P��~��}����]w߭���<�MY���¾Q^���R;��t���>���Qr�m��q���V�k���z��>����������'$���j4���#���o��� ��Ȉ�9b�#9=���]�(�M�+�>.�j   �`U   �J�%�@�p�����lZRq����y�����)��뎏}�u;��Fyݏ�/(��w�����Ȉ�;f z�EJ]s�R�\s�}�J����Oh��!-OL�<9i����9Qp���g�r9���YG�8�������̸v�h�QI?/�O��   ��  �n��4l��M����ZG0H��}���9�0�s��5��B�<�wn�y���(���=%�˩�h�����Q ���a��޽J��{�}��e-OLh��!-<��C��/�;�kT�Y>x�:B[kyyY�J�:JG��E�f\���0���<�w   ��c   h�wY zI*����VUGf����X�:
�d2�ݻwK��VR����x���x|��~f������M���U��u��I�( �X*���nR�M7]xG���cǴ<1qA�}��AgO��f+����}����СC�Q:J,�V,Wmm�:J�U���#�J&�܁�M��$}�:   �@�   ��<Iϴ�׶[.;Xp��XG6���K�����Z9|���%xaxa���WNT�Y�BA�ZMSSS�Q  ��}%�ǕW��;/��:7�>�}bBˇ�����ѣj�jF�q%�R��ԉ��TJ�bQ�O����Q�|^�'�c�]uiI��5��u�DB����1�^�^I�`   n��  �vz�u ��$�I�m����PR��u
�0E�������g�Q��޽Zy�	�WW���g�:T����J%�j5�8x t� �S��[���n�W*Z}�	�LLh�l~bB+����d��T[^VyfFQ�`��J��������	�y�����>�=>2bÄk�!�6�YIC�؎   -G�   �2 �~�@�qm�Υ��'�p��w؊�bڵk����CI^(�g��N�Pun� ]x����ϿD�S�@�CCC�T*Z\\�� �&?�ڷO�}�T|�}�S��|�\�h��Ǵt� ��6*�<�\���<���jbbB�F�:NG��y�f��S��u��D��!���A   ��(�  �]�+ɭ&.��-��ly�rZ_1:��;�x��]�v)���?���U%��ډR��Ƅ��E�b�x\�3Ev/��Ȏ��<Occc:t�V]�	 z\T*)*����ܾz��z���ǵ��c��P�\6Jڻ�&'���F�m�H$T*�499i�#�ܫx2�v>��-�>*�j   ���;   �!��F�@/rm�Ε�{\R�I�Qp�����M��	s9��N�Tu~���v(�(�����Tv�����A��k׮]���P�R�� h��Ȉ##*�qǹ�u�9r�����Zz�q�>�F��v�O���`�X,jqqQ����Q̹\pwi7�'s��&��^)�ϭ�   ��Qp  @;���1�@/J$����EY_RAғgESp����A�r�-}�J����ϫ|�j�eϓE��0��<I%�z�  ��Wr�n%w�^�⍛땊V&&�|�}T�h�Ǵz��h����FFFt��A��_���u3���v�h�_w   �w   ��;� ���<�&Q���T[]���rY]��z�Tjw8���_�bq��K��ܳG��e���U[\ly������<�ɧ� �)�kllLO<�u @��P��W���Uz�K6n�--i���/?��}Tˏ=f�a�����Z,�"�J%�tx��$E���̸0,�r\:n��~I�H��u   �.
�   h�[%=�:Ћ⎕6�ss�Z..)s�����vJ$j�s�R)%S)5�UU��U[\\/]���E�bg�쉄b����C]�~�LF����� �p�tZ�[nQ��[���hh��1-���Z~�1-��?��׿n�T�#�+
ZXXв�'?��u3.Op����{%��:   z�~   h��Ir����k�t�/�{���/L�S��I��V�b1�������>��
�PP�VSmeE����K��F��F�z�7���XL~��ϛ���bM�t������jqq�:
 ��x�ccJ��I/z�$�{�y��}�8��'��522���^�[G1��K���]�:���/H�5I�E  ����  �V�Kz�u�W%	�m���9I�e�s9�����kttTa�޼XLA&#e.�gA�^�<ϩ]*��y����QMLL�\.[� t����)��'�c����XG�Qi``@����QLxA���OOx���)WB�h����J��    �M��   \譒��!�^��"]//�F�.]�=s��@���q����\�t�N��Sn��b����ƚ�� �=��y�uS��B��ܱ����u�rY��e�&\x���   -��   Z���^�ڢt�G����JmJ�����X,Z� p�D"���a� �.���Z��u3�J�:B�8�K��'����u3���&R��u��]+��   �M�  �*wK��:��\+�W��#�DVRx��D���bAhdd�:�K��r��r�1  ]̋�w��)&�_ �"8�K��ܥ���J\;vy�u    �&
�   h�wX z�k�t�,����6�����gttT�X�:��VE�1  ],���'���h4�#t�b��D"a����~�fzuW��q��`�e�ƬC   ��Pp  @+�~P@���k��<I�3_�&*�Z�.+�J���1 \�����m�_  .�r�=��g���<���Q�`�Lef�:�	׎�FI�l   ���;   Z�]�X= Z̵)T��y�M�'i��x�b��Q�D"�'P ]!�L�ȿ �m���:�?��Б��s�-�|�:��^�Y�;�Y[  ��(�  ��<Io����)T�F��cCI�-<�	�h&B�g``�� `[������}vު���: ���x<.ߧ������C   ���i   ��rI{�C .p��V]XP�^���4y���Y��@���a���N�Y�^�y�FGG)�  ���r������y�����c�M�r�}f�:�	��{�u    �VB   �l�b p�S��4����zE�ض�h�d2���~� �!�"p� `������Pp��T*�\.g�-b��0��a��	�[�� c/���:   zw   4�.I/��"�JYGh��ܜu���I�j�8��ϴ14��y��me ��P(P� lImi�:�>O]��Аb��u���<��Nq���|I�  ��A�   ��I�u�.m��+����A���h���řb	t5��4<<̉* ��i4T]X�Na&��g���b�������j���1LPp����"�   ��  �,���Z� \�R��&�%$���}Q���(pX<W��&���H$T(�c  �@yjJ�r�:���/7%��)��Χ���j�]�*33�LPpڪ(��!   �(�  �Y^!i�u�%.-�U�|��'i�K���@3��q###L|zH�TbG �U�=j���6oxxX�����N�{`x�v�t��o�   ����G(   �No� �&�JYGh�n/��I
���Ӷ�$�|��}��x����!� �G����fEQ��;>Eܫ���]4vC=    IDAT��Z�   @���  �f�t�u�5.-�u�@Rv�R�@�b1�J%� Z �N����: ���^p�ZG�*�b��w�	.�Wff�#�p���!|I�b   ݏ�;   ���"��K|�W��1ڦ�����|T(4+
600�X,f@���v� ���9b�ܷ��<[�h���{�	
7H�@   v��;   ���� ׸�8׭����νsy��E���=-�"8!
 p����Q���N�,�J)��Y�h	�O"w���H$�# .��S�!   ��(�  `��t�u�5�T�:B�4*U���clYLR�',��,p�����(� �ӨV���c�1̄ehh�'w�
��������XG0�ڐ����u    t7
�   �)R\�>խƲj·���؁t:�L&c@���R�d �a�T�\��a&>8h�k�b��|oᅡ����[���w�̽�ƬC   �{Qp  �N�%��:�"�
���y�[IJ7�y<�W����ع��!� �(��)�[�  t����:�������Z>���rp�ߌ�ֺ��w���&&��!   н(�  `'�,��V��.���\7��%5c�� ��׃[£=(���<�''� �o���:���޽��^/�4:Zp��˪-/[�h;����Ԝä   pw   �ă� W��8�m���fU��|�I�XG `���ϩ�	 �+s}�{r��]/�L*��Y�h*W�T�����v�7L�t�u   t'
�   خ�$=�:�*��*]Tp�%5s�?*��lpI��(���S� �Ԩմ���1LQpo���A�zhw1��ڎ�� so�   ��D�   ��v� ��\*�w����f.���b���<OE~v �e2%�I�  c�?��j++�1�x������1zB=�C�����w��^!��_�   �6
�   ؎P��Z� \����n)���2M~Έ�2���� $�� ����:������ ���3��|��r��{��Tff�#�]���],!�u�!   �}(�  `;^%�w�6]ȥŹJ���%yM~�0�o�3��1��Y�t�i� �y���={�#���4<<l�)\��^qp�{<��S� ���:    ���   �o� �.�HXGh��u��Ji}Q�E�B��,��*C� :'� ���=��u
S�k����sR���٬u����������lI7Y�   @w��  �����! ׹Tp��	�֧��BH1[T� ����sj� �9��:7g�T�O��Г�~�����&\:�t�7[   @w��   ��VI���9�0�h����>I�=7ܱ�tڝ� 6-��[G  �����#���F�=)î�%�O&�;:���	�C�р��:��0*   zw   l�� �3�Xk++j�j�1.+�z��e�O)[��v ���߯ �c  �l������LF��1�=�P((�򂸫S�]-��r�pC�~�:   �w   lų%��3�\�<U����pE9I^�?��xh�x<�L&c@�<O��� �Y��f��]��27�(y����6��U*��c숫�z����u��K&�� �{�u    t
�   ؊_� `�+����u�ˊ$�Z��A&����:����|>/�� 8c��U���R�y*�Z-��*�j���
-�KR�Ç	�܁��RIlY	  �M��  �͊$��u �\)�wr)��K�!�elR,S6�����A��	 p����e�\���#8app�:¶�:�]����Z���h@�Kz�:   �w   l�+�d�c��0W]X��pII��ƴRT,���+�٬|�C< ���� �f��;��$�Lv�ItA.g�w �^o    ݁�O   l����\'Np������9��Ci�f�R)��>= `�:7��G��a*�d����R�$��cl������z���C   ��Qp  �f�%��:�s\)�u������
mxt�d2�B=�M�9<� \1��H��uS}�x�<v8j�(�T��ϯ.�;q�@��r�"o�   ����   lƃ�X :DE�Y��m�}I��|=*��J�fLo����]9a �y����us�g>�:�s�Ŭcl���;���t��h}�L   ��hD   `�^k �9.-�u�����A�	����Ͷ� � �����: �Eժ����c���z�u�������[B��-.K��nIwX�   @g��  ���V�m�! ��ҶʕZt$e��z�q5�l֙� 4O.���  h���}O��y���(R��7[�pR>�����>y�~�r��w�#��:    :����  �o����Ң\'Mpϩ���Ƌ�6����lG:�V�1  -p�k_��`.s�M��:��<�S�T���i��)p�ĿN&�..K���J�3�   �v�   p5�� �B�,�5�..Z����Ғj�k2�W�ŔJ���@/�<O�L;�$ ���o|�:���3�i�i}}}J���16-�﷎`�2;k��9�t���WX�   @�bT   ��NI�Y� p!W媋�R�nC��jK�������[d�Yy^;� �K�٬f,6�}�kk����Q�����F��ڙ���S]Z�j5�VWU/�ըTT_]U�V[���8�=��j\�}au~�ү���z�r��jU���n�|_�M���Ӓnf��HlL���w�O$��E���|��'���XL�TJ^*�Lʏ��G��dR��� 6k��?�ڱc�1�eo��:��u��A���j��^.���*ߑ�K�;�Ҁ.�FIa   ���;   ��M� \̕E����-�������%(�2�٬u ],�J)U�U�(���yՖ�U[YY�,.���������UՖ�T]\\����������WW;�=\/����%�dRA_�z	>�T,�T�ͮ��I�����s��׷~�d6���z��׾f���Sp� �DB}}}Z8sBS's��.���9r|Ir�XЅ^"� i�:   :w   \N(駭C �X<��J���,��GŢ���[A�d2i@�<O}}}������&iT���ϫ�������/.RH�`��%Ֆ���\�t���{,�Q������\N��K��)��W�Iu]c����:����7���s���Z\\T�Ѱ�rEA��g���)���6܁�Jz���d   ���;   .��hXȕE�N([�����n��S�pu�lVSX�P6���ޡ�kk��Ϊ:7�����+����Ϊ<=��쬪�����ʊult��e��-~�����lVA.���� �߯h`@a>��XTX,**��L�7�|�{�:����>�:Έ�H�lVsss�Q���	��9��C��+�Ҁ.�ZQp  �%Pp  ���: �Kse�{͸���fz���bp�L�:��L&��T�լ����ښ*�O�<5����*33�3������(���4�����M����{�TRp� l��bq�v��M3��k�#Pp�,�RI���=���{'h'
�@G�]�.IOX  @g��  �KIH��:�KseQ�b�ؚ�݇f��qe��+�ri��V�<O�L��'�v�z}��>=��S�T��^/��>�q��}��%�@���������W|��)��
���B���RI��!Ň���b�6��ө�|�:��X*��ӟn�	�P�|^����Q.+�Y��n���{�0������u �%�^�Ǭ�   ��Pp  ���J�a��J��r��/)k��Z�f	\B:��ǤS M�N�)�?Y�����*�:��SZ=yr����e��̌��i�j���?������(VbhHQ������
K���Ţ<�o_��|�����a.w�m��=;�������:v��O.�8�0�Hhyy�:�K�yQp  ��p�   ���  ./�[Gh���kg$YΈ^dǕ��i� zH&��9���5�MN�|��N�\/�NNjmrRk�N�|�ʧO�Q�ZGp�z}����.�	�E������z48��X�z�DA����?���p	�XL�|^SSS�Q.)���/4�Q�ε	�w��=C�S%��:   :w   <Y��Y� py�Lp7Zl������q9��Q�V,S"����u���׵65���ǵv��N�\�z�V���䤓E.��ju��~��K>Ə"Ň��W|tT���.A��Ϛ��.I��ޱ�Ţfff:r���
�IU,=�:�@G{��Y�   @��  �'{���u ��ʂ�����K��K���
��:���d���^[^�(���8�ճ׏_/�ON2y���e�>��Ç/y��^T~O���tޒ����	��##J]s�u\����ɓ'��\R��9Ypw��?W��]�բ�  ��t��8   X�y�  �̕���|�_3&)��W��q)�t'�t�5�LFSSS�1�z]�'Oj��Q�=�գG�r�V�\���Z'����Zx�-<���w�����e�3��]J�ޭ��݊%m�L���a򺝦p��p������V�R��r� ������v�\��r<�b�Jz���Y  @g��  ��$�*t8�����N��.1��F�@+$	���z���ת..n�W���c����U��� HZ?	��1�;vɻ��A����(�'��Ur�n%FG��b-�t�o��5��e�w�eWqv���,�٬u��U�������Q�ƅ�i@xP�  pw   ��%��! \�rՅ��h�kv��vI
���KHM��<�S2����RS��:?�QZ_��$v �E��I�''5��p��^(>4�>�}|\�k�Q��k�SbtT�m���w��r'��a,�L���϶��M��r:}����u����u3��yE��u���;T����Iz���  @G��  ���: ��s��^[\l�kf%m�^�<^,� ������k��O ��J��^.k��!�>|Qy}��	5�����ѨV7~G�~���K��ܳG�k�U�k�ڷO�}��T�}���U��J�s�+?��c`<�S�X�)�1G'�KRev֩�;'�]aD�]��n   �(�  �qI�[� pu.L������Q����w4����x ��J�.��:?���t��F9s��-OLH�z�C@��--i�G���#��vm�Sg.ɽ{���$�����_��A��S|��#`r�����T�T��l.�W��#���Ӏ�zQp  �(�  ���J�C �:&�W��z�2�]���~��@�*��N5�u���[Y��?�C-:��C��|�ꫫ�� �I�Je���4u��dRɽ{�ڷO�T[^�	�A<�W��;�c`�Nq?q�u�wg�p<�?-��8�  �q�  p�+� ��0���.J���;iz�tf�;�$Lp�m��ꕊ����emM�3�������5����g�N��8����Nw�����H��D��L��.˒l˒�<�|���T���}�d��̋d�T���IR�7��U7sS�Ln���)O%�;q2�܉�+o���"%R�A �z��}_ �H �s��~��
��ϏZ�������2 p'�ZM�o��ŷ�6%1��Snd�tl��ࠦ��3�=[���`Lkv�t�X1�H�ݒ>-����   �,
�   ����N�`c�L�j�XpO��vI�����	�@�\�t )��
uE+��FC
7|���q
� �Ty�9��I���ww�rM���E�  �y�   I�&���Ѐ\Y��k�{Ҧ�KLp��\�����Ⱦ�����bB  zo��J����	�ss�#Ċsk U�"������\   �w   H�WM �9�,��Up�W���KR@��6ꀻV����{�l�Ⱦ������1 �ґ#*NL���mJ�w�X���*L@�>nm
� �k���%���    0��;   �I:i:��qe1�C�ݗ���W�:&���(���"u�u���
�uE�vl/?x�2����y  �m��ϛ��J���5��Mǈ]{~�t�X�rM���E�  �i��    0��Z�yHW��qLpO��vI�����a�[�VS��-�>��ٳjMM���k�]��|^����  l��sϙ���1�=	�J�t#Z�Mpw�`�WD�	  �i�  �WM �y�]�==~R��KLpǭ2��r��� �,
C��_W���K�ׯ�^h_��=���  ������Q�1�����f��c(;0`:��ZMQ&�ǥX,�� `k�Jz�t   �C�  �m�$=b:��se�T��I��.1����r�d��_+����P͙UϜQ������H���n�  ����ϛ��.I�wW�Ԛ�5!6�\S,�    s(�  ���Zd %\�6E���jώ�K*���;����X�+�6 ֋���gΨy�j"����B� ��?�Y��E���
��h������#Ć�k �����)  @�Qp  pۯ� `k\�6.-Iaس㗕�a&��f�\�t ;6��;�ƕ+�-��001a:  wT<p@}��o:�(��hxx�h���	��$ܨ�'M�   �I^�  @o�Hz�t [�B����سc{��{v����ey٬�H�,�= �֜�R���j��lJ�ؘ�a8  �v����聡�!���M&].�7ggMG�M�w �-_3    fPp  p��&�+�@ʸ0m����Oo4	C�H���Q��y5�]���t�M��yOP �N��������4h�|8�T���i�&�Kn� ,���    0#���   譯� `�\X��������ד#wOvh�t$w }�fSճg{��Y������  ���x@��q�1�#����<3K�.OpoQp�|�>a:   �G�  �M}��6���r9�z���Г���m+(��f�L��Ӂ�	�ΝS�l���me
� �����K�#��� Ѐ��y��	�T.\W,�5�   ?
�   n�I�! l���z5�'G��-ّ<�lV�L�t ��Zno�MG�&� �(������c��FFF������o�kw���z�t    ���3u   ���  �ǅ��v
�EIi���w�,�͚� `��v[���u:���Xy�>�  ��࣏*;<l:z,�˩����陌����_7:�������  �xQp  pON��C ��R�E�=��%&��V܁t��H��Z��tEit�t  n�祗LG@LFFF��n00`�uMkQp�_3    ��  ���$��bX����n��+i@�7�}�t �иrEa�f:F���� �0^���g�51)
*�˱�n�т�k�]X�+�    ^�  ��U� l�q�./��ez�$e��LG@�Pp��������]E� �4#�<#�T2121�=�Tb�$[-�����qap`�OI�g:   �C�  �-I/�`�\(�w���v���b׎�{�.�cm܁d�:�/]2��(� �f��/������e
�X_��	�R�$w �<I�t   ć�;  �[>#i�� �/�^���];V���KR�R!nB�H��Ԕ�v�t��˖J��� ������x�t�w��{gq�t��PpR�WM   @|(�  �嫦 �&�o�/)m���i�䣗(���Zj]�n:F��.x �e��?//�5���+����;��4�݅�j�垒�	+  �#(�  ��� ؾL&c�B\X�+l��r���LW��LF�B܄�;�\��i)�L��<;�  b��/�� C2�����b{=�'��Tpg�;�zYI_2   ��  ���%�c:���f��dRU�޲v����H��ʑ����Ph�M(����j�Κ��SLp $A���?���0hhhH��rv���?��y�bc���_1    ��  ���� `g\�2���԰���U���C���?��    IDAT*r ؚ���VOo�$߁� ��}��`��y��t���j�6�.\[�I��   �=VJ  ����@ʹ0e�[���]9J����1��� �Q��w�y٬�  �y٬�����H����X^'�K�>p���Ұ�4��X�"�i�!   �{�  �0$�� vƅE�n���x+����6
�@���u:�c����Mu �d��g�2	���T.�{�:^���M~��Я�   �ޣ�  ��_���
`�:](��u�w܌r;�L�9�b�j� ����b:ddd$��	�Ӹ�ε��MG���#����    �=
�   nx�t  ;��"\k��@R�;Qb�4	B�H���T�Z5#� &�����c����)�˱����������nziQ(LG �G$�k:   z��;  ��IϚ`�ྱ>Ii�3�7��$�+��%
�  �F_~Y�X�ĭ���z�>ܭ����!�t    �W�   ��yI�! ����¶֓T�^��Qp��(�	Ej9Tp�)�  L�d���_6�	T�T��~O_#p��ީV�(2#.\[�   �Qp  ��WL �.L��,-m�gKJ�I��� ��jUQ�e:  �|���7	�y�{����Ga��w�K
�U�4b:   z'�k�   ؜ϛ �;\X�����/C6��G"G��i����Oi�i6MG  8j��WLG@��t�+W��ήǤ��# �x�^6   �C�  �n�J:d:��pan��
���F�]v`�t$w Y\)��2� `@P�h��L�@�e�Y������A��t��y�b����1_4    �C�  �n_1 @�����f����&0�7��$G�VS�n��+
�  �~�K���;344Գc�Lp�^�<*�E>+�7   ���  ��^4 @��>�=
Cu��-��/���8�����EQD�H���.�f�f�t ��F�l�\.���H�r�ݡ��.� 2$�1�!   ��  �U���� �����Ғ��BoYR��qb�0 ���#�,o�w @�*'N�t���H������傻K�ym��8��   ��  ������ ���	�-�LFR_����/��	�1�0Lp�[-������� �۾�~�t����<����.���m��8���  ,E�  �^_6 @w
v߳ҩն�3I~��Ď��XK��# �s��s����~ �9��A�<���H���߃2z�g�-�����^ۯ�zH�^�!   �}�  ��Y� t����3�ݖ��R1	��tLG �����lИ�3 ���_��<��w�}���]?f&���h���P����k��2�^6   �G�  �N�I7@wپ ��b�0���M��Lp�(��EѶv�Acv�t �C����H�R��|��W�L�O��C�^�w�8v4  �w   ;}�t  �g�ʝjuK����xd���5Pp���뒣�6��MG  8b��I�2)544��c��]��N��ҳZ��   �Pp  ��� �>�'��[(�g$�{%v�N�ÝQp���W�h--)l�L�  8b�W�t�X�R���]=f�����Eۡ����� GHz�t   tw   ��Iz�t �g��V��E�uB�4	D�0�Ղ{cv�t �#���y�Y�1�b��i``���tv�{����4#Lp����    �.��    X��$��*
�#�T{qq�ϵm����y؁�;`VX���`w @\����<�o�F�v��qW�;S�)�����    ��t    t݋� ��'�o�H��}w�d)�c�s�fS���6��LG�+2���e�Y��2�//����+�y���ok�K%yA�L6+�PPf�go�����-�(Z���Y\���_�����ӑ�h�9�Z��V��Q�|#g������QX�)l��?�Z��X%���W�b:,P(T(T�׻r<��{vd�t����X�I{$M�  ���  `�gM ���å�M=���&ܱ��7����te��+�# ��\N~_�����r����������BA^���_�>��+��W(0��&a����T�h�S��������ZM�jU�jU����U���:ժڋ��ϻ���u�UE������'�Pq|�tXbppPW���	�����ఌ�/J���   @�Pp  �˸��M� �}��)�͚��S�ju��d$�z%vܱ
�9����˗MG@��~eT*
*eW>n�:�￥���SJ�o�F�n	�M���o�h��������:��˓恘��Ϳi:,R�T499�0w|�`e��Rpg�;`�E�  ��  ���� ,��t��&&�$����l�b:��j)�"e2��ĭS���`��ŋ�#`�2e���RnxX��e��)�k�G�������y�S���\N�]��۵kK?�ᭅ��Y5�_WkzZ���պ~]͙�ffV��:��.`��'�������x����>�����X.߀N�����Yd:   v��;  �]>o: �ޠ�������X_Ej����� $N)l4L�0�	���J��ݻ\T޳g��Ȉ���˟W�칡!
�芌�);8��ࠊ���E��쬚��j_��\���QsjJ��5�^UsfFQ����H�L��o�������`w
�Lp�w�j{$=(闦�   `�(�  �##�i�! �F�P0���Z����Mm�&`�;��j�(�1[-)M�0�	��V'l��Wn�.eW���޽��ݻM�6tc���h�ϫ95��q횚SSj�|��u��e��v�]_��J�����ee�Y�Z����])��0DpܗE�  �
�  ��a�! ��oQ��\(�����䱍W(ȳ��/�o�� [��#�i4T�~�t�T��[���ޭ��=���{�*72��
�.P00p�rs�n�53���+jMM�~��/�q���W��y�����1�F7���7�a:,V�T455��c}}�x�"o�q���w�z�����C   `�(�  ��K� �����S�!�	.O���(����Y�tI�"�1�+�Qn�.�Ɩ?��S���J�=��3�H�L,��gϺ�	�M5�\Q��U5�\Q}� ߼�k��,O*/�ױ��]y�Ns�QpW&#�TR{q�;�Rĕ����� �	-oz��B  �x�  ���  z�`y	�S������e+��`�Y@��f�tc�Ϟ5��LF�ݻ�߷O�����7�:?:ʮ+@x�����*������̌j/�~��.���~�W�*�tbLe2����}��1����r*�J�np�a#A?w�1��^A�3���A   �3�  ��'�� z���R��1�0!��7	F��������3��2��ܮ]�����R~ttu{~t�;`�����x�۾��j\���J��R|�]����j��Hl�������_4��J�]�/w)Qzt6���(�NxI�  R��;  �^��Í��ŷ;-�f$��;���t$X��TE�d2�� �p��~���;��r*�u�
���Qؿ���e��#0,�N�uך�o�ͩv��j~����?�����߷a�k_��7�a:���/�����N�����X�s�   `�(�  ؁�u��l_|����$/�(�su��E���
���(��VK
C�1�IK����?*���o��{�*����@����+�?��m�[-��(��;�ڹs��;��^7�6���������ۦc�1�穿�_����>���Nka����R��m�%�$阤]��L  ��Qp  �çM �[�/��iJX9�&�.�c�(�����i4�x����Ri��~s����r{����Q�ߣH�+WT��CUϞU��YUϝS��Y5''̈́5(��:����~��LG��*�ʎ
�.����2��8���iy0��m:   ���;  @��H��t ���w_�ݿs�α9�F�t�a�e:�1�g�(�yz}��US��A�TqbBŉ	�&&��5 �H&�¾}*�ۧ����[�juy����k��-�9����~�������}���|��Q�R��\.��6o^ty���Ғ�� �y�B�wn�(�  �w  ������Q �����:܋�2�F�wl��;���׳c}}*8��]w�|��J��p�]*:$�	� ,�J�;vL}ǎ��xgiI�?\.�����+�K��(2�vg��zJG�w�۽�t@����������e���[�z�gl��d��f9�����    �
�   ����  z/�˙��S�uPK1�0���p؜Z�f:������;��� ��¾}��Z��^:t�i� ��\^��ޞ���������ϜQ{n�Pҍ���ա��w���LGVn��8\p��a�6�|��;`�#��K�`:   ���;  @�}�t  �g}�}�o ����|
��@��Q�ٴ�� 	\.�_{�M=�/�U��P��A�Tqbb�c|\N����8�ʉ�<ޜ�V��-����N����vN�PR)�T���_�]_��<�wC��r�m��=���ۋ��#����������t   lw  �t�/�� z�����&��0�]���~���j��;��т{kiIsgά~��<�GG����Tb/<�������r##ʍ�h��GW������������xs��!���]�/�,�P��k;Q�T499��sy��z;�����l V}N�  R��;  @�}QR�t �g{���;ܱ�ZM����c v�"E��F\��/����ݿ��*NL0� R����w������Ǣ0T����;�h����;j����J�k�����_P�}��4:���
�[�v��n�u6 ��1    �G�   ݞ3 @<�٬�=��؄��ʇ
�؄j��pX.*�L�0��/~!Ix�!��5� ��Sq|\��q����Wo\��\x?}Z�3gT�xQ͙�gg6��?�)74��ؘJG���{4p��r�v��-ۖ�fU*��|>�;\pwe����� ��t���L  ��Qp  H��M ��-�������h6�j��
.� ����vI�Z)�'&' �J~lL��1�<���(@��\p�
yA������X�EQp  H%�t    l�I�M� ��N��H�z���J����wlV�V3�Z�阎`D��h���$I��q�i   �k``@�Lf�?�\�2�������:��|�t    lw  ��z�t  �y�TX�*
�կ�|sqb���0���թ� ���	��o���ʟ/Lp  ��}_�����s�ft&��Г��~�   ���  �^�1 @|l�,��XiץiA��H�EG&���:�����_�$�TRnd�p  ��T*[��x�Rp��:���t��   �:
�   ����  �c�d��O3r���;:��l6�l6M� �����?��$�t��    =���'��ڲ���ێ�f�u6 k���    �:
�   �4!�� �c�d�v�����:Quu�۷��4=��(MG�]��u]�IRq|�p  ���<O�[�A�/�t��G:��R���s6_g��gM   �ֹ�   ��L /�'KuW]4��&�c�o��@w�Xp�������  �k��r�GI�-
C����=g�u6 kz�t    lw  �tz�t  �y�-\��:#�
�ف��2�jU��� #\,��������m0	  @o��ey���]�!����a6_g��QIGL�   ��Pp  H�'L /��N��p��{'�./�c{�0Tu� ����(u�G?Z�:O�  X��<�m�<pt��$u8��:�u}�t    l�k�   �t�t ��<oKS�Ҧ�Rpwmz�$[�"����� +�Vp����՘�]��	�  �v�[8w���^\4��(�Nz�t    l��	   {� )c:��ؾ�֩�$9Zpg�;�aaaAQ���Ǳ���?��[����e(	  @<���6=@���A6��t �{�t    lw  �����  �e}�}iIyI�� 0���n�Uu`�x nQ�c:Bl�0ԅ���[�  ���y*or2�_*�8Mr�(��~����K�0   �G�   }�4 @��٬�=�^Z����.O���,,,�� �ǡ����Ǫ��|�@&#���   �Կ��]�q�C����7    �G�   ]vI��t ���j*�a���ؙ��yE�qtׇ�����I���4   ����Wf�{�MNz��wۯ�Xw  ���  �.ϋ�p�sl�*���M�0����8��:���ժ��U\�i$l�u�/��Ǽ|�P  �xy��Ri�}䂾>go lSp`��M   ��Q�  H�O�  ~�/���u��	(�c���MG ��H��ʫ��17w�c� �K6|N���;�Ʌ	�� ��#Z�)   )@�   ]5 @�l/��].�;��9vn~~^a�� e��ɟ����   ���߯�&��}}1�I����=g��6 �ʈAR   �A�   =r�6@�l�*U��%N�lbj��0��t������Wu��Q�c   ���T*m�<GoJ�T��#����� l��   �9�  ��	I�! ���R�lVrt����st�st�����=(����w�i6o{<l��  0�o��]-�3���4    �C�   =>c:  3l�*U�Ė�����U��T��M� ���韮�xD�  8�����z�.-���s6_k��㒘:  ��  ��q� �a�T� 8\�6��lS�l���~��>X�{Lp  ��f��o��Z�h��S�[������ lJNҧL�   ��(�  �� G�:U���_�����Ip边�9�ah:�~��*r�O�d��E�v�I   ��o��r�T�)I�Da�N�j:FOQp����    �w  �t�W��! �a�[__��w&��[�0�����@�Y\p������}o��G��"n�  �٨���1%Iۯ�d�YyU	�aO�   ��q�  �L� fc���<�J%�L;�izzZ��[�ؾS���:����w  ��b�(�����O��jA�� ���$�{�;  �%(�  �Ó� 0'�˙��u�RI�穵�h:�1�nu��h6�Zr�� ����������w6|^�jŐ   92����Lx�Yہ�56� �iÒ�1   wF�   1 �96.��X@va"�z\���133c:�jK���韪1;����  \t�����y{ہ�5�|�t f=k:    ;  @���I�Ӭ.�;0l=.ou��XZZR�^7H/�Q����6�ܐ�;  pP__ߺ7:�<�݅�A�� �,vN  H8
�   ���$�t ��r9���P(���;ժ�4������S܁��x�]*��?��>�pS����  H��TZ�����v&��v����4    wfߪ  �}�2 �Y�Mp�y��6܁����W��2H''�����ݦ��N  ����3�����Ё�����'��?�  R��;  @�=b:  �l.��\�syz'�"MMM����m�/���z��M?�����4   ɵ^��+�{��Y.$��z�-���  @��yF  �.�M `�M�|�W�X\�څ��O�Co��ͩ�l����e�_~��[z>w  �\.�|>��LF����S����s�Hz�t    �ϮU   ����t f�Tp��T4����#Lq�Ǧ���}M��Ɩ~�����   �Mq�o�I�%mvܳ�z�m{�t    �ϞU   ;=c:  � 0�k>�`:0l=>w���ܜ���@�XRp��H��ַ��s� ������;��Z�@��	�(�    IDAT� $�0    �c�  �^O� �����N��/�<�=Xg:�-Lq�&���#t�����u�ԩ-�\k~�i   ҡX,*�������;���=�w ��I��t   ���;  @�}�t  ��2Q�P(��Xy���D��0��6??�w`l(�Ga�_~����Y&�  �y����鞫wvܳ�z�{�t    ���;  @r�0�y�,�ݶ�w�M�詫W��� �����ǚ{��m�lka��i   ���r�ܽ]�IQd:FO1��

�   	E�   ����  ��e����;����Ҙ��<y���p��Ғ(�����{kiI��ַ���m��   ���~�0Th��`�\o�c��   ��Qp  H�'L �6Lp�<O���]��z=^����)9�199����{@7�����o}K���m�|gq��i   ҧP(���{B�����N�f:BOA`:�dxXt�   �7i   �u�t  �`C��X,��X��傻��T8�W�ͦfvPz\������z�?���	�   ��>��w�݆	� V�$3   ���  �\�M `��yVL����d�B靸�@3����n�M� -������N���c��_�R  ��*}�|�c���(����   �v�  �� �n�! �g��vI*�1���;��0u��5�1�dKi����K�W;>NkfF��.$  H��_��A=���n�@	 ]��    �w  �dzT��V ;bC�=����w��Pp�����:����L&#y�\�i4������+l6�^X�ʱ   �*���r�wx�{���G&���	�   p�t��   ��1� $��mkMo��.��O��Y�/_VĄf`]��Mq�[�����];^sj�k�  H���cx����_�����yP�:   $w  �d���  ���	��ܗ�bN�>�aH���V`]i*�_?uJ���v�����   �n�����N�f:BO�p�@�$�o:   nE�   �>a: �d�a�m݂���w�w�4==�F�a:�Hi)�������O��]=.�  �R��L&#����m����7    ���  �<%Iw� Ҿ]r>�W������wB�&EQ�˗/+�"�Q��IK�����5���]?nkf���  H��T($�}�n�`��_s�u��   �[Qp  H�G%�����O�*�aҙ��`���@\j���_�n:�8�un�J�����Ʒ�ݓc7��{r\  ��)���RIZ���ۯۤ����;a:    nE�   y3 @r�}�T���:KK1&I��	pH���I5�1�DIz�=�t���ծ�{r���TO�  �6��32����0�����~�@�= �;_   ��;  @�|�t  ɑ�iRw,�[����0�IE�.^��(�LG#��_~�ۚz�����;  ��R�����v�ћ�ۖ_�I�57 ]��r�   	A�   y2 @r�y�T6���b��[]߉���H�F��k׮��$����˵_�Bo����5���==>  @Zx�����v�X4��&�p;,  $H�G  �'/���ve2A�V�e:�5�<M�N��%��LpG�LOO�\.���@b'�7��o~SQ��uW����   iR.�U��8z���;�Qp߾ ���$)�ϯ�vpC��R�ӑ�|c=�"'L   �G��b  ����fEjy��Zn,�*
*
��.�*���r�ӫ|�_-_g�Yy��D�Z-�+E�z�.I�t:j6���j�������V�iaa�Y^p_Z�)I���0�.]��ÇW�W%�����O�t�R�_����������  @�W&���Np���$���r��*�����o�\*�n�6\(��n
�t:j�۷\���z����E���kiiIQu�wl�æ   �#��  $�I�`�r��J���h���k�w��r��b�V4���iaaAsss����������477�v��͸���Ŷ�/�މ�ۛ#���.]������<����i�Ip������_c{�������z]��Eu���K���j��+
C�u:
�UE���KK��m����v[�g�FC�7_F����d|_�:��bQ�lV^.'�PP���J˻"��;����LFA�,�X�W((��_*}���@�) ���q]�su���;����fy��J����!��Q�T�u�v�|ߗ�����T*>?��k�7_���������f��$e$qw  @��  �.�M@�y����!�ݻW�������e�$���ڳg���ٳ�����t��U���hfff��6M�I�b�f�:پPz'LpG-..jjjJ�v�20��	)�_?uJ?��ߋ�5�/�|�h���Ya���쬚ׯ�9=���Z��j�Ϊ15����G%����YZR�������岂����~e+���
�����GvhH��Aeؽ �5�(�w���NGQ����v'Y&�����X�^1��kddd�cϞ=ڽ{wjw��<O���\��KKK�����̌&''u��U]�~}u7Q`��%����    ��  �4��t	�@{�������E�RQ&�1-�rY���ÇWk6����ֵk�t��]�tI���S�LZ��M�].��:��w��5
������	i�I�qk�������R�^��u/_���$)
C�ffԸzU��I5o|�vM�+WԜ�Rsz�����j˓�gf���A�����j�=;<���!�FF�۵K�ݻ�۵K^�S> H���.*�jW��ZZp��w�Lc�=��ittT���Ӿ}��{��M]��I�\V�\�����c�v[��Ӻz��._���/j~~�`J��IQp  H�t6%   씑t��H�R����Q���illL{�����[�r��ŝ�~X�T�Vu��MNN�ҥK�x�bj��Zp/nb��咚��ߐ�.]���7܅�U&�Fa����h����_�ޣ�{{~^�T;~��~�W��95������bc�9��椳g7|n00�\x_)��w�Vn���Sᮻ��} �*�b����ZMZg���r]�\.�9���<�3+qn�ٻw�mׅ/]��K�.��ի��.c>%�L�    w  �$9*i�t$K>���Ą&&&��~U*ӑR�T*�2��nkrrRgϞչs�499�(��\[Z��f��"���ʣ8��t:�x�&&&X0��2٬�z�_�k]�����N
�Q��ڹsZ:sF�>P��2{�ɉVh�ϫ=?����4�*�o�
��}�yll�?6&߱� �ts}�{'�݄�M�{����y�������W��H���u�K�.��ٳ:{��f����	�   �,�M	   ;=b: �addD��������O��� X�x��O�V�����:����}---���*�w��������N����sx�ң^��ʕ+3��g���������?0���+W6~R�q��O�V��-�|��=��l�HkvV��Y-������Ua���SqbB��U�� @�����3Il/�'�ׄ�����5>>�g�yF�jU�Ν�|��gϪ�l���4    ˒s�  ���� t��!:tH�p�5��X,��ѣ:z����y]�zUgϞ��ӧ555e4[��6k3���ZI����H���9��y������*c��ޙw����M���2kMpoLNj�7�?�|S�o��N�j lpc
�ҩS�}���T:xPŉ	��U:tH��	'&�s� 0�oh�tcl�~c��������w��5a�J���;�cǎ)C]�xQ|���{�=-,,��3�$I�n:  ���ה   ��:���=�ܣ#G�(�˙���LF�����?���y����z뭷499{�4܋�غ������;RdrrRA�R����&��y�����7Sm�����f~�U�{o���0�n
�M-�:��5����{U��P�������*=��ࠁ�  ��)�[+��n��ittTG�ս�޻�kh���y:p��8�g�yF333z뭷���o'j�O�\Fҧ$}�t   ץ�)  `��M@oy������رc��Sd``@Ǐ����533�S�N�ԩS������m-�۾@z'LE�\�|YA���p�g��ުV����U�P$�"��w����mW��q��f_}����{��|���>��W}�ޫ�訡�  ���`L�^7����vs���ѣLjO���a=���zꩧt��e���{:u�ew7�w   ��ה   �Ӱ�}�C�7FGG����{�Q>�7;0<<��\�?���]��7�|S���=\�K[�=�ɨP(l��w 5�(�ŋu��An΂2�/y����^�n�~��u}��� 6v��>���XP����{�w�}˟�Sq|�`J @�����I���a���ܳ=��uxxX=����>&��\&���ؘ�����OZ�ϟ�o��3g�(���c�e  �HWS  �^'���!,���t��ꡇҞ={L�A�޽[�>��>��O�̙3z�7t��yEQ���I[�=�����׮VcH�L>��H�N��?�PLݟK�vx�\le�������~�k�h��i��Wo���V��	|��?����2�� 6���)'����lP��~׏w��=���:p��2�װ��y�����Ą��N�:��^{M��Ӧ����q   X�  H���;��ٳ:�������n1<;;�7�xCo����]*p��H�ىT�O �o�$j�Z:����ǻ^ �&��J1�]����t�?���� �53���}OS�����
�'Oj��1� �T~�L��Rݺ~;<<���_>��v6����z�!=��C����/�K����j�ۦ�a�J�n�  ��jJ   ����}A��������5<<l:��O?�'�|R�O����s]�|yGǴ��n���,t"����j�}3�5 i�e����5���?ԛ�����U ��������=�<��o|C�O~�t4 @�d|_�BA�ެY�{��u7��t��w�ĉ�b*�ў={���~VO=���x����kZ\\4�W�tD�{��   �,]M	   {��a
�J%=���:~�8�yp��V��ONN��^�;Ｃ0���[�LpҫV��l��y=މ����~�/�EO_���f_}U����ܮ]|�UyDC�>�<�5 ��b��?IӶ�����n�\N<��>��Oj``���f�BA'O�ԉ't��i���?�իWM���w   ��Ք   ��=�`�u��q=����+#~{���/���{L�����x��Z�M�|���}_�|~S��T�=N�\�&o �liiI.\����)��J��?���Y?�g��g��3ͩ)M�ٟi���L��w�F�W����J�� LɖJ
ff�6$f�(��u7��`+n�r��%��'?�|�(�LG��}R�wL�   pYz�   �: i�tll���:y�&&&(�a�*��>����G�믿��^{M�ZmßKS�}+�{�/�މ�"(,�����/ꮻ���EX���zr�����G��+�Ʈ. �X|�m�~�m}�/���|�K�C�]�L� �,(����+�o��U�m���ȈN�<�{�W��Ő
���/����)���?ջﾻ��>�M   p]z�   �:a: �l߾}z�'4>>n:
,P,��c��ĉ��/~����j4�>?M��&�w,_ ��	���.]����1J�J/&����?���?P��t�� z������G����j�k_Ӂ_�u�c b���Krm?����o�wx�?00�GyD<� �vtŮ]��/|AO<�~����7ߤ�l�L   p]z�   ���� Xۮ]��裏��ѣ���B�lV'O���?��_}ݢ��ڒ����xLp�e��������O���x�2A��ݝ�������D��@X��¿������#��[���K�# b�LpwMd�|����X�}�Q��虁�}����'?�I��G?�{ｧ(�L���I�KZ:   z��;  �y���[������=��CQ=���t��I=���z������L�fs��k-�%Ua�����;a�;l����?�P�  kd�ٮ�O}�;�����"&�Vi����o~S������{�i� `9�XTV�'ɥwu�(�y�D__�N�<��z(U��^���������)���ݓ������M  pw   ���0!*���z�)��0�P(�����?�W_}U�����0T��-��m)���w�wتZ������a/�U�ÿ����ٻ��8����OU7@c%A�$���H��(J�$j�D��,ْ'V<��ؙ$g�8v$'���M�Q6*���ڞ��3�=�NNb'�8�sm�VdǋƖ-J�@�;[�F7����H���4��~����spD��>�����~��?��SEJ��z����ڿ_�>�	�o�� *U4�#�J�囯��hT��պ馛�m�6��b��z��t��}�;���ӧmG�w   k�є   �\��5�C�]UU����z�p�\Āu�x\w�y��mۦ�|�;WL��Lo�4��`�E(������K������sc�Y?����ɟh��?_�D �j��i����?�#Ϳ��q  %��%���n�y�\NN@�Ö́1FMMM��_��/��lZ�d�}�Quuu�[������lG���v   �0c�  �]k%��V��hӦM��>�]�vQă�̛7O�x�;t��)��^]]=�Ǉy�{���v��FGGu��1e�Y�Q�9�m�'���{����ہ�ɧ�z�7S}����( �p/������)�TJ����ZZZ(��w�����Oh��݊���k�f�   �;  �]�l�ŋ��Gս���E����^}�U?~\����Lj��+��h�\&�#�٬�;�t:m;
0k���>64�o}��:���W	�;/�ӫ��[��mG Y��	�aSI��������K�x��F�s�N=��ڲe�Ǳ)���   fQ�   B��eV__��o�]�ׯ�(�1F===���W[[�.\h;�[̸�^AGg��;�"������jkkScc��8��ʹ�>|������h���%^6�W?�qm��C5mm��  ����*I�$c5MyUc�N�>���ny�g;P���z�}��ڸq���o����v��Y.�FR�  �  ��v��pG�6m��?N��5>>��Ǐ�������b4U4:���+i��LE.\���S�N����v`ƜhTr;}z��W�����r; IR��O���o��x& ��\<�w�	rAR�J���~�={�r;���M�}�{u�w��*�{IX�J�`;  @XQp  ���u477�]�z����O��hxxX���שS�d���a��w����_nLpG����̙3����D!S�_�����}������!��H�߯����ڎ (�H]ݥ_�l���ꐂ���<x�W�"��r]W۷o��?�+V؎&[m   ���`  �7kl�d��jǎ����Dl�����g�jppP+W�T�eZ˭��zfO0�"���-&�#���d�l�2��!0�Xlқ��|^/�ٟi�_���� &p���½{_��v �]~�zL҈�(e��a�t��	e�Y�Q��kjj�#�<��^{M��/�����v   ��b�;  �=K$5�Q�Z[[����G�w�܎�6::�����ֶY���|&�"��ʉr�9�+����ѣ	SA6��L����k��?ڟi ���r�ڷ�v @D/,��uM�
�\NG�ё#G(���9���7�}�{�֬a�R�m�    �(�  �ö�%ຮv�ڥ���=jmm�(c�zzz��+�hxx���ϸ�Э��!2ÿ+�]�&���� �r&(��߿_���:���[H h���]���� �9�|7��܃2����_��������(@����顇�<0�]6Q���   �w   {��Pi�s?��h�    IDAT�sڵk�\����l6���̙3e[3�(6�t�ɘo��^vA���n�:uJ�|�v`R�Op7���������?h��?k߉?�s�  s���o�ZR��f�|~��'N���K���� V�_�^�=�����lG�D��&  ��0{  ��ѦM�t�wθhTc�N�>���A�^���{f:�]b�;�7ittTmmm�_V��b�=�߯{�i����-'D����F_]�+Wڎ ���U7��$��J��{:��ѣG��qF�\. z饗��/��<ۑ*E��U��X�  :��  ��m� �����׽��K����Ȉ��߯�����3�}��.w�-r��^�uuww�c;p'Q�O~�������̞1:��/�N ���
�aፍَ��uww����ہ˸���;w��GUss��8���  ,��  `�Z��n���z�'�a��Q _�<OG��ѣGK6��	�3s�q o:���;�l6k;
 ������O5��c;������$n����\��T��6������t��A�8q�	��$/^�����\;)�km   ��� (�O��K{{{c��Ǘ8�s���3,I�H$��  ��^}�պ�~���l�*�q�}�v�v�mr]�����ק���Y�F�E.X3�}f��L-����ѣZ�h��`U&���ӧ566��+4��K�#��s�4�ӟ�q�V�Q  ��D�rc1yn�S�=�	�TJ]]]�𽋻�.[�L���7�!djkkw���A��  T*�q���|��u��ncL.�N���d?����Pp��|�3���������ht��yˍ1K�i�Ԩ7vȫr'b�qFFF.Z�1�n��I  J���0��bڳg�֯_o;
(cccz�״j�*͛7�h���|Sn�GFˍ�;0=��t��jɒ%��>̖1F���:����f��V��b���w 0���R�=r�#o5Qyx>�e���['O����6��mٲE---��W�����q������|���s  �߿دQ2���8�������4d�9�8��uO����D"?�����?��tY� (*
��L&WJz��ݒ6KZ�8Nc*���$�u/�q�8�[�ρ>  �r��9�i޼yz�����b;
H�穫�K���Z�lل�3��f���߶�.�78K������5��9���N�u��Y�]�s*N�@����jկ��� �Y���|��
I�����t��1���[�Y[[�{�1}��_Չ'l�	����ێ   .c�q��!YTR��&�q�K��y�\ו1F�TJ���9c̐���^�􂤿��'_��@�(��Ѕ2�c��q��Ƙ����� @p���؎8���ڻw����mG���[���jooW4:�����{���P�uwwkhhH�/f�D>�Woo����&�z|��2'P���Xw��[[mG ̂{��H��0��y'�ɨ��K����2 �"��Gы/���������Ȉ��Ƹ> @ c�$�\��,�QI�uvv�c�$��uIE��(��@2���u�_�<�m�VH��]1Ev  *Ooo����8�n���ܹ�ɭ@�R)���Z�f�����^#���ya.��55�# ���d���k���Z�`��v� &288���n���O���%K�VW����"1F�/���?l;	 `"W�?������&���ѣ�v10w��j���jii�?��?+��>sg�Qoo��.]j;
  (��[/|�)����䘤��~���>��?��ܭ���?�4�N��1�~I�$�80  \�ΰ0�HD{������mG*R6�Ձ�j�*͛7o�ϯ�eY;�A&��g�����500�h޼y���Y�d2:w������u\W�+Vh�С2$P����_)�@@]]p˅v�͖}���n�<y�Ap@�lܸQ����������!�={��;  ��Z�:���I��d2��t�q�����?�Ї>t�r��	�q�u����H��1枑��E��   ����mG���Z=��Cjkk��h�穫�KmmmZ�dɌ�;�	�&�A�	�����y�;wN���Z�hѬw�@8������G3z^|�*
� �����M^6+w�� �\}�:�K�ĉ���.�@-Y�D?��?�/}�K�����zzzlG   �����ydd�����!c̿������Ǿf;\Pp/�g�}vw.��ϒn7�0�  HzcZ$1���ܬ�~X��Ͷ� �q��i�r9-_����ȳ-��y��K�(�L&��_]���jmmUUUX�%�����ק���k6;)�W�.A* a�O�5������lG ����#�\I��Ow���x���G���fT ���ԤG}T_��u��I�q|����v  `�1�Q����ݟL&G%}�����>򑏼`;[���^d�>���l��v�\.�`;  �s�α�������C�����r�����ؘ֬Y#�u�|l,��1���<���m@�)�J���I,��+c400���^�����ujW�*^( �7��Pp� r'8���T��{٬d�T�@����r:|�0�a jjj��#���_��^{�5�q|��;  �J����\no2�Lc���~�#���l�$܋ �HD������p.�[V�C  Nl�:�M�6iϞ=�.�����!8p@k׮��$:��������ࠚ���p�BE���
3c������۫l6;�ף����C�  ��j������ƹ�R���d2:t�PQ޷��H$��{����Y����l�񥾾>�  �58��\.��d2�'������G"��Է"�J�ttt�$��u�[�1�y  @0Pp��Ν;u뭷�����^{�5�_�^���>f����;�R�XtRss�ZZZ(���1F�TJ===E-��W��\W򼢽&��J���##���َ ���$�0�g2%9��N�u�С9��8�Ѯ]�����o~�����N�5::���  `:�%}�����;::^���SO=�o�C�1g�����d2y�q��9�s�v  0lc�V;w���ݻ)�>��fu�����N�u
�C�(����ק#G��ܹs��r�#��<�S����t�ԩ�Otc1մ��5����5��ێ ������r;m)��R)8p�r;�3[�nս���N�`�  (�1&�8�m��|/�L���'?�qۙ�(,��s�H$j:<����8�U  ��6�orG��v�v��a;
�	�r98p@�ׯW��)es)��3�ݍ-��.����T__�0i������_������%]+�z�2'O�t �1��j���ڎ ��0Op/v�}hhHG���I�/mܸQ�HD����ȿ��twwk�ʕ�c  ��Y��':::�/�u�<�J=�H$�{�|(�O�3��L|dd����o��1U  ��������8���m߾�v S���:x�֭[���7����b�~�0Op�0��fxxX��Ê��jiiQ]]����ؘ���488X�m��W��;�)�Z *��~`; `�&*�G�Ɩ�^��8�```@G��4������F���|��7�����mG   �8N�1������cGG�?����b"��@4
�H$�����~���  (�\.�t:m;�u��jϞ=ڴi��( 
p��v�Z544���jN[Ԇ��>�v� �+�N+�N+����I���SUUX�.�1F�TJ)����V�}M �k��A���	˒  ��{v��J?�Q�s9���:z�h�nR07���z�G�����f���X��  �ǉJz����d2�w��ÿB�}b�o$T�D"M&�����z$��r;  (����П�w]W��?�v `<���Ç5444���Rq�~�[]m;����u��y>|XǏ���P�ߧ���ؘ���u��!�:u�J�]zc�; ��)��+�S  f R[;��˜Æ|�����Rnhٲez���|N�Pp  �t�������������H$��v
���'?��������^�K  ��z{{mG��u]�ݻW�֭��,x��#G�̹X�xڏ˅ ��FFFt��)>|X===�N~�����߯cǎ���K�ϟ��%:w �6�ӟڎ  �w�	�a��l�x.���OǏ��T[[�~�������o;  �Lc�������dr�1�^��EHJ&����ٙr]���  �L���讻�҆lG0����ѣ��.iŘ�T�Woo�������Eٽ����u��	:tHgϞ����X�D��U��j;�
��� ����2r
�sVp��U��@����顇R$�}+&�J���|  *ZL�G���7�L&�v?u���g����ٹ_��1���  ����o��6]{�c (�q�ӟ�T�TjV���\p���@���Ʈ(����Rv/��K�O����o�/�۷ێ ��������w ����>�YQn*Ȋ+���u�Y5�<oN�_   
q�������7��cS(�u&��d2�e��^2�l��  �GX�/���[�c��1 I4U>��O~������(Z	��o���ؘzzz��եÇ�̙3��y���1F�LF�ϟ����Qj�\�Ν�# � ッ=y�v @��<�=?�	�TJG��	�0k֬�=��#�qlG�����v  ��,s]���d�ˉD"��CWp��������^Io7Ƅ�7  �&���n�I7�p�� ���6����z�嗕N�~��	�6�N4*'�Ӎ�J���400�S�N����:~��Ο?�L&����\N���:}��:��G����[###��;��k�ҋ� J#�ӟڎ  (�d�#����f��
FFFt��a��@�ڸq����ʒ;w  PN:�o���������y�-7�K��Ă���0�첝  �����e�c��|�Ͷc (�H$r���lV/������:UOr��ra����b�# (2c�FFF422"Ir]W555���U<Wmm�����l6�t:���Qe2�U����65lެ��~f;
�
���O����c  
0Y�]z���g��������Q:t�r;P�6oެ��Q������U__��   ���y����W\׽����ہʡ�o&�$uvv�NCC���  ����!eg��kP�[�N��v�� �,}�}ҙLF/�����ǧ}~���   �<�S:�����u�ĉK��Ϟ=���~��i�+hc����488���n?~\TWW�Ξ=�����*�_�z���# � ï�f; �@N,6�n>�>U�+�v.���Ç+���v�ܩm۶َQV� �MƘ��������Yʡ������7��cL��Q  _
Ӷ��-�޽{C�=%P�&�D<22����gںu�ޯ��dJ����*� ��1F�LF����UUU�����GUU�b�؄7�A>�W.�S.�S6���ؘ2���٬�1����{���g�-�� S9|X���L� ���ʭ���}�?��O!<���ÇC5��t�w(�J����v����  l3�D%��d2�����[~�����L�R���������y��$��  ���^MMMz�;��ۂ���������<�k��f�Ǆy�{���v >q�,><<|���QUU��hT�H�-Ÿ�0��O�q1���/^�j�<�>������ڎ��GG�9yR�+V؎ (�����^@i��ѣJ��eH�O\��<������ٳgm�)����   .j<�L&?��O���0�Pq���?�|������yޝ��   \����#�\MM�~�a��q�Q ��t7��={V���Z�r�_��� �2�(��4��u]��{��~q��q.�a���y�ޘ�xqں�y���h�����(s�� �"}�0w ��Z��FU�/�_��rS~�ĉ�>��F�z衇����J�R����訲٬b1fm  _�J��d2��+V�}��G+jK�����S���5Ǐ?-�N�Y   �V�'�]�����v͛7�v %TU@I��ѣ:wn��
��U�"�ն# � ��i||�Ҕ�L&�L&���Q���hddD�t����,ً�v�
-ܻ�v b��a�  r'ٝ���S��w��Yuww�1 ?����#�<������  �jw?~��3�<��v�b���{2��p6�����Y   &288h;B�8���{�j��嶣 (����s���	o��h�s�� eՇ?�Hm�� *�ȡC�#  
�NR܌��.�O�L2����_�N�*s ~5�|���o���\�
Î�   ������:;;�v�b	��Jc��L&�&�9cLaM   *��s�Nmذ�v %�n�'<�����5vU�ݛfK�J�Rp��R�ڪe�{�� *�0w ��$ܥ7J�*?A�}ttTǎ+ ��b�
�޽�v�����  `2�1插��׌1����H$����aI���  0���!�JbŊ���m� P�No�(���g?��<ϻ��0Op�� �g��߯�u�l� p�S��� P��vg���������9r�9 �hǎZ�~��%3�Υ   >sOgg������E`��d�������㬶�  `:�lV�L�v��khh�}��W��Mx�LJ�t貉��$[Z��T� ���b������ ̍19r�v
 @���I�-c�r��|�믿��]� �r{��QKK��%���o;  @!�9�����>��u�DJ&��*����lg  (DOO��E�D���*�ێ�LfSp��3g��̙3�$��3R�D(?@E���k��O�c ��ÇmG   RS3��y�@���w��ʝ �����C)V��D��  �&���˅�u��8;�L~Rҟ*�� @x���َPtw�u�-Zd;�2�m�]�:�T*�w @EZ��cZ��wَ �2'Oڎ  (@�'��R)�>}�r A��ܬ��O��؎RT����#   ̄+�O;;;?e;�L�8����o%=b;  �LU�D��[�j��Ͷc (�ht������W^Q[>_�D��Rp�����W��	����`���r�QE���,4��x��rE�q9Ѩ��jE&(�9��܉v�2F���|:�N��a٬򙌼�Qy���������-ҟ~G� �a���������);6���.�Q L{{�n��}��߷�h���d����>  �lƘ_K&�k�|��lg)T 
��7�L~�q�;lg  ��Jڮ���Uw���2 ��2�]�2���64H�#S�T�A� *��jSg�^��G5��َS��U��AU����mlT�����^�pkk��q��'*�������f�O����������S�7>�����������0��

� a��.�Ց#G4~ٍz P�]�v����:Y!�y=�S*�R��  ������R���D��x�?�N$5����:���v  �٪�	�HD{��s�@0��~��Vέ��}�"$

� P�"�}�9���S�{�E�qǭ�Vռy�-X��y�T5o��,P�¯c--�͟��y�mn�㺶#��[S#����t�3�R�}|p�ү�}}���eϟW��W�CC��� �R��J�	��[�fg �亮��>��_��2���8E���K�  �1f[}}��D"�1�H��͙��D�����5IKmg  ���
)�q�jii��%ź��<��̑#rΜ)���C� B������N��?��/|�v_pkjT�d�b���Y�HՋ�QboiQ�BY=�`A`&���\�a�^6�lo�r�����)�ݭl_��Ν�عs�vw+s挼���|:�\���  vLUpw�F�=_�4e�t�̎�S ���z�}����W�b;JQ�������v  ��ZU__,�H\�H$l���o��=�\c6�= i��,   sU	�U�Vi˖-�c ��u]9�S��F�=��"�>+�r�y� �Lq PYܪ*�y�)5nۦC��{ʧӶ#��[U�Xk��/׫-z����g=yV���j��T��6����9wNcgϾY|?}Z�S��9uJ�
�ɬ�FO��� >�����*��^]-s�}RHv�PZ�֭ӦM���~�Q�l`��=0 ϟ4�    IDAT �B-jhh8�o߾k>�����3_�;::Z��쫒���  P###�#�I<׽��[�r+��)���K/�y�9_�Rq_�ǜ�*�  e���{հe��tt���߶gvG��f�R�,[v��,Q��E�8!��MM�ojR���~=�Nk��IeN��Tz��1v挼��X�̩Sj��r �&�Ko\|���p��el� PA��N�>}:��Jl  `�Yh�9��ѱ񩧞궝�j�+�'�z�uf���  *B:�V6��c���=�ܣx<n;
 ����>z�w�=xPΫ����h��� ��T�d�6�ۧ�o[G�{N�c�lGz'U�ҥ�]���{�e�Y�Ln,f;"(��~����̹so��/�އT�/�?����:e; `��y<�]�7�Lr# �V,���߯/|��<�v�Y�  �X�;��j"�X�H$|u��
���g�T�1f��,   ���mٷmۦիWێ���Op�$Ǒ��w+�o�4<\���ʁ n�o�]�v�V�/���oJ��J�3D�(�/]���v���U�t��k��s
�庪Y�D5K�H;wJ��lV߽�.y���p�d(���9Ӽg�����hj�w��S �P�-ҍ7ި�}�{���Z*��  ������~������7[�����矏����:���v  �b
����F�z뭶c ����%��Q�;�)����4��# ������r��J�߯��G���?){�|Q׉-X�x{��֮U��]�ի_�JѦ������������ڎb��ɓ�#  ������e�QR�#s���1 �Ѝ7ި��.uwwێ2+� @j�f�'��b
�/
��7�L��8�
�Y   �-���ў={TUUe;
 (Y�]���:��X��I��4ݔ7 @�4lڤ�M������4��K�я4r���Ξ�)`��؂�]��2{�ڵ�66��O _�M7Qp �Z
�f�f�\�PZ��������y��w  P������c�:�c�M�/
�������8�m�   (��!���3#�6m�
.d ��uݒ���w�NΑ#R�7��D���v ����7nT�ƍZ��c�$/�U��Ie{{�e2�g22��HM�"���SͲe���ZW�֭�#X���<O*�{o ��Mw�z࿃���m��N $-Z��۷륗^�e����5::�Z�� @�qgugg狒v��b���L&�_c̍�s   �����3��u��ێ�GJ9�]�Lc������/�t��� (��)�ޮx{��(@Yխ_�F�;������Sl��I  �p��y=���]w�p�>�2��[t�ȑ@^K��  *�M��SO��f�7�wvv���o3  @�q�����6Us!�eJ=�]�̭�ʬ��ͽ"�  ����(�j��Ve{{mG  La���+�)O��ko�Y��v
 !�F�g�9N�{���ێ   P2��<�L&�63X+�wvv��1����>  @��R)�fd���Z�n�� |�w9�̣�JQ뛍��SUe;  ��}�
� �o���icu��l�b���v
 !�|�rmܸ�v��  ��~����m-n����g��n�����  �-H�X,����v >�n�&蘅e*��tS�    �,]j;�U���
9�b���v�T_o;�������mǘ���A�   J��?��?����e?�N$����/H��{m  �r3�(�NێQ�]�v�� �R�����KZ���k���َ   �{��mG  L���{�.����\{�� B���F�v�cF(� ��pc�ط�D�/����^__��ǩ+��   6�R)y�g;FA����m�6�1 �P$R�K�Ѩ�(�e�Pp  �Vu[��V�lG  L�'��;�ʴs Le˖-jmm��`��ö#   ��1&^WW���1e=�-�b���_����k  ���w�qG�K� ����u�̚5e_��"\  �XK��V�َ  �B�Mp_�^&仧 ��qt��ێQ0
�   L�Y�o߾�+�e+��۷�Ƙw�k=   ?
ȅ�+V����v >�vf�y�|�di�R`�;  ����Ϸ�*&�������i�U����۽�v
 �²e˴v�Z�1
222b;  @YcޑL&�c��+KS�駟^���?[��   �$�Jَ0-�u5@�Y�ݡ�M�7�Y�\
�   Ӫjn��8Xɘ� �7��A�)f��^jl� ����oĎ�� @H�Igg��r,T��kc�[[[���8�R�  �7A��u�V-X��v >fk��$���jj��_4�+' e   ls"E�q�1��� ��VWO��@������i; L���Q;v�cZ�lV�\�v  �r�Hz!�H��^�¾}��$iq��  ���a��TSS�]�vَ��N˩���g�������   �s+��Y�ڎ  ��t� Lp7��*UUَ ���TWWg;ƴ�0�
  �،1������z߾}�4�<X�5   �,�Jَ0��;w�&�� ��9�]��m�I��[�0Wn�M�   
5]q�����< @�}�{K��5��N S��b���mǘw  VƘ;;;�]�5J�Rx��=���R�>  @���؎0�x<��[�ڎ  l���{���f�+�S�  &�wy��l�v
 ��inb��ws�-��؎ �ڲe�mǘw  fƘ��H$�K��%;���$Ɓ �P�s���nP,�@ X/�K27�(��؎1kLp  (\$�;�y���#  ��VUM�u�/��ʴ��N q]��S����3  @�U744|�T/^��B2����8ח�  �į���:mٲ�v ��a�W$"o��)fm��n   xS�'�K�Sp _+������y7���v ��i�&555َ1)&� ��3��L&�.�k�����k��Q��  c�����馛�l	� �����.�\���j;ƬPp  (w
� �kA-�/Z$�Ze; ̈뺺馛lǘ�  $I�D"�\�-��u6����p�}  ���=ϳ�-�y�f�1 ���蒬�ʻ��)f��;  @�(�Sp ?s���Lr̔��V���k��F��ϷcB~��  ��buuu_.������g�y��[���   A�ש�v�R$�@@���.�l�.�d��3��}  �`N��J�Qp _+���y[�̊�S �����]�vَ1���a�   |�q�[���/�k���H$����Q��  :?��q�F�1 ��
�r��ﶝbƘ�  P8'��e�\�v �
9�����C�P�֭Ӽy�l�x�QnN  ���D"Q��E;�nhh�s�q��z   A��m	���:��U���Ef�V���1f��;  ���=h9��q�  S(d�����.X �|�� 0'��hǎ�c�w  �79�SWWW�ߋ�zE9�~��Wc�[��  �~ۖ0�i��Ͷc _��2�w�N1#�  f �wy�� �)m��ٹ��� *¦M���mǸB:��1�v   �p]��~z]Q^�/����X�  P)�6�}�֭��b�c _�%��n���Ō���  
��]�ʉ	� �o�*���ˬ_o; E$�֭[mǸ��y�f��c   ��1Ʃ��y��5�c뎎���1ۊ  ����i�.q]W۶������XLf�.�)
�w  �y�ݣ� ��VUM���$3�]'��� �����UU���r�ێ�   �9���������u�|4�8���k   T"?Mp��k���`;� ���Ls�mR@��Lp  ��-��ێ  �JP&��b2�^k; UMM�6n�h;�R���   ��D>=�טӱugg�KZ0�   ��Oܯ��:� �o'�KRC��Ȃ ��    8B^p���N  �B!�}q6��k��j�) �访�z_��f�;  ��tvv>9���;>c�����   �ltt�vIҊ+�p�B�1 ��.L��qG 
PLp  @��� ��	�wו�}�� PMMMZ�z����iGg   ?1�$�1�>D��;;;;$����   ��/ܷm�f;� s|^�1�ˬZe;ƴ
��  �7�\�v�x� �V��i�gSV��m� ��ٲe���0�  `Ru���4�'Ϫ�����ǌ1�>�E  � ��؎�x<�) ���wI27�d;´()  ��fmG����.J vnUմ��}6�\{�� PZ+W�T�On����+   �����?��gu��ĉ��f�   @c|Qp߼y�\.��� |1۶���ڎ1%
�   �{�]��� �)�~�{]] v���pG�7o�C�422b;  ��Ŏ;���g�T0Ƹ����l  �t:-��f���= ��	�v찝bJ�  
gr9��r(������n6o�0�  ��/C���  05�u%�H�������%��?p�f��  ?��Z�l����m� p�(�K2�vَ0%JJ   ��w��#��ܪ�ic�l��H=���Z�r�����  ����럞�f\pw��f�  ���C�}˖-�# � �)�/Y"�|���b�;  @ἰOp�# �Z�w+gT�/�ij��2 Xq��ڎ@�  �01�̨�>������E  !�����Y��j (7s�M�#L�)�   �3!/��5l� ~V�H6
' Bf��ժ��[c��  P�ڎ��'g򄙵�]�7g�   �FGG���q�FE"� T��Lp�$s�uR,f;Ƅ��	  P8/���*
� �s~-����0�@ȸ���7Z�066fu}  ��p]�c3z|���'>q���'  !��6X]@ep'PwUW�X��1)n:  (X�'�GjkmG  L���*�qe?��n���h� T����[]��5A  � Y����@�.�7�t�.  @��<���РE�Y[@�T���m��r��  P���a���� �V�.m�>�b֭+� �����?���=�S.�7�  ��>���{2�\)��Y'  ��6��
�����l�$��؎�VLp  (��<�C^pw��~ pI���:K=�Y���+���]�����t���   ��B'}Z�Ww��.j   Ae��n{+F �#�wE�27�N�Lp  (L>���<�1�b�; ��/'��]+�e����lذ����  
�H�d!,�(���g  �L&ceݦ�&-\���� *O ����#�E��  �.74d;�UnM�v� _+t�{9Ϫx=r---�?���m�  �w�i��d�$1.  `l�7l��B* �	���a�TSc;�(�  f|p�v����mG  L�w��q���\��o���	�   3R��3ϼo�2���E  *cccV�]�n��uT�����\{��W��  P�w�  �(t�{٬_/��n� �kÆ�֦�  03�|���{̔G����/ic�  ���	����Z�pa�� ?2[�ڎp
�   �a�;w �;�Mp7kזi% �y��i���V���.  @�m��Q�Ԕ�|>�;*��i   �"�͖}�U�V�}M �-��u�⮏J宏�   ���А�VE��lG  L�O����L[�� �����|  p��y�y�LYpw�狛   (��e��L{���8���   ����n; `nUUA�+�؀+$w�K� *���ٸ.  P��Oz���Oz��%E�  �\���E"-[���k�ߙlG�����  �n���v�b�Ͷ#  �Qh��,z WX�l�b�X��+��   �-�L��싓�GFF�Ki�   T6cL��˗/W��$�"s���+s�5�#\⫋�   >6��m;�UQ
� �{~��ݬ��  �亮��P�  f�q�ߙ�k���y�4q   *[&��1��k��r |m�"i�<�)���N   ٞ����� �Wh���cZZdJ�
 ��kf�  f��}a��>��EƘ���  P�l�Ģ� ��w�G��   �l���� �i�e�6�9a ���kf���  �Rc>��3K&�ڄ����'K	  �r����u���F5s &d6l�A���/  �-�S��y�)��� ��c|
� 0���F�+�ΞLp  ��|>�щ>?a���Hi�   T�l6[�����T��i��Y�Nr'<�-+�\�  ��^��lǰ*��d; `N��KzV%�Y���+ @��\����1�  `N&쬿�*"��cV�>  @e�d2e]oٲee] ��Z��_��  �.��k;�uU���\?�ľx1� `
mmme]�	�   s�����Ǯ��[�z�p��a  �Y*w�}ɒ%e] ���`�7�  ���==�#X�����؎ ����e.n@�,-�Гr��  Pa�'N<��O^�	c�{ʓ  �2�sJC}}�ʶ�pq��n�]6~(��    ���E�lG  ���{)Ϫ
� 0���:566�m�\.W��   *��y?��&:��Y�,   ���ro� \*����n;�?Lw  𹱳gmG����  0
9�/�YǑY��T� ����r���a�	  �l9����GމD�YҼ�%  �@�܆��; ��Af�|�(�  L/s��VUSV���z�?�TSco} �r^C�<O���e[  ��߷o���8�nhh����  �<���V���~�L�  (���-� P '��1%��ti�^ *J������   @%�<�������1���  �<��PUU��e- �TI[��U����  0��ٳ�#X�� �aq��Y���� $---��be[/�˕m-  �
���s����2  �H�:��x�b�6��P�*��.�w�[�  ���)��k;�UՋێ  (��	��� ��hI�gRp  ��+:엮�c\I��  ��VkkkY��J`-��Q�1   0��s2�g;�U5� 0�����4����y�g~�_���g8�C%Q�J�(y�^�k;~�N$@�dÈ8FbA ���ȉ8�"F� ��I��țc�s���]kq��cuߢ$��x��9���]��!Q��ǐ쪧����%9�~�$�ͮ���{6�Y������������� �FY�m���?��M��������?�L �JUܯ��J�h�N'��Ү ��J!�,���#Y�}۶��-}��ڶm[ek�� pu�������ƹ���=�f�H  �2*Y�ʩ�x*���N�Hx�w��  1���֭��vS� `��q�_ʮJ�EM�6���n�; ��˲��.��~���� h�*
�N'�n�Z�: mR\�c� ����c�����o_�8��G���pe%u4(]������<m�˖ML$Y�Pp�,[�n�N�y�����; �H��|��~Kۦ� �P��[�l��D7Q kǎtk;>���WW�䣏Ɖݻ�����#�#��\}� \�Tw�.Ϲ�Qǎ+}�*� ��[��`2"�(������̧� �ULp��HE`|��!��������r �ǙW^��_�b�s��18s&u����e��#�Uɲ(��fԯ
�z۶m���n�; ��˲l�(�N�e�dD�����~6�I�  �Pńw�+0?�qcD�"af�; �������~�|��Q������ �Id������~]���Ꞛ	�  W�(��?�����F��'#"��_O�	 �5Lp���"{����Upk��c���N���Q������� �I
������; @��ÿ�
��a  ڤ���[���@Q��0���o�HPpOr���<���ś��{���������7�� ��X�u��wU6o�+��-[�T���; �hLLL�?�
�H� �U�</��;�N��ϗ�@[[�D�Y�	� c���;��o�F�z��Q���t�1}���c p���K~���6������|t:����U��#m    IDATq�3 �8(�ⶈ�
�EQ�9 ��pX�����E�$`�+��w��r���_���;�:
� 37�����I�],,T�&@t:��������R�)��  ��>"�ܕ��  #R��M&� )��,	w Jv��ߎg~�W�ہu�p�-�# p�RLpWp�r���r?  ��("":����7�{�� �zeOh�b���Dw9�ño~3^��"����Q�Qph�u<�>�{̛Yp��e�; �hdY6���~cgÆ?�: @��=�A��JQ��Vlz��33կk�;@�߽;^���2�� u�afo�5u .W���وnw��0V����� 0:6l��N�e?�: @����E+�Ql�R��&����={�_�u�v��̘��J#�U�'pU���V� , �q211qO'˲;S h���
�@U�Zp��[�_�w��Z;u*��G�(��˩� �A��q�� ��;@}lڴ��5Lp �;;��K ��
�@k(���������GS� jbn.��\�: �i=;&#�U������
�G� F�(�[;�N��A  ڢ�ͫ����� �x���ƒ{�qc���c� �s����8����c 6��O�� ���qR�HwT�	\�*�)� �N�e;:EQ] 0"����ן������R� ��6�S�^��� 4�`q1�����:�pswޙ: %�J133�W?U�_Sp ����H0� ���޼ڰaC���Q�,��ͥN @���S��:�:�p�wܑ: W`=��tGž0�U�)�a!w ����D�ǽ F��ͫ�7� >J�}4Lph�ށq�K_Jh�ک���\���H)� �ԆNDL�N �&�m�Ƃ{1;[��
� �����Q�q��	� �e���wS�\����y^�� ���NDtS�  h����&�Ukc�=�w �c���x�k_Kh��֭�ݺ5u �D��¾0�Us� �Q�:Y�# 0"eAMp��ڂ�%nD�Zf�;@k���"_[Kh��;�L���t7%�"��p��.��r/  �,�&:EQT{W ��Lpڦ���݊3��P@y�K�# -1w��# p�.� �HwS��#<8p��"�ʽt �D���:Y�.; ����y5mRP�<�SG(G�'b��h�Ճc���S� ZbV���F��R�C� -U�=6w ���Lp ������>�G���^T�~��r�v8��C�# -2w睩# p�.q�?Ҋ�=a���|��; �He�2 ��7�܁��vS~r�����w��8��#�# -�ML��Ν�c p�.q�?�q��F��{l��K HD� `��޼*{��G�u�{Vu���+�Xz��)�����'�3=�: %Qp�w �fѐ ��7�&�,dD{7�
og
� ����[�v�d�@Kl���� �
���Wp�w �fQp !܁���#����2�� ����3�# -2�kW� \w��)���; �h�� � eO� ���n�Wy"�	� ���쳩# -b�;@�]j��HwS<80&� 4K�, ��)����;P�<�̱����T��܁�ɲ�۹3u
 Jd�;@�L�<�D�
 `�:�z� ��+{���>��w�����Xٷ/u�%6�|sLnܘ: W���~��;@��� �,R   \Pk� p���%&���x�=�# p�*-�+L�D�tF F�(
w �Q*{�J��Zk��խ���μ�b�@���# p����_�N�}��^� ��Ȳ,:�-+  $Pv���P��(�Yr����� c��K/�� ��§>�: W���#��W��>@��}��w ��2� `�܁6j���n� cfI��lr2�v�J��t�	�#�	h�@
�  ��� �9ZY2j���*�޻m�ĉ�=�:�sw�����1 �Z���c�wCO FB� �Y:Y����  �FٛW��	����?S #K/��:�"��d� ���f�c�-ܗH��!R
�  #UtZ9�  �N�S������������B����^z)u�E��A��y�"�� 0Z�  ���S���k�{O�'b(�4֙�_Nh��O:u F�"��q_ ������  F�w �*{�{+K�@�q�{V����&�Pog_y%u�%fv��ޚ: #`�;@�(� 4K�, �1S�����j��p>�|�fe�����i���G����Ė�~6u F�b��#�E�'0e�cSp -w �*{�j��B&@D'���vz@#�}�5����l��=u F��	���)� #P�=6w ��Rp ��7�z�^��p>m���-/W��r$@#�}�����ޱ#>���1 ��"{%e�d����!R  ͢� 0B�N��܁Z7����ʗ���� ���믧� �Ď_����"���P(e\5� �E� `�&&&J}}�%��6��HPp7�����ٓ:���6����c 0By��þ0�U+{�T�� ƍ�; �)�mTE-*hg)&���!��P��wo�@��w�nL�Φ��eOpϜ�	p�� �E� `�܁�j�����	 h�ޡC18s&u�᦯�>n�;'u F�B܋0�����Pp hw ����,����a��������y���H2��E �b���SG Z���O�33�: �v�	�]���pU��~�{ܝ�
 �(�t 0Be�#Lq�h�ww �ᬂ;p���sq�_�K�c P���$e�dN��*����� 0Z
�  #�eYdYV������>���i�{�8Q����@}��ۗ:�`37�w���: e��>Ii�'���J��� FK� `��>�P�H�U�S��� ��Xy����������ߊ����Q (ɅNj+m�Ğ0�U9}�t�k�} `��t 0beOhPpRhS�=;y��EMph��7�Lh�lb"��w�.�v�L�2)�4�	�  ͣ� 0b&�mԖ�{����U�n���(k�NŠ��n@�t:q�o�Fl��gS'�d�Op��#K���
�  ͣ� 0beo`Uq�"�G��F�8~<ͺ-y@ `\��z+u�a��ɸ�������ϥ�@.Tp/u����+�� �<
�  #�eY��o�;�Bk&��<�f�$�p���ۗ:� ����ݸ�����Q �J��#">�b
�  �3�:  @�LN����ٳ��yt:�U�SE+�{�'������qa�;�^���?�[�n�5u *t�	�^�|pE���byy��u� F��� �*{+�sS܁$Z1�=Q�=�"ͺ \�w�R�,n��_�������0��Sp����,�	� W��{j
�  �e�; ���=�="�ĉ�y�������pSSS�c\����4+�4��}�# 5���[���Oc�O�T�( �P��^�X�T�4����+Y��{�  u�� 0bU܏;��~{�� |�`0H��>�d�]@�y���O����뮋���ߏ~�"3�`|]�!���ǎ��@+������V� ��Pp ��
� UK�U[�lq1�̙4������G�硫���wĎ���㺟����0��쏔>��{w_c�ƲWh��� 0Z
�  #V���;�B�������6��1z��� ������/�����??�c�� P'�&�GDv�X
� �E� ��� F���S�N�p8�	G�jz��s�p����c5�@��d��pCl�瞘�ԧb�g>�;"�RG���T�㽂�m�U�@;���XZZ�d-w ��Rp ����?b�yǏ��۷���9�A�jK�r"���P?
�7���+u(M656��ƍ1�eK�\w]D��: M�p�{8��;v,���f��n%�  �w ��jBñc�܁J��B�)��=�����Ŭɠ  �u�	�
� �s���Mw ��2� `Ī��Q�@DDQ1��M����G�-_4�� �q2�ܳN'fv�H ���s�_DE�'λ> �W彴�� �w ��j��;�S�: 4RG�"ّ#)�����^p����: pA�{�}��K��|�nU�K3� `�� F�����Ç#7��XS���I�7��9V�I!���nJ ���w�_�nIv�`��4�`0�#^�+� ���; ��UUp_[[3��\S�Y�{f�;@#N����r�Im����  j�?�k��(��ˑ#G*U��A �q�� 0bUn`t3�Xc���%]�w�f���&� \�yb�t����*Wh��_�� 0Z
�  #6==]�Z��l-����O��8y2iw�f��|�� p	�y�F*�-9{6bq����{h�N�w �Sp �*�UO� hb�={����o���; �%�kk���wK2f\TQ�ܕ� FO� `Ī,��={6M�*TE���1.K�o_��;W�ÇSGHn�RG  ���<����3�O .�ĉ���*[���V� ��Pp ����J׫r@D���`�����P?��GSGHjbÆ���O ��>z�?����m�'pQ�t=w ��Sp �*'�GD0��X�&��z�8��h�C c��D�IM_w]�  ���k�$W�ǏG���be�FPp h>w ��z���}�*]�Iܳ�^��+���1&�4�ژܻ
�  �4��?��$�$y��)V���(�͊�#� FO� `Ī.�/..�ɓ'+]ok*kg/��:BDD�;g�^p�Qp ���^��)���ѣGcyy��5� FO� `Ī.�G��T�Q�_y%u�����w0��<��N�N��	�  ���Sڒ]���Q�V���̦��+_ ��� F���F�S��,w�J��0u��9|8�.'\(���کSy�:FR�۷��  P��Ovf�ٳǎ�Z���Lp	�  ��� P����J�ۿ�&*͖�y#J�u�����n ��Z]�Jh�w �K��)m)wH2�O >duu5>\��
�  ��� P��7���a�߿��5��ր�v��˩#���@�>�:Br�k�M ����""�@Y�)� u��oF��t������ h;w ���԰ϴ�B�?5�ߏ�7R�x�	� �7XZJ!��͛SG  ���#�����S� ��T��Lp =w �����F���@��}�{��5*��P&�GLnڔ: @��(�'����>����(��7lؐd] �6Sp (A����ӧ��ѣ�����OpϞ}6u�Qp���Op������s  ���k�:�N�^{-u�Z8p�@,//'Y[� `�� J�j#��W_M�.0~j=�}0��R�����_ DD���b�IM�� �.���k�8�޽�:T��ڳgO��� FO� �333I�}�W�(�$k�%����c�W����^�b�;@����Iw �u��Vp"۷/u
���<���h1;;�lm ��Rp (A�I���q���$k�gP��v��ө#|La�;@�ΞM!�Ʌ��  ��C새��Fy_�pj1@�߿?�����?77�lm ��Rp (A�	�i�`��ZK���Zd/��:�ǘ�P��J�IMmޜ: @#���^�+�7ވ��S� H&���T��  �L� ���EQ$[��������S|��;@��SG  h�s������0��{S� H"��x�גf���M�> @)� � �F���R>|8�������g�I���]�ay��:BR��#  4¹���v��9�So��V�^�OMM���d�� �J� ���"|�W������{���^J��Lp����r�IM$<�
 �I�:Np��x������M`<�I�����t�� �J� ���"|��c8&� �_��z�ɞz*�����c�;@�WVRGH���  ��{���{�}8��� e�����3 (��; @	ROp��z��k�%� ��:Mq�}4u�Rp���O�̦�RG  h�|m-��r�sϥ� P��_~9�O�4� �
�  %H=�="���Ou)�g�E��T$����5�7-� ֧X[��~r<q"�C�R� �L� Pw ���ͥ����S�N���\m
�?�:�E�{i�	��0u��� �'_[�~�a�;0.�9G�MC� �$
�  %�������������
������][�x��).*7���ƽ��MM��  �����gO��j� �{�RG��z�� �F
�  %ٰaC���/F��c -6�(���g��le%i�KRp��q/�w� ֥��c0��WR� (���Z���˩cDD=Nu h#w ��ԡྼ�{��Mh����s˲GM��z
� �7��n7u �F��Q�O��sϥ� P�={���t�0� �,
�  %�ˆֳ�>�:�rIo$:�o�[��� pi���3� �e�	���١C�S ��g�I�}7nL ��� JR���[o�G�Mh���;>�l�ˡ�� y�:ARY�V1 �z��db�dO>�:@)�~��Z�����K ��ܵ  (I]
�O=�T�@�%��~�tdy+�� ��,K� )c �OS
�����N�N0rO�������  ZI� �$u*����+����:�R�� ���|��CE���{%
�A���&&RGHʿU  ��kJ�=�3 `�N�8���K�CLp (��; @I괡��y<��өc -UE��P���#�T��U�Mp�=ww �K��<����^x!�^/u��y�'�[�� ʡ� P�:�#"�{��7e��8k��G�XY�tͫ�4P�^p��[ pI�^/�A�"�}6u
��X^^��_~9u�����n��: @+)� ��n�~��?�|�@KU� M�G硇�[o�&��S��d�I)� \Z��k�5~����a� W�駟�a���6lؐ: @k)� �d�ƍ�#|�SO=y����P�ܳg��8y���F�i7����Opw� �%�z�țv�����M<�\�~?���
�  �Qp (I�KKK��/���P�ߏ�(�_�(��o��ΈyEͦ�a�>��0� ���8�=""}4�����~����z�c|��; @y� J�iӦ����G���@�E�
n�fO>q�P�딡�7�����L�I�� pqy��j�E�⋋���B� W���ǓO>�:�y�q� @[(� �dzz:���R������x���S� Zhuu���<�(w�)���ĘO].-��  Pk������G"�_O<�D-��G(� �I� �Dsss�#��c�=Vɤe`��K���=�xd�S�e2��:c^p_;u*u �Z[YY���{�g�Ff�	�0�^/�z��1.H� �<
�  %���M�Ξ=�>�l�@˔Zp���o������RG �"�}���; �ŭ��4�����"krI;�?�x�U����B�  ��� P��Np����~P�MA�y�A�y^�kg�>q�x)�]�B����� .fee%���./G|4���J�5�� Pw ��yckee%�y��1��)���� ��Oo���WWSG �":
�#  �V�������#"{���9��k �M�6��  �Z
�  %���O���XYYIh�2n8d��nd�O��u���z�# p�5~8�
��[ P��{��m(����%w�;}�t#�4-,,��  �Z
�  %��������x��S� Zd��3g�ӂ��C�jmŗ���>Q�c  �ҹ!!m9�-{≈���1 .h���1SǸ�,�j?�
 ��� JԄ��?�|;v,u�%F]p�|�k-�|n�;@�M6�{��� KK�c  �ҹ�{���8Ɉ��y��) ���ߎ�_=u�K�v�155�: @k)�*��    IDAT ��	�<���Lh�<�c0�����?�k�@+�1h��1���z�p�  �SE��{h�U��{�D�ߟ:��4����\�  ��� P��Mؔi@3�j�{��{#�b$�Um9����}�{DD�С�  j���E���D�
��y���<O�}M:ux�ƍ�#  ���; @�65h
��ݻc8����(
���OG�w�����io ��d�>��eU� �cVVV��qѲ�{��Nt^z)u
���X]]��~8u�u3� �\
�  %��������1�������SO������N*_[��W�:�05b�;@�M)�G����  j�����6�=""����6����y�G>�PQݙ� P.w ��5i��������1���_����7�q��Ճ�;@�u�mK!��ÇSG  �������ʂ��rd��~���;v�X<��3�c\�&�� �D
�  %kR����Ƿ����1��+�"�Wx�7;|8:�����C��Pk��11;�:FR�C�RG  ��~�kkk��|�Ƃ{Dd�<��|�D���o~�W54%w �r)� �laa!u����oĞ={R� n�J��E��q�p8�@5`�;@�u��6u��z��  P+��(��JQD���ݓ����C|�z��ͩ#  ���; @ɚVp������+++�c v%ܳ��l߾ч����;@�M�y�}��k'N�� P-�����ĉ�<�x���Y\\�Gy$u�+�� P���  ڮ�������w�?�3?�:
�P�~?���,����٩Sѹ���S���z�# p	�m�RGH��޽�y���1��G���[o����,/G1���LL�����B��v[Lnڔ:& 5��! E['���裑���σ@E���\Ѱ�:Pp (��; @ɚ����/��w���rK�(@E�~?������ٟ�iD���ED��?@t�oO!��{c�O�D�pU�Ǐ��k����^���_�3���o�����n���;c��xl�ɟ��O~2��0\�q������e����yd�gQ��/F�sh��z饗b�޽�c\�n�6lH ��� J�����x����_���v��� ������{�䓑��b��Rp���;RGHne߾�`݆�˱�o_�ٳ'�_=ξWj_;y�_s�ĉ8��q��G#"bra!�������\,�؏�*: ����cPp��8t(�瞋¿{@����c��ݩc\�����  ZO� �d[�lI�-..��������/��4��:
���bt�4�)����M7����rC���bE�Ç���[��o_����o����E���җ,.ơ?��8�����7�ʯĵ��\t��J_��Ξ=��_�k��ߍ��#����w���>H��#  ���; @�6o�Y�EQ��\�g�}6n��ָ���SG���GQ�]�H뢈��0�<7��h8&7��l��SGHny���8��]٤�c��?~<z��Go��Xٿ?V�|����z+�5)�,��{~�7������������o�-�?h��Np_[K�$�����w_��K�N�4@�<���gϞ�1����|�  �g� �dSSS1==�^/u�+RE<���˿��1;;�:� EQD�ߏ����~=۽;��_�8U:�2���fn�!���(���Q��8?�����tb���c��bÍ7��1�cG��xc����m�".��G1D�С����
�y���W��������Q��k�[��SG`���yO�+��i9z4�G�ⳟM�h�S�N��ݻSǸj&� �O� ����-�GD,//�7�������Ob8�����ܳÇ�s�}	���P��dt��.VL%�<�����;x0N?��Ǿ��v?^~߱#�w��뮋�5�$MJ���X=z4V��#G~�����;t(�G���ᑕ7ߌ��?��~��b��zd�#0"������������?���(n�)u��<���?�-xXH� �|
�  XXX�w�y'u���o߾x��g�ӟ�t�(@���f�`����#��%���n�I�}�~?V�|3V�|�_�t�ѽ�ژ޾=�����_w�|�1�u�BpC���/������ñz�p�}��~�PWVR�L�ȗ���Ÿ�����t��� 0+�w��k������#~�W���	} ������ÇS��͛7��  �z
�  شiS�#�{����c۶m�� ���EQ|��Η�q�P�Ti|��8��馈�K���~?zD���~O���Ԗ-1�ukt�o��֭�߻۶Ew۶�ܼ9�6o��M�"�&52E���ԩX;y2�ǏG���X;y������ɓ�v�D����'#o��Ų��x�������-n ��ٳg����6�=""Μ����ٟM�h����9���lْ: @�)� T�-���a|��_�_��_�	7�u(�"��~L�7�k��T�����Jc즼4Ԇ�nJaly�~��쫯^�{�N'&7m��͛���M�br���n���7���BLm�7���������;SS������pi)�c����/.��̙w|���S������[������o�f�������z�k��=���Wc�ƍq�̙�I���zq�}�Eޢk��  ʧ� P�6Mrx�w������Z�(@C������t����'6o��"u�$��&8@�(��S���O�\�n�C��ɍcbf&�n7&fg�397F61�7F65�������N����+,O��E��|���~?��Lw��D1���׋�ߏ�ߏa��p��rE���w��һ���./��̙��\Q�^�|�+1s�q˯�j�( \�Mo��	��yǎXݿ?���SG�(�����c�k�6��������1  ZO� �[�nMa�^z�رcG���h�(@�z�ؼys|򓟌�+(����;@3L�xc��X��G~�D��8�:
c�������㎸����Q �g.0��(��.�O���w�/��R>����<��ño߾�1Fjaa!2'6 ��s�o �j�����o;<�:� kkkq�w���|L�̤��L��a�*@�m�馏M��,E{����U�� �t�	�kkcz*]��D69�n7n����q��ػwo��?Hc�Lo ���; @�l��N�>z�y��w�#i�K���k����LO'N���w�ڛ�����Oh���3���Wph�~�k�Ҟ�������������ǎ;'��ԩSq���G���6mڔ: �XhW�
 ��&''cvv6u��[ZZ���/r7������n�)Ξ=�1���+�4��Ν�# -���3�����c pΜ9s���(�������ϯ��zO�������_�r�[�`Ж-[RG  
�  i둅o��v|�{�K����ɸ�;"˲ܻ��'~����7u �fV���������J�u:�q>���z�#�,���n��1?�8�o}�[q����1J�y���  Ƃ�; @Eڼ���O�K/��:P#�N'��Θ����w�����Y�1��9��RG `6*�#���������c �EQ��������C���˙���;�3&''$���k����[���  0� *��#[���?��?��L��s뭷���܇~��M≙��jA���܁:��#q��S� �VVV"��~}���0�������;��Q; "���?�p��Sp ��+M ���y�{DD���|���N�s�7�w���1��<���� M2s��1�aC�@���/�%���&H�ܾŅ�u��"{97n��n���0@-<x0����GQ���*˲��kR�  
�  ���~?��ދ��۶m����?��Ξ=EQ�u�=_]M�u�:������1�Y޻7޹���1 ��K��������ٲeK�ر��4@ݜ>}:���p8L�t�����vS�  
�  ٶm[��X\\�{�7���RG*�����r��>����D�a��: �4�sg�@˼����)� 5��y�.q͞��~��:��p�c1���������86��6mڔ: ��Pp �����SG�̑#G���܍{6l��o�=�,����={62�h w`�V�z+N<�P� �Ǚ3g�(��~O1����:��v�m���Pr�.��a|��_�S�N��R�-[���  06� *2==����cTf�޽�{���1�
t��عsgLLL\�{Ϟ=33��'w��ظkW�@�?�'u ���ٳ����8Op_g�=˲��'>1V��0��<��~��q����Q*�
 ��(� Th܎.|�駕ܡ�&''c�Ν155���_^^�0���x�=�MN���̩���7�L��8s��%����9�W�aÆ)E_���c�޽��TN� �:
�  Ǎ�'�|2{��1�LNN�]w�3�9�}u�˂
� �љ���wݕ:�BG�/u >`ee%��%�/��+HSO��(�G���޽���_Q��o;^y��Q�ضm[�  cC� �B�Xp������O<�D��MLL\�4�^g|/E�++�# p��GSG Z��W�Q�c ��Lo��k��
N㛚��]�v)�C�<��C��Ϧ����; @uƷU  ����#���|��R� F����w����W��W;��:�py9u .��;P�ޡC���۩c �����T������n�;w+��@���0�N�3���  ��� P�q��PE|�[��c+�-Ε�����E��b\���x�@m��Kh����SG  "�A�z�u}o���k��Lp?gff&v�����#LT����{,u��bbb"u ���� P�q.�G�[r��׿{��I����W�:Y��Z����(�;vD��kR� Z�w�@� ����GDǹ�~��7lؠ���O��ݻS�Hn��ͩ#  �w �
mݺ5:�����y�����/��\�N�w�y�U��#":c\p��g�S�Jh��	� �p9�|u��$�v5�ϙ���]�vE��A"�*�?�x|��ߍ�(RGIn˖-�#  ���nW Tlbbb$�Ц��<x��xꩧRG�abb"v�����#y���L"b0�Wk��g�ӟNh!w�􊢈�gϮ���q��>��{D��̌�;4DQ�{��x衇RG���[���  0V�DD��aP����]�N�ژ:GjEQă>�~?~�~*u����b�Ν�aÆ����{7EW"b4����W�uv=@sm��Oh�ށ�# �������|��?�����^���Ʈ]���W_����B������O��R+7n��S� �	Ûa�)������H`���+�C���?kkk���_H������뮻bf�71#"��
����P��q��'&��c���:
�"+��GED���0��.��	��������VΝ���/��R;��{�߹��{N�`��o��rD�n��H�r ��k����?�w(RG���v���y�=��W�ݣ����M[���tb�g>�:�2y��'R� kgΜ����	�#.�GDLNN�Ν;cvvv�\��p_��W��/��  Ɖ�; @�^I���|����׾�� u{���q�=�D��-���k]ĻS�ǉ�;@3m�	���ۿ?u�����kkk��{�y��D	"�-��ڵ+6o�\�������O��O���_O���Eĩ�!  Ɖ�; @�Lx��W_}5��O�ı����͛c׮]199Y����R�*����۟�܁2�H`l]���(����r�4@V��s:�N�q��}���� .�������q��Ӌٗ:  ��Qp ��+1L��:�'O�L��������o�N��K���~���I��b��Q�ӟ�6��S[������;@:�������1����ae�����o�,�J_��s�dN�8�:J��M  `�(� To5"�Qg�O��?��?����c�[n��&��y�[ry��j� \�,���ϥN���![ )���E�2��8ܳ,:�n%KU5|x�Su/�k�  �W�  i��:@��z���?��x�WRG�V�t:q�wƵ�^[ݚ�)�R���0p������O�� ������# �������=�<�}bz:�©�7o�]�v���dek�8z���k_�Z��Q����  ƍ�; @�����0���x��G�(��q�u��n�}�ݱiӦJ�����w�����|e�*� ������L�F���2�$/���������4;;��sO���V�6��`0�o|���|�}���R�   �� �4e�NEQ��?_�җbuu5uh�������cÆ���MLD�S����wMph��-[b��S� Zd������R� +�� V����q.�O|dPAU�fضm[������������_L�i��p�0 @�� Ұv��x����ǎK��믏��+����e�LO���4��w�����?�:�&y���N0V�dz{D�p��=��JY�ŭ�����'��4%�*o��v|�_�#G����DG#b)u �q�*  �1���S��_���"p�:�N�~��q�7��rނ���;0����|���# -�z�`� cei����c=��#{8)lݺ5v���n7uh��(����/~�l_�J�K  `)� ��jD8��
����7����7#���q�1fff�{�-[�����5��~�(����X��dLmݚ:�"�RG �� V��T�|uu�i�#�I�|vv6��XXXH����W���x衇�O�:�� ���ޝ��y�����e��C�p'%n")���p;���i��@�<-��E���&���i� AQ�E�E�hN�i�x��h�v9�DQ7�E�9��̜}���Ő#�8$g9������`0�9���HQ�������(�  �hI��:D��;wN����c��l߾]�=��������*Y\�}�L �K����[�e@�ԙ� ]S*��;?��	�ZO�f�:r����c����)=�䓺t�u�$��:   ��(�  ���:@�MNN�����~�ӟZG")���СC:p����h��K�r��+�o�	� k{��?S*��� !(�@��J��\���?}
��T*��{������]e}	p]:uꔾ��P(X�I���   \��  �[.ZH�f���{NO?��|���~�g~Fccc�QV�Yeҗ����Lp�x�ݵK�~�W�c H����� �	�﫺�����-��ĉڱc�u 2J��������?��� ���$g�   ���;  ������ŋz��'u���(���S��;����8�t��_.T�}&�@�����:��h0� ��T*)��|
�єN���~>|X�l�:`��ŋ�����I��%�[�   pw   ;�$M�Xd:	���ק�ǏkϞ=�Q(�˭�y
� �8�ٟՎ����c H���"�@�J�M�|�����5� JFGG��c�ixx�:
�u�fS�>�,��v�Il8  ��  `笤��ª� ЩS��������tE*��Ν;��c�i``�:Κ�ksԓ��m�7� I���L�u 	Pg�& t����T*�����3��~�\.�cǎi���J��A������?�s}���Q��#�    ��  ����)�I5;;���˿ԫ���V�e蘁�?~\?�p�6�2�������L��d��ܩ��w�c H���u H�b��0�ܜ�^oS��I����ڱc��q���ZG:�Z�����SO=��*�@�=   `$k   �q�$��TA���������h���֑��I��ڽ{�v�ޭT*eg�R���U��UR�~UkC� �c߿����u�Ο�� Ƙ� �U,7}���	��RU===:|�������lZG�"C}��z��WUw�ƛ.�`   �U��  ���f�    IDATLm��BA�������O��D�c�=�={�Ĳ�.�s4���mc
� ��\N������ 6��; tN��R���]����a����[��ĉڱc�u`�
��������c����Y   p�  l��:�K.^���ׯ��_��}����ᮞ��۷O۶m���i��U������k5� �6�ݵK���ҹ��])�� ����u H�vLo����2i'��)��h�������`Ď�yz�w���o��<�8���w   3Lp  ���.�V�z��g�����$%�D*��Ν;���'��.I����>^�v'J�Lp�����/��o$n��Lp��)
m�����^p�mxxX'N�СC����cX���q}�[��o�A����ZZ�  �&�  �:k�U�������+=zT��˿����H�����u�����ZGi�m��������<
� �H{��U�$]�/�E
�z��NhLMYG �Dj4j4m����S	)�KKC$���422���iMNN*�f& �gffF���
Cz�]�   �2^�  غ))o�Ua��ŋ�ַ��7�|�	(��|>���ڻwo����ڦպ��BPK� ��_��?��(� X�Z�W*Y� ��i���0�Zm�Vep
_e�Y�۷O'O�����u`Y�Vӫ���	��q�:   �˘�  `_��2����o���_�%;vL�T�:U�T��[o����
� �7^�װ9Z��K�t<Mw�Lp�D��ۿ�t�.���(��� �QsfF��a� �(�b�-�q�F��)��b��7�|S�җ��%�ر�:�l6u��i�:uJ�f�:>q�:   ��(�  ػ 
�P,��3�護������������5�ZM��N�>��Ԟ؂�6GC-Mq�x��
}_A��t.g �!;�74t��~�����eN4�`��i<�u H�j��V����F[�WkYÉ��F�\���W��СC���H�]�y�Ο?��'O��P�(z�:   ��(�  �;o +��y=��s:u�~�~AG��莎���:}���}��U��$���㭫J^�]Z��N� �m��A=��o���Ϛy�i�8 "�13c �]��%ɯ��v��I��(�Mn������0�����\���G��_��FGG�!ɂ ��￯7�|S�J�:V�	�   ���j   >N[��������Ok�������y>|�:��l��ٳz��ո�$����:��������x��U�l�j �a��=���i�?�'��7T�x�:��jRp��	ð�������jS��0�ŋ��G��ѣ�җ�����M� Ї~�7�x��O�#�hiy   F��   ��w%��QSSSzꩧ�w�^}�_СC����V�:s�Μ9��6H�ZpOe2J�r
V�Z�iUI#���UA�f �E[>�y}������_��j��[G1��i� ��Je�d��ry�{f�
�j���m���.]�������^۷o�b:$I����￯��{�b{||`   �u�  �$ݔ��:�orrRO=���l٢�}�sz��ǕM��h�B��ӧO�ܹs�*�'��.-m����^Q�
�G�{�i����T�~�75��˚��wT<�aN �0� �gqq����ն^/N�^p_ˍA��p�P�n�jUgϞ��ӧ�4��r�:   ��h�   DÇ���BA���N�<�'N�s����c!�&''u��i]�tIA���'������0����Y��O�=^�l `$�ӣ�����뿮�ŋ����|S�>�6��dh0� ���}������S��	/��o��jn@پ}�~�gV'N�P&��P:���ܜΜ9�.��D	t��    ���  �K�U�X�j��S�N����:q℞x�	���Y�BA�K�.�w���&�*I.�g�����%���Sp H:vLCǎ������bQ�'O�x��*�/�z���ss�t	��=
���0l�5]��N�}usssz����[o�'�Љ'400��t�� t��5�>}Zm��]��u    �Qp  �����q����ٳ:{��v�ܩ�|�3z��G��嬣���������i�3���l��$��K�]~�b 1ّm��_��_����y����/�2>���K�������\�_�*C9 6eqq����.�'�ߥ�N�.��������'z衇����ȑ#J������(�����t��Y�pZ%b�&�u   �Qp  �&A$��̌^|�E����z��G���|F;w��}_�/_��������}2�F'I��z&�Z�U�X���J%� ��k�'4��+>ߘ�^*�_���ի�ML�z�����FI�CczZ�Y� �ت��j4m�nP����q�a���A���	MLLhhhHǏ�g?�Y�������� t��u�?^�.]R֑�^iiI   �(�  D�YI���,1�ͦΝ;�s��i�Νz���u��1�%|S�%��Ӻp�>����l�޶�IRQ�^G�]�*JP��	� �M�ݵK��vi�_\�y�Z]*�_����v�j
:��
��h��Pp�M���vi�{,W�����	ð#�n�rY�N�һﾫ��ĉ:x�Y���`nnN|�A[O�D$��:    (P  DE]Ҹ�c�A�~333z饗��+�h���:v�}�Q����{�|^/^ԇ~�����<��y]y��.I%�N �\��  H�����O����w=���߸��v���Ǔ�R�O��~͹9� [a�X,v��.�3�:��knAh||\����f�ڿ��=��G�Rv���k�/^T>�����8k    ��   $�yQpO� 499���I����:p���=�GyD�\�:��z#��L�H���(]�Qp tYvdDC##z챻��O��7n�~���͛�OM)��#�r۶�w���٣�={T�qCs/�h�Ts~�: �V�T��)x~�֑��A���:B�ts������/��#G��ȑ#:x���t�r`�Ţ���u��EMNNZ�A��c    �  �䬤��:�����M�L&������:x���9-MMM��ի�|���K&�V���;)������T��t� Q��бc:����A���ܜ�7n�9;��q��ǵkל�l��eGFԷo��[n�v��ء�}����]aO�t���b"( l���bǮ8�}N:�'PZ�h6��p�.\����>>|XЁԷ��2�ǝk�W�\���u$�	%�m   �  �����}_�/_��˗%I[�l��Çu��!=��CL��j���ׯ��իW=BSJ;5},
��$�%5$�}��	� �8I��.��掠�����SSjLM�9;����Z�����j-,����0��۸"�N�gtT=۶�w�N����w�N��޽<��w�n��yJ��#�t(q|4)���x��jK�.Op���{q�S���r�=�Jiǎڿ����Ϻpܹ&|��e5�H�����   (�  D�I� ��B����{O���r��~�a<xP�����ؘu�Dh�Z�����Ą�]����Y�ahkUQ�l��7Iˊ��	� ���U���1�����rٽ��/�o}|g�9?/�R�Rz�s9�lݪ��[�UntT�[?�Sn���	�=ccJe2mϐ۶M=��j-,���q�w ؘ��Ŏ��|R��	�P333���ѩS���߯������ڳg�FGG�#�^�����nܸ��W�jnn.�k�0��u    ,��  3�nJ�c��l6WLw��rڽ{���ݫ�{�j߾}�t�\�4�jUSSS�����䤦��c3��jYG蘍��Iq�a�w ��n��u���6h6�-.�9?���rY^�$�X�W*�/��*��ˏ��E���f���hI�rJ��);<������;�2����z,34���Q�mSf`�:�$i��-���u3�`c
�BG�����Nߋ�����j5}�����%�.��JE7n��͛7u�ƍH9A���   �%�  ��(��>�ͦ&&&411!I�d2ڵk���ݫ]�vi���ڲe����6�M���innny�X,Z�ڰ��7"��"U(�"i��i���;  ���۹S��;��s� �_.˯���j
j5y���z]~�.�\V�j)�����x�T�$y��B�_z�Se��^W�Z!���m��R)e����tvxXJ����W��G�f��U$�Y�}��W*�UvhH�>e���Rf``�Ǚ�!��`��a����y� ;�JE���z��7��������p6��Ν;�w�^�رC۶m��ؘ��JeyMxzzZ���*����y�:    �Pp  �����b�����T����FGG�k�.���illL�v����a���@�RI��󚙙Q>�������|�&��m�m=6:�]�ʒ�$�ږ��|6�  �T:�4��VI����C�L�A"nV �nY\\����j��׏�ͬ�D]���<�[u]x۶mڶm��o߾�6�ʍ�q�j����5;;���9���kvvV�z�:��u    ,��  -�Y@�A���y�j������l٢��amٲE###��GFF"9ݧ^��X,�P(,�/�J*
*
��n~[�7��g3�\{����z{"l�7�  ֫��{���
���ZG�X�<O�[��tJ�x�=���wj�v"O�A���Y��ή�|&���А�lٲ�622���!j˖-F��v{�I�PP�RQ�RY^��F���&����q�   XB�   Z�=�W�VU�Vu��ͻK�R��������߯��>���-��߯��^�r9�R)��i�r9IROOϪ�f��0��qѭVK�VK�z]�ZM�z}���?��j*�J=b:.���v[v``S?����%�+����  ���	����)��-..v����j�~�e�n������rA|5�\nյ�;?��rJ��J�R���$e�Ye2IR__�Z���@�F�!i�����u��P��\^�sm��5b
�0�SI�  �
�   ��:��93�������򦮓J���f]��$o��7Yp�K�%eڒ���rY��ۭc   DF߾}J��
��:�����y�: D^�Z\\����OpO��(��c�c��f��f��b�h�v�:    >q��E   X
�4!��0)��Y�7��}}J�2��B-�W^��Q  ��t.����|�: �B�\�����L�u��b�*�X   �'(�  D�i�  �#��T*���#�7����8�I  p/��;�#�jQp�5���vI
j��<Oe6y�^�%y����i    ���  =�X ��YG��n������w  �����a�w x�V��J�ҕ�rz�{��Lp�)uIg�C   ��  ��	 �%}�T;6K����~~�6�  �$�z��X��  �����0��yn�������:*�kn ��$�|  �
�   �sN��kh��o�eڰYZ��9�^�l   rr۷[G0��=" �W�*
]{>&�'W��� ���    X��;  @��޷ </���k�fik@�  ���w�T��  �V*���V�r�=��	�I_s�n��   `%
�   �Ĥ ��?M�]����N�>L�  �[��uS�����|~���狒t�'�7� ���    X��;  @41)�����m�H��L5&�  �-�e�uS�	 ��h4T��Du�'��k�&�Z��u �Q�t�:   V��  ML�  )��m�6N�۬K�K   w�q���w ��|>������Mx�=�C% ��I�u   �D�   ��+~]M ��{;���$��v��c�;  ��z�n��`��; ���}���?���3mJEI_s�.g�   �n�  �)��� �K�4�vo�Ʃ2N�  �n��a�2�f�fSA�_ �F,,,(��?���t��I_s�.��   �n�  ��u  �� ����1:�����s��O�  �n�T�'�>S�`�0���`��~�f�Q�i�{QD��ް   ��Qp  ���� DC��L��fi\�@Lp  X]�u� �R�T��u�v���R��5�I�gI^o�.I�C   �n�  ��u�  �!�n��,�J�����Gq	  `u�>���� +��y��uyz�$�~�Y��� ��9�c9  �9�  ��#I��! �K�ɝ�,�4v'�VKA���  l���)��'�ժjFEs�Z5yިH��ǍF�:�h8e    ���  mg� ���R����\�,)�ȕۋ)�   wK����� ����.I��ܳ8u/J<ϳ�  ް   ��Qp  ���� �����$�a��  �ݒ^�{�� @���eÿ=�'���i�r9����6 ��c�    Xw  �h�;�  �%y�{��O�tg^�ơ�W*�   "'��g�TP�[G �HXXXPڝ�8\p�8p�w �nJ��  ��Qp  ���%�! �J�[*�L�
LIQ��c�;  ��:u�O\��@Ahqq�4�_���p��B�=�% ��{�   po�  �mQ�� l%}í���Q��{�G�  DU��{�hXG  s����}�4�˧��PpO�@	 k��u    �w  ��{�:  [I/��;�iZ��u�����   "�S'��EH����0��u�oJ�ZG�0�o� 	g    �F�   �NZ `+���CC�v�hOq�JQN  `#�w� `�T*Eb-įV�#�Iz����� $_қ�!   po�  ��5�  l%}�{�7M�Zڭ�"&�  �-��XG0���� �����uInOp��0�(H�Z�5��h�F  pw  ��{WK�L ���ԲN�v��H��4w  �U��޺`�; ���e�#r�����#tw �NY   ����J  ����! �I��[7��.k��5�B�:  @����Q= :/*��%�g�{b%}��59i    �G�   ޲ ���$U:�,��w  �U8>�]Ao��Ϋ�j�Fhj��p�=��)����u    ܟ��   ��c�  �$��ޭ�`%IaW�i�(�  �-�����# ��(Mo�$��[�#��	�I_k�@yI�C   ��(�  ��KZ@�AI�*Ս	��K���%�  �b��u �f��R�dcY��k5�f��Vc%�km �u    <���   �1'�u 6�>U������*_�*�#   Dw� �usss�V�U��}�Mx�=�km ��    x0�W�  b�u  6�>U����-IQ���W�
=�:  @��2���?��V��b�N8��e��2�:*�km �U�    x0
�   ��w� �H�T�nO����m�  Xs��0�N  ]���F��>�Z��`*34d�����ྚb�;  @,Pp  ��W� ���M�t��[oQᗢV�  ��J��u�|��S|����u���.OpO����N�QLp�vVR�:   ��Ub  �xy_Ҝu ݗ�M�L���S�f��
�   �$�����!�|^AXǸ��p�=;8(�R�1:*�km ��-�    X
�   ��u  ݗ�	�J����S��)�^1Ju{   {�㥳t6k �"-,,X�X�W�XG0���I{���~^�   ����  /oX �}.l�Yl�F�VN�  `���;��b~~^��[�XU�p�=��!��8+���u   �w  �xy�: ��sa�-cPp��w
�   +��(|�f�	� \����܇��#t��$ �ꊤ)�   X
�   ��w�F@���1�<�B���;  �J����O�	� ����;\pO!�6�I X�I�    X;
�   �R�t�:��r��n�y�)�-
�   +�Op�� �>�]��r�:�����u����8�U�    X;
�   ��c�  ���@�'k8̺^�w  ���R�:��L�u �|>�c�    IDAT���9<�=kt�^7y�g��Y   ��Qp  ���� �.6ݬ&�K�S�)�  �Ԛ���`*���\ �
�@�|�:�yOp�B�-Lp�4)�u   �w  ��yYR�:��i�������eŜ�;  �JM��Y
� ,��%ɯV�#�ISp�LoX   ��Pp  ������! tO��R��1:�z��r�;w  ���1���I��~� �q��.I��܇��#t��$ ��5�    X
�   ��w� tW�7ެ'�KvS�)�  �!�ZX�Na*�w 	���a�� ��0��¿CLp��#�    X
�   ���u  ݕ�{&��$���V�(%|B?  �Z5��z�uS.�'N��=���K�X�鴤���˜��Z�   ��Pp  ��$E���I�d��l�.<g�y�k5�g  ���ĄusQ�� �i~~>��%ɯT�#���){���u6 wy�:    ֏�;  @<Ŵ	�)I�,��� Ijhi�{��
�g  ���ի���FG�# @[������k������tw�9�Y   ��Qp  ���X �=I�x��t0���_*<+  @�ԙஞ�[�# @[�iz����tO�R��u��K� 	 wy�:    ֏�;  @|�b @�$}�-��)��cC�ԔT��s2�  `I��5���$H�Պ��v��{f`�:BW$}����X�   ��Qp  ���$�! tG�����������]|6  ��9^pO�rΔ�annNA�%L��{��f:Ʌu6 ��Pw�z  �&Y�    ذ���%}�:��sa�TfpP��E�������wk[��;\��*�9��ŋ�\���������k5y�ʎ�(��)�}�r;wj��!=��#G4p�RY��  iB�S}r�:����Q� �6�fS��X���̸Pp�P��Y� �=�X   �ư  o���;�&Ke#��Z�4 )Յ��T��5����UU>�H��8����97'}��򯽶�X��G�i��9��c�4x��r۶u��  ���
/�Qp�$���
�����U�f��6�	����T ��u    lw  �x{A��Z� �y.Lp�YGX��T�ԍT�N��"h65�쳚��wUz���]��R��E�/^\������)�G�j��Q>�t.׶� tF�j�x��us��ۭ# @[��ucz3���Dsa��e3Z:	   1D�   �~$�)���p.����r{�{����J~���VK����>��?Scf�k��ZX��ɓZ<yr�s�LF�,�����#��o�>�2��e ,i�̨61��Ą�׮�z����ON*�}�x�zwﶎ  m1�����W*�̸Ppo4� t���   �q�  �,鬤/X�Y.ܣ6�]�|-�E;���a�;�d�'?��o|C��	�(����UWu|\��?���tO�������C�o�j��A&��&�ժj�ML�z��j׮-���5�ժu�H�ݵ�: lZ�ZU%�%q/��7+�k3�F�p�K�   �q�  ��5QpυͷL'�KRIҐ:;��g�;��Tt��_�����u�5	Z-U/_V������߷O�w�V�����{
 ,xŢjׯ�~�[��U�~]��Y�x�E�@�����\��`ƅ�<.� ���    �8
�   ������:��r���)a�����|���b�t^������=�''��l^,4?�X��^[�P���8xpi�����}�!�?�����Q*�2��i��/�W��~]'�tD���� `S�岪1?���{vp�:Bǹ��@�tU��   �8v�   ��I5I��9 t�ӥ���Z���N�����8�}�y]������Q:�15��Ԕ�|s��S��z��Q��/�zH������ջw��==F����fS��7U�yS�����z��{?��8�� ��0��̌u�M	=O����e"�6�.�g�n    �C�   ��ޑ���A t��(o���
��u�����R*աg :��w����G
��:����U�~]��׵��w=����C|���۷����2��"h�Ԝ�Q��5gg՜�S��ծ_W��5n�t���(I��(�k�u ذ���ؗ��R�:��lDO�k'�� H�^�   �͡�  ����;�hq� ^�(�%���)��v�jɯV#�{ ���w��K_��u�X��EϜQ�̙��R�ݹsi�������Sߞ=ʎ��A��4y}rRͩ���>n��YG�:��ۧT&c 6$�%���\��`*���.��P(�9�   �
�   ����?��s\�|�Ơ�]���C�n-.RpGl�<��.��1�/՘�VczZ:uꮇ3���۳G}{������={�۽[}{��g�V�� �%h�����̨q�9=��~fF��7)�'L���� `�����y�u�Ms}���.���EI7�C   `s(�  $�O$-H��3\8>9�MԆ�&�wb�YkqQ}��u��@{�Ο�G_��� ���x~��ʥK�\����������;ջk�zw�Vn���ڥt.��� �"h4Ԙ�Vsvv�F���SS˥�f>/��uTt���� `CZ���c����8�,
�^�   �ͣ�  ���J���:��pa�-;8(�R�/r$�KJ�������l�|^��U��M7q��j����:>~ϯɍ�-���,�S�:����[\\1u�9;���)5fg�
�1A�����쬂�� �r�=��)��c��\Xc�g�   `�(�  $ǏD�H,&��2ez{����Q�˓T�4����|E��� Ї��j��XG�:4�y5�y�?��_ӳu�z�mSn����m۔۱��cc��ܩL�����E5�y���՜�WkqQ͹���Ԛ�[z|aA��[GFL<h ֭V�����|��١!�]A�H����C   `�(�  $�S���:��pe�-;<���$%JJ���u׿�M-���ut@kqQ��EU/_���e��W�o��{��Գu��[�*76���Qe��ؠ X.�7�����j��.�����z>��������TJG�X� �u�I��^�l��+w�H �{KR�:   6��;  @r\�4.�u ����[vxX��Y�h�侵���(�#�Jg�����u�k5�&&T��x�צs�����r۶)�u�r	�w�6���.��g�VeGF��+@R���V� ����o߼���Z��j-,HahXֻg�3�B �Q,U�V�c������p�Ϫ�&W�� ��d    �A�   Y^w �\����Q��,iH�{a�wDU�h����^�u	�M5gf�\�D��Ȉ��ß�������(3<����ǕJu�W�n�MyŢ�Ri�7���K�u�'�"9����  ���fcp��z�\p�:Rp����@ ���   ��  ��9I��u ��J�=N����EI��t=
k���v�u8�+��ҍ�����ae���W������Ko�=�������L����P�hȯVz��RI��)����j�U��R	�RY��Z�_��/���zܯV��뷮���;��YXXH�$l��{�%��-�es�NY�   @{Pp  H�g$5%嬃 h/W6�⶙Z�Ԑ�ۆkQpGϞ��'���<����T*�Q��O��{{�޲Y����J��O�+�J)30 e2���)�[�-y��W���ߦ��Ye��J���b�y
��{f<O��O�I���˫T�>n6ܺ�ίV�*���� X*�7��+���W*)\�� �c��;��}_sss�1:�	����	�Q�ii.	   ��;  @��$�����A ���y�}_�L�:JG�qj]Z*n�G�4���?�)�� &�[Ep��A 8a�3���  k633#���ct����7o&w �~d    퓶   ��{�: ��pa�{6���-I�6\���І� �s�O�D��q�  $^ߞ=�m�f ֤^��P(X�舠�P�jY�0�w 1Jz�:   ڇ�;  @���u  ���\'�KRQ�fg������+Wt��'�c  ����~�: ���Ԕ�0�����'��uMf�\X_uQ҄u   �w  ��yCR�:��sb�{L���6;�.�:�s��7��g  '?��u X�B��Z�f�c�r;�g����ɬ��k��^�   ����  �<��W�C h?&L�y3�"i���Z���l��K/)���X�  �[�x�: <P������Q�R�:���Аu��pa}p��Z   @{Qp  H�g� h?6��\p��EI�9���;��������c  ���А�}�: <��ܜ�����^p����Z���8�"��   h/
�   ��I�u ���ʙ�A���}�ڔT���o-,�+
�!����Rcr�:  �������fS�|�:F�yܳJe��1:.��ߨ8�5--�   AX5  H�9Ig�C h/'&L�R�?� )���e�;,5����e  �l���# �MMM)7s^Y<�\p��|-f��X[���u    �w  ����u  ���&\&�Gb�Z*�owX���UA�n  ����/ZG ��*��T*�1��+��#������rempL��S�  �0�  ���Z �^ͦ��fc^p���6v&�G�FO����/[�  �)�?��Ç�c �=A����]����Ȉu����$��&�C   ��(�  $��f�C hW6ᒰ�J�HU�	�0������u
  ���W�: �����Z��u�����|�� �i�   	E�   �BI�X� �>�l�%�X솖&��wX�}��Ο�� �s��ʯXG �{j6�����1���{B�b�^�[G �~?�   �Π�  �lO[ �>��45� )X��SpG��&��O�S  ���ؘF>�� pOSSS
�����?����u��pempHQҫ�!   ��  ��)I�u ��h4�#tE�6U}I멬SpG����T�r�:  ���4[4 ��P(�RY�d1���e�f��s?܁�yUR�:   :��S  �d�Kz�:��pe.i��Ik�5����.
Z-}�?��u  �4��/[G �U�����i�]�W�
�X�L��b�^�[G �^�Z   @�Pp  H�g� h&��W^R����U��� {�?��W  ����/��u X��̌|߷��u^�d�T�bV�������Y�   @�Pp  H��� �=(�Ǘ'��֯e�;� �<}�gf  '����P�\�: ܥZ�j��פܓ��W�� G�+i�:   :��;  @�]�t�:��se�Tvd�:BG��Tt���et��3Ϩ19i  '���߲�  w	�PSS��)�Sp;O[   @gQp  p��� l�+�p١!�Jʯ��(��む��  :~\C�>j �2??�̺�j|��tZ��]��q ��g    �E�  �?� `�\لK��(��g�#�*�
���^P��5�  8��� ���lj~~�:�)�\��`&;4�T*e�+\9p�ǒ�X�   @gQp  pÏ$�C ��6�2	>� )��㭅�nE������  pR��O;�7�c �]����{��|��ܓ��i�� ��u    tw   7x�^�`s\ڄ�I��/�~3�)���
ﾫ��1  pҞ��me�}.�x*
�Tt�X�|��K�6���$�  8��;  �;�� `s\ڄK�����{��l��݌������:  NJe������u X��}MOO[ǈ�'�gGF�#t�K�#	V��u   tw   w�@R�:��si�ǁ�ռ���o��w;
ј���k�Y�  �I;��?Rߞ=�1 `���i��o#�B�:���Аu��qix�`/��.   'Pp  pǂ���C �8�6�\8��Ҹ�Ok-,t;
q��'�`��*  @'��Y=�;�c V(��*8\��4�'�Sp/�V  �
�   ny�: ���@��Y��

�T����f>o	�W�����c  ऽ_����﷎ ˂ �͛7�cDG�+�v�\Y��(�	�I���!   ��  ��I�u ��F�K��y����E�0����U�  8�glL��տ�� +LMM9s�Z�ժ�?\Z�qe]H����C   �;(�  ��#I?�`�ͦu���8���I��Px�Z�_�Y�AB�����#  �#���ND_�ZU�Px�:����vIʎ�XG�
�@�1�  �!�  ��7� l�+q=���J���/�-,XEAU>�H��c  ��m_����+�1 `Y�����9���n�re]H�P�_Y�   @�Pp  p�_Z �qLpO�-��HRc��v�>SLo ��z��t���: �033�V�e#r�R�:���Аu��qe]H����X�   @�Pp  pϻ��Z� �1�L�riz�m-I�Eg�;�%h44���1  pJ:�Ӊo|C��ۭ� ��j��^k��[\��`�gd�:BW�a�@���:    ���;  ���� `c\�4�P*����u%IMI�|�:
b����F @W�R:����F>�Y�$ �,ݼy�:Fd�~͔����ct�+C#���u    tw   7��u  ��f\*��CGd�Jʋ�;�g��#  ��TJG~������$ ����37�o�W(XG0��	zά�����s�!   �]�  ��i� �ϥ͸�C��wjI��q�:����ŷ޲� ��i��?Ԟ�~�:	 �P�V��&���E�f�##����<�X��    �>
�   n
%1��!�6�z�d����i�j5�����^R�y�1  H����N|������i V�@7o޴�yN�:=�^�[G �q߱   ���  ��Z �~NMpwh��Ӛ��&''�u��̳�ZG   ���������g �2==�ԍ��
��d:=���ؚ���   ��  �g%��{ĔKӦ\����j6��������j�̨x����޽Gɚ����Ե���{����(�JDWHtEtEV�K$�I\�$q�Zf���4���ƃ"D.�@BPP�.CF��={�V}���>�\�սg�ww���>O�ޯ�zUwW��φ=�]������c  0�R)���������: �dkkK����1��ڲ�`ƥ��Kkj������  �1Y�    0�I���W[�{NMpw��.Iը���?k���8  �Q<^����ɗ��:
 �RZZZ���Q�#�Ѱ�a&;1a�o(���a�    ��w   �}�: ��qi3.��&덂z�j9yaaAA'BҔ?�Y�  ����.������=�� bmiiI��[�H���]��ڋKkj� Y���   ��w   �}DRU��c���qi3ΥM�Ea(�ZUnrRAhqqQgΜ�����uU���  ���N����?�cʎ�Y��;���T����^�^pg�;����$��  pw   ��%}Zҫ�� ؝v�m�o��n_{�Sp����-U�U�;��	vg�s�SĴF  �Y��9�x�+u�U�r�wS ��y�VVV�c$Jgs�:���C?�(���߭   �w   <$
�@b���S�v�_�\���Ғ�Ţr��Q"$��#�XG   ����:�������|�K�T�: ���Ғ� ���(��-��\���y�u {���&   8��;   >*�&i�:��c��;n<&=-,,����F��Q�����1  H�TJ�S�4��h���4�i�[�U�,[' �g}}]�z�:F�7��vJ*��ؘu��i6�� ��'$qD!  ��X�  @KҟJ�A�  �Υ͸�А2�����_�s�M�F��r����)�DH�ړO�[_�� @�;��ŋ��>_��-�_����u4 �g�VK����1�V��]�VʡS�\���   �w   H�E�H�6�r���J喟_]]�qr<    IDAT��Ȉ�����I���#�  0uS����T�xѩ	� ���E�u�D��kod'&�#�U���% ��%}�:   lQp  �$�����Q�  �̵͸�Ą��l�D�6��a�T*�J��}N���<��u  �"���;Ev .[YYq�b�^rz����u��rmMH�OH�C   �w   HRKҧ%��:�;sm3εib�
���n������'O�1�.
m}���1�!���׼F��E�/_V�TR֩  {�V��9ϟW��y_�����9e������Z������v��ރ.�ؚ�kkj@�=d    �(�  `�E��=��E�R��u��pm��Z���cssS###wl�n���
�M��0����O��Տ#�WsvV�+WԸrE�������vA ����#�tI�3gTܞ�^8}ZC'O*ŉ5 pK�NG�1��ܴ�`Ƶ�܁�ؐ�)�   �G�   ;>"�.i�:���P��ihh�:J_�v\������>fiiI�bQ�\��wկ|�:Bl�x����8��j��%_�t��C�S�g�e����Z|o-,P|��MN>;���yΝ�ޞ=�4�� ��DQ����RtO�(RP�Y�0��P
�@b|BR�:   �Qp  �����)��w{  [�vۙ�{nr�:��Z��H�ô� T*�t��yg������?n!�:��Ѯ���5���j��Ͻ���5?����33jLO�93���̮.> ��i�S��iN�V�̙g�?w��������h4�c$^P�)r��V�~6Sp��   �  p��w �Z���لtm��Z��+h4�����fSkkk:z�h��!���	��N|��+����s������p�_��U*�q��W�\}�93��	� \:�W��ћ
�ӧ5|�҅�uD x�FC����1�_�ZG0�w 1�&�S�!   �  p��J*K����\ڐ�:��z�N�rׂ�ԝ�722����>�B5�����1�R:�W�Ȏ�kt|\���u�;��枝�>?��������dH �q�)�ӧ�;t�:" 8-C-,,(�"�(��x�ݵ5��Ӏ�CI�u   �w   \�#��^k��!�wl��F~�*�:��ǖJ%]�tI�L�S!�jO>i!&��T<��k�s��S�oz�Z�R�m~���{kaA��$��ؘ�N����^<sF�3g4t�ҹ�uD �m,,,���X�~�b��K��u:�\t$��X   @|Pp  ��> 
�@��Tpwm�؍:���~���ZXX�ٳg0�����b��?�'�n)��k��E_�x�}Q�[Yy��~C	���2H �R����S��qN�����:qBC�|���a  񳱱�-~7�)��QΡ5��Ҁ�����!   �  p��)iY�q�  n��n[G�T>�L���эȽn��j5��eMMMP"�U����������1�,�Nw˧'NH/y�M����Z���KKj--�����Ғ���j--�S.�`%75���G�?vL��'5t�x��~�
'O*䈔N[� �X����ʊu���qx�{vxX)�Nm��$��K��C    >(�  �F��?����A ܚk�r��	g���l_YYQ�XT�X<�D���������_ٱ1�=�����ĄF_��[�z�������Zw|�����͙�F�Sثt.��Ą�G�*䈆�U��i�y�s'N(3<l �ga�T*)C�(���a�Lv|�:B_���$���    ^(�  �V~G܁�rmS.;1!-/[�0���q�Q�T*��ŋ�d2�
q�Zj/,X�0w仾�:��t>����*�>}��t��g'�_����-Ɨˊ|���w�s9e���9�};vLCǎu�[G ���ҒS'���_�ZG0������W���	�w��  �x��  �[���I筃 ��k�r�m�^k?wI�t:ZXX�ٳg{�qԸrE����iM��e�)b+75����m��KR�n�[[�:	~g����ښ�jU���qb8���NV߹͍�+�]^ڹ��a)��� H���U�q�v�sy��ck-���	�a�    �
�   ���H�)� n�ڦ\αM�k��Pd��jZ__�a&������̍�7:W�����]'�K�'�����.o}�[~/�孬toWW�)��˒�^ Qr���MN*�}�����������䧦�ʲ� 8X�fSˎ�f�/.Opwm�ŵ�4 a"I�  ��a   ��>Qpbɵ��].��w�����U�E�(�5;k��!���M�PP��Y�vBD�+����P�RQ�\VgsS~�rݭW._}?t��F:�SvlL��1e�ƔWv|���������S� 1�J��"N�90Q��ڲ�a&;>n��(������[�   @�Pp  ��<&�IIϳ�z�mʹ\p�k5E���)�Q�T*��ŋ�2iv`�WV�#��z�K�#�F��G�(�Ȯ�H�ju��ժ:ժ�jUA����[[�������s���e�o��Qe����)�o�w�~�X�� �=[XXP�ӱ�1��JEr���Z\[K��   O�n  �N��[� p=�&��vl�u�H~����Ծ���}�������J�R=��h//[G0���s�k=�.4t℆N���[-���F�[�o4���
�M����Z���A�!�VSP�)�<ͦ�fSa�s�¢�^?��� J���$e�ƔR�XTfdD��Q���ǣ�ʎ�(]((]((7>�t�ؽ�X��ٝ�9u ี�5�j5�ϯT�#�rm�ŵ�4 AI�  �x��  �;�o��/Ii�  ����)׎;Qgs�
��l6����cǎ�(��[]��`j�E/R*���cW������Z��u��ͦ"ߗ���-�7����$IQ��.�G�����A������h(
��;�����Q�l�����l̎�*���W��Ȉt�����2����(3<�T*���X�y�ƤT���LF�bQ�\N�|^�!�r9&� p ����֬c8���i��kk-���	���C    �(�  �Nf%}N�ˬ� x�k�r�M�Q��ʭ���X,jl����������������+�   ��T*)�"�(N�/��[ka�;[�   ��b'   ��� \ϵM���uS��*���(o{�0�_�(t�{F��<�   �=��H�RI��[Gq��x�=�X��y�ӑ ��K��u   �w   ���%5�C x�k�S��2Ţu3�,�A�R��0{����r|z�$�>�9�   �{����F��~��k��
J���1�ʵa@B|Lݒ;   pK�  p7[���:�g�Vp���c�Ů��M�V������>'�x���Le�Ǖ?v�:   �o�jU����1���w�X\\K�}�   o�  �,41�⦜kGg_� ��U*���?/�/�լ#�*^�`   طv����E�Nry���k,.��1�(��!   o�  �$i�:��v��(��c�����;j�}eeE5��у t|��p�u   `_� �����0���$
�n�����K�    ;   v×��! t�a�N�c��\<>{�Am�GQ���y�w Ϗ��m���(�   ��(R�T����(�_�Z�0��w v�c    �G�   ���  ����\v|�:��R�hb?�/p�{������    ���ʊ���ug��B߷�a&���k�h@�����e   �G�   �����[� ��vlj����vDA �V;��o��Z\\<����r�����    �I�RQ�\���4oc�:����u�������Y   @2Pp  �^|�: �.�6�rn�^���y��_�V���~�_#t�b�e
�   ���Z----Y�p�_�XG0��)yQ��<� �|I�  �d��  ��x��� ��Vpwm��F��%ieeE����:���Fi
�   H��5??�0��8����̵5�������H�(I   �
w   �ł��Z� @��5=�}���S�&t���4K[   ��(�����N�c�:�Op�MLXG諶�'�1��    Hv  �W� ���{nr�:��~�&��ZG06�   ��Z^^V�^���m���<�\"�l6�# �*K�}�   H
�   ثJڰ�ε�{*�Svx�:��~n���m�J%EQԷ���KYG0P  @�mllhc���8q���)�.�c�܁���$Ǐ"  �^Pp  �^�%��u�u��%){�u3��|��jZ]]������VL��O�   1�h4���l7p���spm��54 ��e    �B�   ��� ��\�>�����`�S���k���3e0���^�YG    n��<���s:V����"���
w �Fң�!   �,�  �_���u�eN��2��7�.����:�c���{ka�:   p� 477� ���:_̝wpm��;�c    �C�   ���� ���9��&���ӣ(R�Tr򂊤�
�L5gg�#    ��y�y�u�B�y
\S����x.��1ӑ�^�   H
�   دߒ�N`��±��h�Z-�F�Ah~~�Ƀ1�v��ޘ���    \gqq���b�������$-Y�   @�Pp  �~-K��u�U�f�:B����.�n�{����yEQd���z�ݯV�/�    >���T�T�c�:������ 
�X   @2Qp  ��x�u �U.Np�;�	{-�o�����i�,�us�˗�#    �V�Z]]�����~mm��	�.��1�,�#�!   �L�  p/�@҂u�E.N�rq�ص:�T�T���n�:~�:������    ǵZ-.N���i]<��54 F~W�o   �D�   �"��߭C .rqs.w萔JY�0���$����Z�Z�����#R���
w   �}_sss
��:
v�	��pq��P�;�C    ���  @/<��B%�>j6���.��*;:j�L\
�����8Je2�>l���W���2   �a���Y�>�i�"N���-S((](X��;�/ 3%�u   $w   ܫg�]��G�nι8ilG�6��0��ܜ<ϳ�ICǎYG0�om�q�u   8&�"��ϫ�n[G�x1zm�o���4����e    �F�   ��n� �k\-����`&NwI
�@sssL*����#�   ����E��u��#?f���)75e���kh��uIY�   @�Qp  @/���5��K<�S�1���icR�
�R����ܜ�0���<w����   ����U*�؇8���W�TZ��u�EI��G   �
�   腎�Z� \��]���XI�lnJQd�&�VK�RIQ���p�usտ�k��   �Z__���}�M�u3���;�    �(�  �W~C�F��\<b��{��ȯլc�R�V��Ғug_�d�^�����)   0�j������c`�:�uS����u�5_���u   $w   ��W%=jp����ԔuSq>J}ssSkkk�1�4r���ba�ӟ��   ��l69�*�:���L�84 �"����m�    �  �K��: ��Xvu�؎8�%iuuU��,�Uvb�:���Gq��  ���y������u��'�:d��Z�� �U��~�   �  �K���N�G.Npwq3�ZI،_ZZ��֖u��w�usa���?�S�   0AhnnNAXG�=��E��š.����T�  ��@�   �Ԗ�A��+\ܤ�NN*�v��l�SGQ���'�}Z��~�����OXG   � 	�Psss�<�:
z��;w ��   08�m   ࠼M�5}��&]*�Vft�:��$Lp��%���yJ }D��k�_Usv�:   @E���w���r���)�.�c�]�Ѱ� ���l   ���;   z�	I�X� \��&{��!�f�m������Yu:�(N��-����Y�   � X\\T�^���r�����vIj�Z� ���u    
�   8,d}��&]�Ⴛ����N����Y��oe��<�yJ���1ba�U��>   ܃��EU*��$]4�kYG�R\X���   ,�  p��bt�ݓ��x��477�0���t>���?�:F,��V�����  ��ZYY���u�Z���E���G��ߕ�Y�   �`��  ��Б�;�!�A��&��w�VS��X�سV����yJ�l��/��=$E�u   $L�\����u�����k��Ąu���}Jz�:   w   ��J�C ���M���u;Q$?�����J��"J�f���#�F�����_Z�   @�T*-//[��I�k�^a�;���.[�   ���  ��2+�ϬC ���hXG0�u��.��ذ��o�ZM����1���^�T���s�~�u   $����U�W.[G0��ZJ�ղ� ���   0���  �Aba8@�n��ݔݑ�M�J����%�);6��K��c���׾��/~�:   b�Ӧܐ��{!��wW�΀>Z���   L�  p�>��$w ��M�����;�ؔ�����ښu��4��[G���w��:  @|E��JE�R���� �V�N�W�fS����0���Enb�:�	WO?��%��!   0���   0�BI����A�A�l6�#��ML(�N+
C�(&:���zbuuU�tZSSS�Q��K_��}�:FlT{L�<�C����Q   ����_��jO=���O�1=�������[>>=4��'T8sFc/x�F��|M���ʎ��9��j�ۚ��S��kK���Zz�\������'��_�  ��E�   ��%����u`�8;�*�RnrR^�l��� ������N�599ie`L~�*��+�<�(�1����|�K�Js�!  |��5._V�T{�)՟zJ�RI�Ä��VsfF͙m<��$)��j�4����}��*����=���쬂 ���>����)�.�c�����JZ�  ��E�   m]�H�Q� ��i�Z�̸\p�ئ���$Qr�L��ɗ�D�G�������'?�c��}�Q   z&���x�iշ���˗ո|Y~�v _/�}m~�K��җ4������_�ӯy�ƾ���$��433#������\]C���R��kg@��:    w   �ïIz���u`�A�N��\.g��o�Z�]�����N�5>>ne z��(���7�I���[��~�w_����U<{V�L�:  �텡��W��7�~Z��]���=Me�i$���>��O}J�^�2������^`�e�:��fgg)�;��ܴ�`��5&��˒��:   w   �×%=*�[�� ���l:Yp�:d�Lgc�[dI�5CQia�{�1%�{w�;�SO��-�1b%
C5��Ԝ����Ϯ~>�ͪx/]�ȥKy��4r�}*�:5P�� �d�U5�\Q��5�\Q�'T���S�	�?��Gѱ��^]�������r{�ӱ��>�<O~�n�L~j�:��F�aT�a    ���;   ���E��f��d!8Υ��v:
�ueFG����N�=�Jill�:N��:��K�Ըr�:J�E���v�l��g�ǻS�/]��s�������}�)˿M  ��rY�+WԜ���.2=���������'���Oh���s��&��o�Nt��577'����7�'��Evb�:��V�/�,�}�!   0�(�  �_> �%��W�Z�;<�]�n���.uK�RIgΜ�� ���i�;����=�UU{L�����CǏ�xႆ/^�ȥKW�w�T	  p{���n���g�}�rE~�j�@t�e��O��μ�u��?�T&cI��fgg�n����H�񂻫�W<�S�1�A�I\=  �G�   ��;��笃 ��Ղ����;:岊g�Z�8Qi~~���=:��߭��1L�����jo�+    IDAT//k�_���ى	_�x�[��N��R)��  �/�P�RI����+W�|�5��4���/�4����~����+��L�h'���Pnw\bOG�WO�su�8`���Y�   �(�  ���*�g$孃 ��գ���ܽߜߙ�~��Y[�I���@�s�Ԝ�����RQ�+_Q�+_���b�;���/^����tI�3g�ʲ, @����Z���McoNO�1=��������뫯�����լ\�!��!��{nj�:�	
�������   p;i   �%I��j� ��pu�.�������u������(�߃c�x�f��N�N�M՞xB�'����lVųg�+�o�Ӆ�QZ   IA���5E�����O?�V��(��%��׾�����Z/���Pfd��_{����E�ޠ_$~7C�����f��Z   �;(�  ����(�=��f]fdD��!�N�se�\�����ٳgU,��$����
�1�����u���R:vL�s�T<{V��g�E�s�T8sF�<��  ���5?�����o33�����jO<����O���v�����5w��^��\�H��R)e�NQ��.@�=)�O�C   ��  �o%�I�f� � py�>75�`q�:�	�J7Ahvv�I��P<^��{�jO>i�Ej//�����G�������/^��}��p��շ��� �-x���)���j�Jj�Jj\��������Qy�1}��o�s��kQnǭ���F��q�r9�&�> ��ۭ   �-�  `�m��k.o�妦�r�����ajnnNgΜ��Ȉu�D9�=�C�}��ժ��?���_G:��M|߹:uJiG-  ���KK���|�vnN�����z�uBl[��'4��:��;ԏr;n���a�Lnj�:�� =U���   pw   X���7K:cH:��[�>l���X�]�U���)��ѱW�B�>�(��� ��Zj-,h�_���tZ��'������N)�ey o��U*�97�l�}������ӱ��]z�WU���*�?����@333j��=n$[�騳�e�L��!�f��u`��[�Q  ����  �_һ$��8�x.�so҆���VSft�:J_�Lr?}����Ƭ�$B��QM}�wj����:
���Z��Z��6>����Je2*�:��ٳ:sF�ӧ5t���۬c�c  v������ו�WV�(���=O_��_�7��o*�N��y}����,�v�Rgc���!9����f���   @_Qp  ���J�YI�����-�<�]�Nq/:X>��H�R����|��)�㖢 PsnN͹�[ޟ���Zv/�:����ݷS�4t�ҹ\� �*h6�^\�z������E5K%���uD�I��_��G?��zUO��r;���Ю��p 
�@����y�   pw   Xٔ�AI��u �\>n��MZI���U<w�:������S�4>>n'�&_�RN�Tkq�:
ƯT�U�h�o����R��G�^-�_[|:qBCǎ)�e� \�ZW���ś�읍눈��w�SǾ�������t:�����y=J�A�Y_��`*?5e���C!��5�    p�L   ���%��zw.5���Q�|̶$u�BE�E�&&&���Z*�։�AM���Q0@�0T{yY��eU{�����9��ɓ����:qB���ɓ��� ؗ��P{iI�[Naw}B2��[]��C���^���܎�r��S�Ⴛ�C!�zDң�!   �&
�   ��w��L�wY���iT.O!�(�Kݒ���TrJ�wv�~@3�|�� ��W����y++�>��-����Zx/�<�����	��Ç�T����=a�}��%oeE������r����"�V���S��t�5��׉/��inn�r;v����y�O�sy�衷Z   ��(�  ��w`�\���Q:�W�h��s����Nr�����[��Gu��/�ڧ?m�ʯTT�TT{��[ޟ��?rD�c�4t���G�>[~�~?��R�L��@rD����G�׽��n�}eE���p������|FG��?�۟�<������J�A�|�����\^3zdF҇�C   �]�  `���Nr�u �\?n9?5��Ғuܯ����05��d�;9��?J��v:j-.��}R�-��:rDCǏ+w��
Ǐ+������S�������>�Uykkݷ�իﷶ'�����)���uT��?��=�[��fggp*�������Q�r9�f��ܳwH�I   ���  �8x��_�$Q��VEJ�R�QL�.��>��V�����=j%��_�B�������_[Gz'�^YQ{e�K���=ڝ�};t����G��Sp ���ݾ����)�_Sbo//+�׭�����cj�̨x��]�h44??O�{�r�=���܁{R���Y�   ��(�   �%�?H:iH�(��j�T,���py����!E��������� t��	�(�t浯����k����*��*�����𰆎Snj�[|?|���#G�o�+;1ѧ� F���Pgc�[T__W{eE��uy��j����]^=�:-�7���.��O��1�ZM�RI!�`��NG���^3�(���=���C   �m�  ��ߒ��� I�r����ڰ�QgkK��q�(�����0u��IgO7���/�
gΨ5?o����PczZ����c����9��ؘ���W'�g�Ʈ��WvlLyN� R�n˯V�NY�����W��?�VW���P��i�&+��.���R:}���ժEQ��ax������P ��;p<I��:   @�   q��J�I��A��i6�:t�u�Ç�#����)��F�RQ:}��ҷ)�8)����=���X'ϯV�W��zl�PP��!�V��!�&'�S�VnrR��I�''���辍�+1`!h6�)�孯���)sS�5�������:�:�ln*�}��@�WV��裚��o�龍�---� �66�#�rz(@��D`�~_Ҭu   ��;   �bC��J�	� @Ҹ<�*�h��W.�x�u�ت�j���י3g(�_��+_��w�[^�lpF�j���������d��)���+;1�����s;����n9~|\�B��&@�Ea�`kK�JE~�����(7����!E8�����M���u���% ����w��ʀ{Ib*   b��;   ��%���r�A�$i4�̸>�������u����ܹs�d2�qb!](��k_�g��6�( n#
y��ϧ��n*�gGG��ގ�<{;>~���ϧ���o�M��
�[[���Bzp�b��ǝJE�֖��-�� �h�/�BA����$ieeE���Ʃ0ڎ�;r����Zp�>#���!    ��;   �eF��$��:�$�V�:�����;�o��V����̌Ξ=�\�k�$��?�������ܴ����v[���9�6��>[�S��b��%��Ȉr��J���
ݒ�А҅�������=��!�fSa�y]1=h44��k5������f�[X�yL���^�_�)l6��8&h6�����x�������葎���\pg�;�o��u    `w   ��/I�AI)� @R��u�f���J��Ζ���{�v��$�|>o�\fxX�_�ZM?��u 1��:��=��%32�-��ʎ�t�����+��w�
J=�~>��ؘ$]�X��������J�rR:���H��+�e��&a(�V����������n����z����uEA����NSo6v:
[-����^�ZV�)�+�,�� n������ߨ-Na@�^p�;<�	���|Uҧ�C    ;X�  @�|I�Ò��:�NO�J����Rki�:�	&��M������Ξ=�"��u�~H����J�:
�����t��2e�-�g2Je��KR��N_}|�PP�6=��������rJ��=�)�� �)�_�qp��W�;v:
�)�G���R�	%]���u���Ջ��^�~͜���+	��Z��f    �w   �ѯ��;�k�O�ʹ\p�ذ��8AhvvV�O����4`We��u�u��3o�u �(�W��t� o��5I^h�_����n�H .Op�NMYG0��i��>�$��u   �Z�?   軏Jz�:���>r�+��(���8aj~~^����Q̝�������1   ࠎ�I��Ǜ���a���;��5y��Lp���%��!   �kQp  @\�� @R��i�?|�:��(ԩT�c$REZ\\��ʊuS�|^�~�ǭc   �1mI���IW{�)y��F�0h<���Kn��H� ���n�   �
�   ��ߖ4kH׏]�9>����n!���׵�����I�ǿ��5|�u   8�)iMRp�Q����G<�_+g>�N����oJ�Z�    nD�   q�Kz�u 	\���z���M�^�T*���S��QL�2]x��c   �5u���͛�;z����C���Ppv�.�-�!   �[��  �8{P�}O w���]��M[o�o��P��533#�����8��k�[��:   XE��]Ӝ�U�T�G8��Lpw{�؃��=   �w   �YK��1��/�;�i�K�VK333�<�:���~�g��f�c   `�D��%Uw���/~� ���/�>l���ke�.y�~�:   p;�  w�&i�:g�z�:�������u3�o����y���vr3|��%�����  �JZ���YʕG=�4p����>���2`�>$i�:   p;�  w��k��f��(��c�I��w���6���@333�Vw;crp����P��Q�    ��I�=���ܜZ���.�8\p�
���1L�x�:�G���  ����  �$�e�}?pF��<�:���Ó�\޴?HQ�T*iuu�:J_e��u����   H������>�<S�qO�H^�l����%���˹��>.�k�!   �;��  �$X���u �\߸�;�y���
[-�kmmM�RIaZG�c�x�&�雬c    ���$���_�b���E�֖B��>�n���d�.0�   �G�   I�K���Q`���q�?|�:�)�)��Z�jvvVA�ȏ�TJ����)��Z'  @�T$�K���C33j//� \䭭YG0�?r�:�)��������	.�s�!   ����  ���;Il�+��o޺�y��fS�����8|�N��Y�   @BD�۫=|�ʣ������/�9>��52`~�:    ��  �$?�{�f�i���޼���4==�Z�f�/ο�*�=k   1HZ���J�&w�����FB���/J��   �nPp  @�|E�'�C q������:�o��S���W�\��r�2Ţ�ޛޤT��#   �ZGҊ��<w��y����t�/w��;ׇ@ w�    ��%   ����=��5\߼s}:��+�"-//kqqQQ4�?��_�"�����  �j�[n��k0���w��H\���>f   �-
�   H�/J��u n\߼K
ʎ�X�0��潕��M���+C�(��ߨ�s�1   #[��$�o�
���/O�����Na��52���  �D��  �$��b�;p6卵������j5=��3j���QL�P��{ӛ�4�H   ��$�%m�?3���V��2����s��J�r�1L�~�!p+��C    {��$   ��Ie�6嵐�G�#��ln*
���<O333��ڲ�r`�_�B�}��c   �P iUR��_4����c���H�����j�1����G����R@R��  ����  ��z�u  Nؼs{���P�r�:�ӂ ����VVV����ox��x�:   �%-o��[��;����rG�XG0��&�%=d   �+
�   H��H��u .ؼ��o�z��� i}}]sss
��:Jϥ2=��~I��I�(   裺��ۭΌ�=�^�b�:��6r|mD���u n�,i��   0�(�   �~�: l�Qp�8>�.Nj������y�u���;����Je2�Q   p�"I�����m���&@�x��6�:d�C ��\��>�   �~Pp  @�}L�Tb�N��[G0��xi�ۚ��V�^���s���mzο���1   p�u��׬�l�<��v����9�/��4��Á{�1�   	E�   I��� q���]�RGAhnnN�r�:J��+u��~�:   @[���m\T\�,��#)\/�9~���Ӓ�e   �/
�   H��H��u��wRvlL�|�:��7��*�"-//kaaAa8X�.���s��_Z�   @�՝�X������׿n	����Lp���u .��$�:   �_�  0���Z-E�O�K�����Na��M���T*���V��9�����_�ox��JYG  �=�$mH*o�G�����p���t>���us�IҌ�w[�    �w   �?���u�R�j�Z�1��>��[_�\��!���fffT�V������/��_���(   �_Ҳ��u���|���wQ�N�l��L��.>w`ۛ%u�C    ���;   �/X �����������ڲ����@�RI���u���.=�ۿ���﷎  �=h�[nOB������u�XgsSQX�0�s�T�k�>芘�  �@�   ��c��h����wx��$uVW�#`�6775==�N'	U��y�s���ާ3���Ki��   �,�T��&)4βU���<�_9|���v��0L�w5�@�Y���   ���   $Lq�Ӛͦus.Op�����I�j���3Ϩ^�[G�t>��?�S��~P�^�2�8   ��@Ҫ��u�}�Pp��^pg�;� I�%��:   ��  0H>.���a�T�ݯ��w�7�(���jee�:JO_��ox�[�>��o��8   �֖��}�D�'�T�k_�F{�^W���K�I�(��  `@Pp  �������<H������O����s�G�"=<Z���UQ�.�D(R'T�
��ǔd���� q�;��f3�8)(pT�NcS(R�yĳ���Ν����}��>�䏞陹w�ޙ{g���������<��w���s�?�&��7��upp�����}�Q���>������}���Z��oQ�T2	   �ZLn�My
a���˦c`Dy���F%ggMG0��;"�MI�b:   pU(�  `����ϛ��"����V̊�[ݨO�w�mkmmm"OV)��z�����������~�r�=g:  @$�*��B�Y�B�K_2#ʉ�I�)
��~����  0A�    ��G%}�t঱�'�	%�e�ժ�(F0�}�y����u���kv�	V*��~P���$�=8P��W�~�55_yE�k�E��/  �u�I�J��}�Z/�,�������E�=q̲���1�8�? �^��  0a(�  `���?��u�� 7�E����ld���E�	�����d۶n߾�Dbrߤfg5�u_���;�����Q��W�~�U�^}U�oȫ��  ?�����&cj�I}ۖ��ʿ���(!���c��(�K&M�0���������  ����R   D�'4(���DdPpH��J_���F��/�Z�7�سm[+++�}��
���87&����Ғ���_��o6�YYQ���~�5uVW�Y^V��  �&_ҁ��'U�O���;N�� 0Ø�$�G�eI�e:   p�(�  `R�{I�����
�Q_����Sp� ��kssS333ZXXP,�����J�{�J�{���WwcC��^�����ʊگ��   $�+��A�}����e雿�t������F���LG	LpGD}RLo  ���  �I�II�d��
�Q/w������n:�X�ZU��ѝ;w�J�L�	�DB�^P�N���﫳�*{yY��^S����Y[��4G  0�BI�4�H    IDATI-�AnH{yY�m+�ϛ����홎`T�O�?±1D�$���   �u��  �I�ǒ~G�_6�	L�HG|jY/����q���iiiI�R�t�����Wj~^���x����,�+_�����ʊ:��r&  x�X"��[�28�������j�w~��s��$�Fj��ʩ�|�6�R1�������;"�M    �w   L��􍒒�� ׍E��d��nķe�t��kkkK�v[KKK�,6)��x6��߭��}��~�%��=uVVd����++r��%  Qu�Ȟ�sG�Ýjro}��;�8��*�ے꒢�WM��_����������qLG n��ux   &w   L��H���K�A��F�} E��t܀F�!�qt��me2�q�V�XT��P��8u�W�����Y]UguU^�f()  ��\N��S���%��W��畽sG��ɋ��w�}�Y���I�����/����E|�;��v�m:pSBI�4   �N�  ���W$�M��mۦ#��x6�D.�~D�=
����������Y���)���41���*�ר�5_s��~�9,�w��e���������� �sS �y�ҰȞ{���4��S��-�)_��>�����EYǕ[�ʹ_�۷MG�p�>�}~�t����1D��J���   �u��  �(ؐ�����t�:��+��L&MG1.97��Ɔ�Fx��B�S��"!CU*ٶ�۷o+�J��4���J�}�J�}��ϓ��'{yY�������Uu���w��� ��K$�^\T�ΝA�����{W�;w��s�ʿ_�T*j��B���GZ��B�
z=�[-�1��g2���c�
@ҏ�   \7
�   ��OI����� �u�v��%�ԍh�]a�^�2����v�Z[[�����8�c%��E�~px�mo���������KowW
C�� �E�,K�%e�yF�g�U��g�}�[�{�Y�������8��߿�^���K/Ezת�گ���}�t�V*�~m�ZX0adt�w��I��!   ��F�   Qq_�/H��� �ɶm�J%�1�K�͙�`���O�=�|�������nݺ�x<n:R��,����_{���;[[�޻'gkK�֖��  DW�T���Nc�ܹ��s�)������ժ���xc��y�j����\����k
�P�X�t��홎`T:��@�x�'�uM� ��+�GL�    nw   D�ߖ�m�fM�[1D}zY/��Q�j���tt��-�E�qp��KR��TwsS��uu���ln'��L$ ��ųYe��N`ϼ�-�>��r�>���(�y��߿�D��������m�Y_W���LG�A�J�t���%1���K��4   �	�  %MI�Pҏ�\��>����7����{��ijjJKKK�,�t$\B�TR�]�R�]�z�1�Z�s��`���k��=�ժ��  ��XL��ye���Hvt�޽��̌��h4���+���|����*fY
������֫�Rp�87�����#��> ��   "��;   ��'%}����� ׁż�T�w{_�ǱF��N��۷o+�˙��+���QrfFů��\W������A�}kK��uVV���QxNA �qb�RJ��K�J��=�x6k:�S�}_���j�Z�|^�XT����YY��d����+Z��o0���,��@�pL�ӒvM�    n
w   DMO�/�gM��yQ_܍��:��y�666433���9��O0+��������~_���CSߝ���ܿ/�� �Q1AS�/��ji{{�ܩ�*��=�%�o������MG�!Q?�;��@���!&ܾ�   @dPp  @}Z�Hz�� �Uc1o�J��,��5���A�
�Pj�Z�u���#(�H(��3�>��x��l���Vo{[���������Y  .#��>T\O}|���T�t����vww�h4.�y���j���o_S���;�:++ʿ���(0īTLG0*57g:�H`�&�ߓ�6   �I�  E���-�L��y�Rss�-��m[~��8%f<�u]����\.kqq�i�J�J*�J*��ҙ����JE���`�������ˍx� pZ�TRjnN���S��SssJ��+s�����9�ͦvvv.<�����ަD.�>':�����#ʷ�H�H���?�11L�5I?c:   p�(�   ����?���A���bޱ���1�q���}�Y�10����:���qaV:=,'������m[����)��﫷���ޞz�����ȭT>Aq 0�,K��y�o�R��me���^ZRjiI�����L�tʑ��������S��,��.տ��+L6�گ���o�&�1`���g:�Q��Y�F�b���$�t   �Qp  @�����[c�01X�;�-�{{{��HLs�U���ʿ����S�@�����m�������}9��rwvԫT� ��� ��,K��Ye�����WfqqP^��W���ܜb��c�i��?����Pp��y�M�a�;DN/�;	���MG}��zYү�   �@�   Q��H�}I_o:pUX�;���"��E~\\�^�mۺu�����8�T�����c�m�7�r����ߗ[���ڒ{�vog�I� ���2w�(57�����v��vzqQ�KG��*��?����\��g�NG�榲oy��(�aQ���c'qLꓒB�!    8J	  ���!IQ��0X�;�)f����#��icc�i�0.Q*�P*���w��x��r+�vw��j��jU��=y��p �ZU�4x �,%�����UzaaXX?*���攜�Sjv����j5���_����Rss�ܾ-���+������?��AQ?����1v5�����3   0��;   ��O4���#�� W�żcQ_��E|����4���%
�q����q��^\|��@����rXzw��O���]�k5�w3���,��'>N��S\q��jgg�ZOF.����%��xCs����aQ����Ob�&L 飦C    &Qp   ���W$�M��y�R���YVd'�2�O��<mnn�P(hiiI�d�t$��,kP�������G>իՆ�w��@n�"�RL�?8�W��S�K������Ai}zz0Y}zZ�����rY��Y%gg�ω����
�p8�=����w�S����~�q`���0 �ܓss�#���a����?6   0��;    mK�I7xZ��(C�b1�Q��%�J��r�U�Q�p+)%�_�j��Z]]��ܜ����w�D�{�[�ܣ��W��_��wp�~�.��c
�@4%����%�SSJ����J����GL�N�����z��~���]�����q�U������+R�0�'w�)�Qp��H���   �i�  ����I�L�F�v���r������\d���k4�,�MG��}_���j4�u�2���H�Q�r���?��a8(�?�_���j��l*��"$���s9%���8,�/SSJ���"�Q�=Y.+��������U��� �|^�瞓��r��w�o�A�=B�z]�癎aL"���͚�12:����U�I��C    �Qp   lI?���c`�ٶM��Pj~^��6���>w\	�q������i���˲,ӑ���]����I�fspi��5�[-y������u��~���u���G̲/�,��׉b����ǉbQ���aQ=Y.�J�L�ǘj����ّg�l[x�;(�K���5��_k:n�[���`'s�P�㘎\�=I?n:   0
(�   �~N�#�]�� Oömͳ�)������r/�h:&D��V�j��Z\\T�P0	�8V*��ܜRss����qN�O���}�VK~�#���]�ݮ|&^b�X�⹜⹜���٬���`��ai=Q*)yXZO�J����|��q]W;;;�m�h��;ߩ���=�FAgy�t� wo�t��~��$۶����U�1I-�!   �Q@�   8H����5xl�|,��^w�tL �u����B����%%�Iӑ H�2�3iaቿƃ��~�5�}���q�s\��v���o6�?�۽�.��)�H(Q,�J&ee�ǥ�lV�BA�BaXZ��r���y%�yY٬���9��b��	x�0U�մ��� L�Qᥗd%
�}�Q��nn*�<�x�	�����1��L�d\�?����C    ���;   p��I���?o6��X�;���bo/���p���VWW5??���i�q \�D�(�W�������W�ݖ�`�q�8
\W���w����}_�mKa(��|�VKaʷm��?�\�S��)��z�|�Q��Gz��J��d�3Y���D� Y��nK�%��g���s9�D9=~XN?�/�HJ�鴬TjP@O$�(N}O J:��vvv���LG��i�^xA�7�0Ũ�����T�LG���I�O��Ϥb�&��5�   @�  �����/Jbl ��z�2_�u+�0�|���Ύ������LG0B���ҍ�0��xI�������Q�~xG8(�? �<��D�=���g��R�?��dΝ:|4%]:<AR,W<��pF O��}U*U�U�Q�Tx�;#_p�${y��{DD�=/�c{�����6   %�  ���I�%�æ� O�E�c��Y�,Ka��GQ�f���8����555���%r`N̲*֟]��	�P�ZM�JE�s��K/��0:++�#���ߵ,��`:���X�\ �c�C    ��2    Q���G`��w,fYJ�Κ�a�{p�p�8�<�FC������W���   <�N����U���t�]��o{�bKܣ!�#���M�����!�ܯI��L�    FG�   ��ݗ���<	�NKFx��0ԏ��?n^�T*Z]]�  0�����߿���u�z=�q.��d�}�Y�1�s����x�y�ݭM����L�t���n3�c˖�I�!   �QD�   8ߏKZ7�,
�����MG0ʉ���0���iccC����<�t  �	�P�jU���j4��\ZᥗLG0/���0�׬�������=`��O��   �"
�   ��z�~�t�(���^\4�(w�tD\����ʊ���Dx�"  }G�[vww��uK᫾�t�����4�,��u��#�
�S�����   ����   <گH�C�!��`Q�T�'�G}��!U*����u<  9��w�q]�t���g��$ɡ�>�܈Op��~�31�~H�c:   0�(�   �����st"���iQ����옎 �����Mmll�qX�  f�����=���L�NX�RI��%�1��nl���k��`��8�1�G�~�t   `�Qp   ����[�C �ԪӢ��ۣ��d۶VWW���%��L�  ���ժ���upp�0MG�R���*��s��&���E��n2��=��;�L �L�    Fw   �b>*��0��z��%r9�1�q��$�Q�fS+++���S�Y
  �~�v[+++��ݕ����\����f:�q���abE��7�'�?�a3�*鋦C    ���;   p1�%����E��}��k:�HIEx���8�M�1�sA���-//�^�3i  \�n����umnnN����[�j:�H�nn���k�5��tcb�R���c�۶MG .�%��C    。;   pq?.���E��wZjq�t���]������������;Q  �+�y����"�#s���T�t�(�O����M��K���##Cu�]�1����%�   �
�   ��9�~�t�"�Rܸ��o�݋��?Ƌ�8Z__��Ɔz���8  `LA���}������b��ܳϚ�a�s��*��q��K�Y�Q�c �.��   �
�   �����k:�8�OKQp7�4۶��������}�q  ���P�jUo���*�JdK���7�8w�����?ۨ�x�b�|T�!:    . a:    0��O�Kb�o��v�m:�Ha�;w��0U���h4T.�577�x<n:  Q�fS���r]�t��/��}�!���Ja(�b�������LG0*��8Đ��ߗ�/M�    �	�  ��{E�?5x�N�D|�;�]�I�{{{���
  �f۶VVV���E��P�LG0����5�c�D�=nj~�t���w�W��   �
�   �����aha�OK��*��n��19� �����|�MPt  �l����666���L�)��%ųY�1���옎�k���Lp?�c`?���    �@�   x2uI�t�<�v�t���,�fgM�0����j��\����������u�ah:  �A�nW��ؐ�8�㌤X,��3Ϙ�a\oo�t\1��T?�f
8ށѶ#�S�C    ㈂;   ��~V�M� �B��a��E��br!&��y�����ꪚͦ�8  �������-���ɶm�qF^��]������I�E��4Q,�bw�S�}��	I��   <
�   ��%����A�����T�'��L.���z��  �`������Z^^椶K��.�"^��DQ�3M�ϛ�0rx��EI��t   `\%L    ��J�MI68�Ž�E}���wD@����Ɔ�٬���T(LG  O�u]��h(C�q�N��{��Гȉ���Q?y�,È�%}�Cr    <
�   �����o�T28����R�r�wDI����榲٬�����MG  �ຮ*����&����wɭVMG��E���4����m������/�   �3�t    `lK�	�!��X�{X���^@4Mt_[[��E  ƀ뺺��VVV��~Ţ�h����
��t\��O������^#�@��4   w�  ���^68���E}8�% D��D���5�M�q  �(�_��3Ϙ�`T���o��o������Pp��[��   <
�   ��$}��5`\�ݦ� +����¾m�g�������E� �A���en�2��~�a:���n������#��<`�|QҧM�    &w   ���;I�a: IA�q�1FNfq�t��������j�L�  r�~///Sl�f��Y����u�pE���6��w��1B|I�'�6   ���   \��T3�آ�,��o��2 �n��{��iyyY�jUA�F,  \�N����MvS�Aɹ9��c����{�������1R|�W��38�iI_0   ��  ���'��H�ϒ��w'�e �<��jwwW�����ߧ� �k��Z[[���:�SnX���\&�O��ܣ~��Yl�f��I�0   �$	�   �	��J�vI�3����,-��`��2 �8�~_�JE�ZMSSS���U"��3  �D�j6�:88`��A�%��&F����8'Ma���$~�    W�:   �ꅒ�[�I�΂c��aܣ] .��}U�U�j5�J%���)�J�� �X�@�z]�jU�癎yɩ)Yɤ��Y�k:�H���F���Y���$���   ����   \�/J�eI�a:��E���MG0ʉx ��0�h4�h4T(4??�L&c:  #��	b��#��R33�~/@�}rD��c�cga�F�+��L�    &w   ��|L�7Ib?pA��a�\N�bQ�V�t#���|�V<�7;�v[�v[�BA333���  I�뺪V�j4
��t�����
���t"�^��F�#�%}�t   `Qp   �OU�'$�c�AM�ϖ^Z���xooO��7[GE�t:����J%Y�e:  7ζmU�Uʅc �h�^�t\7���c�s��xǾ`غ�O�   L*V�   ���O$}�tDE��E}�Y/� ��z=moo��7����<�3	 �k����VVV����{�1��;��&���c:�Q��y�8��!�a�_��1   �TLp   ��wKzYR�tD�|gKG����w�U�}_�jU�ZM�bQ333�f�� �-�    IDAT�,�~_�ZM�ZM��K�"��$t]�p�~�vԏe��c_0���;�C    ���;   p�ޔ�S�~�tD�|gK-.��`Tԧ��%C5�M5�Me2��̨T*)��� �sG�jU�fSa���'�x��	����3��tďe���D`HC��   L:
�   �����o���� ��Ζ��Գ����T*J/..KK��Y���x�DpG�������fff455�x<n:  ��Z��j��:���8��d�t�b�e:.!�<9;;������UowW�Ύ����������p�)I�M�    &w   �fx��Wҿ���*n�|gK/.J���	�~���믫���=�,�.�^(���y�vww����b��r��|>o:  g���j4��j�x=Q�5�(+�6=O��=�vv�;,���J�Zd߯?J�O�?�`�%���   @Pp   n��$���΁�`��lV&��Ԕ�z�t�������u����z,��+�������J-,({�2�<�x6k -0>�0T��T��T:�V�\V�\��4Q ��m[�z]�VK!�҉8��F%J%�")�}y��Ⱦ�'woO�֖��-�*)LG+��Ʊ/�0O��H�   p(�   7�I���9�A0�<ϓ�J�R�������K�۶���ꜱ-|�T:������2��J--Q~�������J��b������*
 �aG�����܈O����OpONO��0��nW��}����"{��{p@���X���sJ<�����/�   Dw   �fU%�-I?o:���m
�g�,-����cL�ٔ�l���=�(�e���A�}~~8	>Y.K���Āy��^��^�+��hzzZ�R��� �k�8�j���ͦ����o4LG0*}��cͫՆ؏�ݽ=9{{�7���EBja���g�P�n�tDǺ�5   �
�   �����o�����`��mM3��!��E�"��l��lJ_��C�Y���33J���������J��LZDd8����m���\.�\.sr ����?�����Lǁ��=���=���#-�}y��p��Ⱦ�����|�11�2KK�#�$۶9Y7%�`g֎�    @�Pp   ��.�3͘���n�MGI)�GB��K�W^y��D.�ԉ�{rnN��E%�畞�S,�4��>�����@��r*��*�Lu \Z��t:���j�Z
��t$���(Op�,e�y�t
�����JePZ��=���S�Z�(	����#�c^�A�R��   Dw   ���%���>e:&�}gc��x�w:꯯�����������`���|j~~0~fF1�p��t:�t:�,K�BA�rY�|�t, ���<O�fS�ZM�癎����H>�!��$+�6�������^�ȫT�;*���˫T��>�R�Bw&۶MG@4�%���   @Qp   ��1I�"�ݦ�`ru:�{���b���)u�+��j�j5�7z8�+5;;(�/.*Y.+Q.+����Rssx�� �l6�l6�N�U,U.��d �� �n�U��)��!�3^+GI��MG���ɫׇ;`�G���rww���D�ܺe:�H�wn�J�1   �"
�   �9}IU����&Lp?[,�TrzZ����(�&����W^y��x&sj�{jaA�9�������H<Z��S��S�RQ>���Ԕ�Ţ,�2 `��8��jj�Z�}�t���W�b:�Q��^2�B|ۖ{p0(�N^w+��e_~�k:"J/,��0�8��9I��p    �(�    f}Aҧ%}�� �LLp?_zi��{�����Ɔ�g>��畜�Ujn��r�qrvVɩ�N�f۶l�V<��ԔJ���٬�X �k�y�����\�5�.�~�u�)���{�ՒW��*��'J�L`�y�dr��w\3[�w�   Dw   ���I�O$�`:&ӬΗ^\<s�7 I}�V߶�-�[ɤR���%��Y���'��Kp����}U�UU�U%�I�J%��e�R)��  W��}��m5�|���ښ�j�tc��R70�:�v�V���ZM^�2���pB
�Pj~^��L�I��5���5�!   �(c�   0ϑ��$��$V�p�X�;_fi�t����������9��e)Y.'���ӳ�J��)53�x>é1�<������N�U,U.��L&MG \R�J�a���1T���MG0*��sO�5B��֫U��U�*y���JE�Z���Vi�]����p�� ��   Dw   `4���~C҇M�da��|)�q�� �[�>rbf<�VrvVə�gf�����%5;++���Ԙ$�^O�^O�JE�\N�bQSSS��㦣 ���:����Z��� 0	�,)�?�����Zm8e�;|��V*���f�f��H/.��0��k�J�I�]   F�   �/�/J����,���)h0����߿/��}��yN"�S�잚�Urzz8>ux���x�N��N����=��y�J%�EY�e: @��[����|�7���/�W���aTrvV���a���$�����H�Ǳ��1���'%��!    Pp   FIM�G%��� �,��/=?/Y�D�#�����ȹw���$�E%�����L���L���U�\���0�n��n���U(T,���)��
�P�nW�VK�fS�~�t$L���|�t�6�LG ����1/\��%��!    Pp   F˯J�/$}�� �Lp?_,�PjvV����(�S�Z�Z�nl��+�TrzZ�rY�rY�%���}��i���X���$���h4�h4dY�r����Qj�Mj����o�a:�+�a���8�+�K�.I��     (�   ��$���Y�A0�Ǒ�yJ2��L��%
�����Soo�������4��������̌�l���&A0��~Tv/�*�������
�P�NG�v[�FC��(Cm��n:�+`%�J�̘�1�Z����,?-�ߛ   �w   `��H���~�tL�v����i�1FRjiI��M� FB����uy��#���畘�VzffP����ߧ��(��MM)��t�쾳��l6�b��R��D�C� �8A����l��nSjǍ;��?Pgu�t W ����l���$2���H��!    �ƪ   0�~IҷJ�K��`�Qp?[}�׷m�m[ν{�|^"�ޓ����RGS���?ڎJ#�NG{{{��r*
*
J�R�����}xrP��V�#!��z]���M� pE8fq>~��
���]gL    #��;   0����W$�L�Sa���X\�a~k��᧦���^'J%%gf���R�\�oX��m[�mkwwW�TjXv��rL�9�^O�v[�m���(Cӑua��_�E�m�t W$��h:��j�ۦ#`r���?0   ��(�   �k[�'$��� o,��/�b1`�E��V*����SS�&�'��rY�bQ�RI�x���G�뺪V��V��,K�\N�bQ�BA��L� ��v�n��j��y��H�){��_��/���
�8)�\��Y��q�!    ���&   `�}ZҷH�z�A0���~�����DBA�o:
��\W�����&
�A�XT�\L�/����RrjJ�bq0)~jJ�T��O� �n��n��ŔN�U(T,��dL��'�����7۶����H��0�Z�7��M����jU{����x �X����8օ+H�I�A    ���;   0��[�˒�L�xb��|1�Rjq񱓣��~���'�Yɤ������J�ˊ�r�ۉ|^��'�e�b�kN?��0��8rG�JE�TJ�|~x�,�tD 8�єv۶e۶�1	z����NG^��~���m˫���j���ZM�fSa����dn�6adq�W�$�k�!    ���;   0�6$����1�m�-s�6w ��SP�˫��\+�<5�=Q*��OM)Q((^,*q�b1�\���u]�j��t���{.�� ƹ��N�3,�3�O-�Z�[����z]���뇷�VKn�.�ٔ��N`%r9%��uq�u�)�I���    ��;   0����Lҟ7�c�E�G�ܺe:�1x��jU^�z���� _,*^(���;yl�'����~pp�x<�\.7,��R)�D@����m�V��7	#�h��QI��j&��w��fS^�%1e�SJs�⑘���h�c�m:   �G��   ���Z�˒߄Ka������u9Y��^�s�dR�|^��i%�e�s9������\���|^�\N�ryl�����V�5�=�L&�e�|>�x<n8!�I��	�=�eG�o���u����m+8���uy���Ng���s�q���8օ������    ��;   0>6$}\�ϛ����Gc��(	<OA�~�2��L��'
���BA�|~X������'���t��T��U?��S�����p�{2�4��8�@�nW�m�����*Cӱp�~PBo����v[^�9��~j�z�%�{�S� �,&�?Ǻ��V$}�t    C�   /����J��A0>�j�h�[��XL��`���V�W�]�s�������D>\�?|<Y.�ͼ���u]5�A�DbXv�f�J��7��h�}_�nw8��qӑpI���n���~4U��t��>5Y���5<��E���(��	���C�m:   ����   ������fM�x���hV&�����j�t �Q�Ò�X�p
�� _(
�'�]��Aq>����>]�~_�fS�fS�q��h�{&�y��`<��}u:�a��B�hgX>?����O�ԏ������N�tt I�6�h���)I��t    G�   ?;����_3��qy��d2i:���ܹC� ."�o6�?,�_J,�D.'�����﹜'�;�(��\N����*�g���%��Ȳ�������Q�ە�8�t:�<�t��z��ݮ�nWA��~�#����;������`�z�;��h�z��0L� 01b����#�	�$}�t    �C�   O�.�?���M�xh�ۚ��6cd�oݒ��e�1 `���`b�e�Ɵ`%�2�uT�?Q�?*�ݟ)�T��V~vV��i��eşr�<������E��R{@q��ǑT8?����*���Π�~Tj� )��,�'C�O���J���5   �1�;c   `|}��HZ2�������7 ����W��%Y���r��r��ޓ�����lV�lV�Bax;��*^,*����f�����YY�����$�	A �q��;������X�+�r�U��
轞Bו�8��]Wa�7(��z���=x��s�'&�+M�T �+���#ٶ�	p���A�M�    py��    �*�{%��b��`ıu�x �H�I�۪�n�KJiP|?y�+���EY��p�|�PP���BA�\N�a9>Y*�J���dK&���Ǖ(������9Yf?����p��ف��ͻ������t�z
<O�m�.�;��^�tY�u�����Τt �dn�2a��Z-�0>�$��L�    �d(�   ��%��������ߣe��5 `�/�{x9r4�=���y�S�yO<Y�q���V*%+�>��RJ�J���LF�����K�e����s���N+Q*]K~DK��New]W�^O�^奔n�y����*����=oP&?��^����bzx�sN~�ѵ��*d2, ��̝;�#�4�8��I�&i·   &w   `�}����DC�b���Ţ����k*& ��p����,�'58�j�D�ÂŔ(%I�BA��N�����$��%)���JN���5���<*�[�p��L*��n�%&�'������.�;�~o\��u8��v���;8�#�}��=|^��ɒ~��0��:ͦz��^�/Ƕ�t:
�pX|�@���P����NG
�S���W�8�� �f��#q��)I��   ��Qp   �_]ҷK��n�c�1����ܽ+��WM�  ���J��q��d�=�1}Q��)��5��*���aq�AGS���fK�=�X����ʑ8�#p��B�9N������G?�p��e�N�8�:a"�`�wx韸/�U  �E1���8ƅ�I?i:   ��C�   ��F�?����`41���2w�E� pI������cY|Q��E\:]^?Yh  7#9==��g���ǨK��Ĺ�   �أ�   L��J�s���t��/{��� �	�?�<8���q���?q�NG%��$���  0+s���#�!x��!i�t    O�5   `rx�>"��҆�`�Pp�w �$����U~?�X�b7��+������\4  pi
��1.<�oJ�g�C    ��  ���'��;I?a:Fӭ/s���I!; �xT�]:.��u<�=��ǘl��׏.G���S�y% ��b���q��ؒ���C    �:�y    ���I�zI�t��/��*5=-�Z5 �3�����w�k���_�?���m��� �l�;wLGyLp�I�)�n:   ��C�   �<���HzYҔ�,,�]L��]
� ���x���U~?Y���ٻ���������Ԫ�[j��v����$�sI�s2	K��b���f��X*�!Da�:��0a��@0vLX0v �f�m����j9���T�%��ڪ�[���zի��VOKXu���ƛ[��ք��o�sk,�7�ڙ�  $&�oC��wH��u    �E�   �M�K�F�_ZAgXZZR�\V4ʟ��2p��Z���  �\�h]��>�)��W��=�M�o|4,k���:�^gJ�jx�U��^�݋�:  ع��b{�U�
�X�{�n�   ��h6    ����.��t� ��lV����1:� `c�&ϭ���^	�\��p����  @'�3��y�)��QA�s$-[   �|�  ��v��GJ�Y�� �L���&�]d ��A�  ��ąZG�x�|^a��Wѧ�X�w�C    h�N�,   ��[��<I%� �Ǆ��\t��2     h/&�o.��XG@����Y�    Z���   @�����X��=
�s������1     @�I<h��QpǊ㒞-.   �4
�   @x��Sm��8	�5ɋ.��      ��7��H
%�T�Q�     Z��;   ����J:iv8	�5�    @;�����[��xo��[%}�:   �֣�   �%�\\��oqpk(�    �vJ\x��u�������]I��!    �w   ���.�6��A�}k(�    �6J:d�+Pp�kK��-i�:   ����   ��k$�c��I��I\x��h�:     �Ƀ�#t�7��)I�Z�    �>�  ��S��,I9� h/Nn��D?�|�     �O0�}k�з>%��    ڋ�;   П�Yթ7�#�ܺ��/��      �ܷ��}鈤�Y�    �~�  ��u���Y�@�Pp�:&�    �vpA�ā�1���S��I���    h��u     �^(�;�~�8� �ϫ\.+�O�͜�ԧj�c�#Zz��Q��U8rDa�h     t�H2����8tHɃ5p�%r��u�������FIwZ�    `�V   ��U����I�LZ��rڻw�u���S���ОG<bպ��\���������W�P0J     :MtpP��ϯ��/�H�C�4p�E���/�u��㽧��_�4m   �
�    �"�M�^k���d(��RllL��1�<�a��S|    ��D��?p�"{|�~�"{���y�ah�qJա,�:    ;�   H�i8�%�q�1�jL�j����œ'����Zz�������C*�rFI    �v���S��A:�ġC�B��C�[G��L�:�#�t���Z   `��;    �:繒�#i�q�'�/�����k��_���˩x��
G�h��-�<.<���D2     ڮ6�=>>���.R����m    IDAT!%�Ǖ��Bɤu���І���>a   �=
�    j��rI�gA�p2�sD��4p���R�5,�岖��Nz?zTţGU8vL�G����`�    �n�@��1%�?�~�8��(y�r��uDl��}��n�   �3Pp   ��vI�I��:Z�����E�J:��Cڻf�/�T���N{�|P�ǎ�xℊ'O�3�    ��\$��y�)>>^-���WK���J<� ����`hC�[��lIe�     :w    k]'�1�~�:�������b���+>>���=lպ��{� ��w    @�	�Q���;�Ğ<tH�/��8a��3���%�L���    ��   ��,�i��� �.���u��{����ܺ���'%��    ��bgJ�T����b���9gmD����*���!    t
�    ��CI/��!I���!����F�9�}��	���ѣ*;��[��)��    ����٣���W���_��Ptd�::�i���%�z�    :w    ������k���y�v��\,����J<x�:_��t�t}�{y~^���j���	-?n�    �-�XL��1��ǫ����j�}|\�.P00`]�ϴz�iI�K*Z   �y(�   8�WIz��߰��`���E"N~����K���|�v№|P��e��    �v�)~�@��~�@���r���/9g=�ϴzN(�Œ~b   @g��   �\BIWJ����Y�L�B3�Xl�����{��qO�<3���	���%�m�    �,�w��㊍�W'��LaO��+z�yrA`}��{ϙ��q�    :w    �yPҳ%}ZR�8viiiI�JE�H�:
z�s���)66&��/��ڗ�*��Uo�����'N�)��<)��Ap    �/k'��FGSb|\�/T�LZG(����Iz�u    ���;   ���Sқ$��:v�{�\.�={�XGA�s�h}��z|�������Z>q�|��Iy
�    �����J�=>:����
	��9�>�BO8&����A    t��$/�Y`�9�3  ��0-��I�]�إL&C��E"�	��^z�z
�    P�^��6�=1>.�[Gv�vEBt����Kz�:  �l�9�=u6�����D�I ����y  �^ҳ%}K��mSt.�^�i>U��S��)O�T��)�N��>?uJ�S�Tf�   �V|�>���W���طO���S���߿_��1�1���ϲz��%}�:  �|�{���uΕ��1�$ L��  ��1/�Y������'�\(v�y��w��~���ƗJ*��k��q��檏W�����U:uJ�B���   � �~qwtT��������⣣�_p�"�1s9���>#�u�!  @נ������  �  �v����$��:v&��ZG :���W|||�m*���Ǐ�8?�����Ǐ��R�/�8��'�0lcj    �":4T/���Ɣ_�<���ׁM-,,XG������z�P  ������ �{   l߻$=Aҕ�A�}��.24��K/�F3}���ܜ��N�tꔊ�N�x��J�OW��̗ͩJ   ��ۻW��1���Sl�߷O�����\$b�	\���-Iz����A  @W���9�})*i�: sE�   �+]%�%���A�=����b�8���n�K%��Y���|�D}|�$��ɓ�L�   ̹HDё�������QEW����W�HXG���ڤ�oY�   ]�N+��sŨ$ƈ��  v"/�
I_�4b�۰��h�+.��c��4p�nW��T<~\��y���U^�_>v�Z�?uJ�B���  �����|tT���jY}lL��e�����s�Q4`XC�z��[�C  ��D�@&*��;}�{��  �Sߓ�2I����.A��L��!\z�α�/������U^� �T������   :A��_��k(��
�ׁ��gY]�I��  �k�e�@���s�   ��W�/�j� �N
���b���+>>��6�X��S�)�O�������*/.��r_:}�i�   �
��aE��O^��<n\߷O.��
�E���uNI�\Ҳu  е�}�9G��$~  �ݻF�#%=�:6G��m.W������sn�K%��Y���U����W�'�ðM�  �/�CC����QE��_)�Gk����S�LZG`la�S�]�"���~b  t/�����[@_��/D%�[`�	�  �	J��.�ے�g�&�٬���!���X�:�rlL��Η�*g2�"|�˩4?��J	�V�/�<I   g�����퓋D���Lp�*���)�  ��A0ｷ���B�{�R���Z   =�I/��7���Ypa*��jdd�:
�.�ѭ��P充3S�W
��充�D�LFa�Զ�   ؽH"Q���g�b{�*:6��޽��ۧ�=g���8���(�w�;$��:  �~��c� �;��!������  ���)I��������)�h*[*�K�/�T�fם
_Yy\���>^X���
  ���}FG:�xp���A� ���ҒJ|I��'�ْ�  ���!�6}�h��� �oι�3  ���&I���	t���E:t�:�>�je�m��+�|u�ܜʵ��\}yinN��E�0l�{   �Dѡ!EGG����QE���<�����\|@�[XX����-J�\�� @S�e �A&����	�  ��^$�$=�86���t��2|r_̩M���r�"|y~^�l���\N�S�T)��   v.���NR_)�G��_��)>:Z/���V z�au�P�K$��u  �;�0|(� y��Rl�D�Zg   =�(�钾!�|�,Xӯ ��Zl+*��J*/.��ɨ�ɨ�r_�d�������E
�  `עCC����o������E��>_YU�LZG S����pno���  �������u ��sG��\r���QR�:��s�寻��zի��  ���SUK�wJJg��l�: ��*28(]x��Y;!>l�_��S%�����r*-,H\= ���8]=:4T��VdpPѡ�U֣{��E"ֱ��Pp�h��4m  ��뮻����lN�֦� �5�l6{$z�WV�������u" ����s�3�  �U�*�zIa�1� vf;�%ɗJ�I���p�_��S%�[��<7�r>��w   ֳ��RllL���Ue�h�r�Y�����d�#`}�I�B� @�9�|:����_���ĿNOO������s��;Ї�s?��   zޭ�-�*� 8��� �.����ƶ�O���J6����٬ʙ̙����a>_-�g�
�y�\� �u�������aE������ޏ�PV����� �rI|�  Z�����HRT��s?���J��� �v�Zҿ��k�AP��A �\A"� �P���F���+S����Y�++��Tjѻ `g6-����^[��/� :�au�Pҋ%��u  ���}��io��n��	��  ڤ$�i��t�8��A �E;�_C9 �
�� ��gX���>j  �X `�6��Vp�w�?�a�]�  �oU�ҵ_�4`���qr Ш���|�z_(����J>��PPX(���T]�˩R((\Z�$ (:8�``@���"��)20�������Y���\,f�  = ��XG��K��  ���� �����Rp�t�a v|,��:  �+ߐt���I�[��r��*��"��u @��M9��W*��{>_-��J����*���2|��r>��Ғ�ʶ�|^�� ���j�|`@.�P$����P�L�.���Ճd��6+� �	�#�껒�o  �H$rO�R��2�w���=R�:�>&�Y" m眻rr�g�s  ���vI�X��w7�|����k ��
��d�����Ҽ_^�����׶����+����"ey ������x�\$�
�zY=H&I$��j)=����I&:�>�~G  4��^/zы��u�~wRң$��:  �/�t�~I[� �>��SSS�3�%�^I�m	��=Wo   V^%�%=�:H?[\\�� �9A2� �lʱ|���X�����j9�P�J�z��R,V'�
���R��_�X]���P��T��@�H�^(b�j�<���bՂy2)�U�I+� ���W{��W9�� ��r��v{EI��v  `�Qp��s�;�Ǎ�{D��+ι{�3  ��Jz��oJ�y�,}kqq�:  ��b��b������%)U�����j1�\VX,*\^�.[ZR�
W�=��Ru��6a�$_((�T��?�o�,��,I*�r-y����䜂DB.��F$�s��E"�y4Z/��h��.��}�x����F��@��� @��+s^իp~�:  �Oι{���Y� �V�Nk�����s�& a~�:  �k�&�+�F���%N `�V�mU�~=�����\�/��Pa>/I���aX�4�+U
��~��佼���l/��~e�f�0�>,���3�K%I���W
�>���b1�$�)�K�Ҹ�j9���ʿ�ιU�>G�����A��A+�DV&���\<.9��ʱ�����Ū�^  �>�2w���b  �/��7�3 h�z��^p�F�_�pY\���a��  @߻W�%}DR`���p� ��S+G�sl��T�����p�eE���:ˤ�R����S*�R,n{�F.Qd�%�`�~��DB���.�P��^�֋��}k�r  ���d�#���$]o  ��H$�5:�@����x���t:���ڞ����R���  ��M�n��o���+���      ���������Y��G?��(I���   �����{�u mq<�J�_{�jB�s�i�@���u   ���t�u�~�,      t*>�21/�2Qn  �{O��_m|����8�@o���  �I��+%}�:H?Y\\��       ���{ە$=O�?[  ���
��U�ֵ�/�7 +��/Zg   X#/�ɒ��/(�     �S-,,XG�'^�u�*�  ��A@��ι/6>_Up��rߐD��}����=�!   ��SIOW����     �N�gWmuXҭ�!   ��d2ߑt�:����ݸ`U�}zz�,鮶F`������:  ��.�E����2�      �T|v�6wH��  ������s h�/^}�ե���-��_h_ �s�� �N�aIo������J���      m����[�3%y�    �@��}g���Up�D"�2 z\�R��:  ����X��u�l�:      ���^�\�:F�{@ғ%��   �K�tZ��Y�ֳ
��J��v`�7�p���C   lы%}�:D/[XX��       ���d��u�^� �2IY  ��J��>� Z�9w���_�Ok��Up_qG�� 0���u  �m(Jz���X�U�L�:      ����u�^V��<I�X  ؆OX �2��knTp�У�s�| �ns\�S$qV�8Y     �N�gV-�%�J�'��   lGtހU�T���^����f�N�G�^t:��~�:  ��#�
U'���8Y     �N�gV-�vI�X�   خ�.���%������d�K�X��>==]����F`����u  ����?Pu��daa�:      �
���[I�[�   ؉+���"�S�9 4ݧ������V�[p�$��_�. ι�a�  `��-�u�^B�      ��Ϭ��^I�I  ]�{O��=vZ7,�g2�;$�W#�;Ng2��[�   h�)Im�W0      ���{S������A   vcϞ=��t�:��Y�`�+3lXp���.x�?ޚL ��{�����u  �&�#�k�Az����u      `
�M���TIZ  ح����$���������VnXp��H$���`��g  �c��.�t�u�n��B      t�:�eU��m  �Y��t���qΟ�s�?/�XS� ������/[�   h�9IO��ەL&#�u      ���6�J��   ͔����S� v�X6��¹68g�}zz�,�}M�����uzz:��  �ߗt��/[�s�P�L�:      P��U�v���u  �f[����:��q��������Yp_9�{$1��^�s��S  ���%�L_�ۡ���      �$)�˩T*Y��fwH��:  @�8��-�b���y���f�lZp����Oҗ���ϥR��X�   h�H��ѭ(�     �S,..ZG�f�(�b  �a���?u�}�:����)�J��f�mZp��S�t!~~ @9,�ϬCt#
�      �|V�c�I�}I�    ��!�8�Km�ӺՂ��%��U" �d2�  �F���:D��!      :�U��IO�t�:  @;�r��Iz�:�m;�G���
�K�޹�H ��9w���t�:  @��D�g�CtN     �S,..ZG�6�Nn��u  �vY����u �㽿u����-�%)���$��@�X��6�   ʒ�!�[�A��ѣG577�r�l      }*C�������M
�~z�u   ��,��P�D"����n;G���y�s�y���ݜs�MNN��:  ���%}U��Y�&�x\������p���e���S$��     �W*�4??���y���i~~^�\�e
��:n7)Kz���X  ��N�o��R� ����T�[�8��#G"���aH��|�9��   ƎIz��%���t�b���Ǐ����n�Q~hhHCCC���ݻW�m�;�      �@�RI�\nUI=��Ջ��|^�lV���:u�*��u�^�%M�r;  �sA�=×h�Þ�_o������N�ӟS�$�s}"�J=�:  @��UIwJ�c���b1kppP���;�_+ɏ��)����     ���zc9}mq=��)��knn�:.�7H�c�   � �NBғ�s 8�ϥR��������aRp:�s���   :�ݒ�%�c���Y�V�T��ܜ���t�ȑM�_;~m1���      �MYo����y����0�����KQn  ����aRp:���Î ���wy�s'�h-��g'''�:  @z���K
����b��FFF422��{�jxxX������p}Y���Ȉ"��ul     �-	�P�lV�L�~[���l~~^�LF�R�:6Z�IO��7   ����J��9 �뫩T�7��ӎ�����O�d_ ����	  ��}P�!Io���*�J:}��N�>��}�񸆆�488X�_�_�5N�߳g����F     ���h�z�V[����癰����LQn  8KoÐ�;Ё�0�ӝ��k����J�����%�.�J=�:  @��Y�X�@����ke�Z9��߸|�޽rn�v    �.P+��������/..�R�X�F��O�c$��  Щ�����o��*_K�R��Ɏ;��.Ia��];�@�y���:  @�F�IWXAw)�*����ӏ��-�S+�ixx���񃃃��S�    ��ڲz6�������z��9�J%���}G$=Q��  6s��W��d�!�s;���9�N������1 4�GS��3�C   t����Jz�u�Q<��𰆇��g����hdd����|dd�>9>�LZ�    ��,//+��)��*��iqqQ�LF�LF�l�~[XX�/+�ֱ���U���    �`vv�����Y�  y��vjj겝��	���a���`7��kIl  ��%=Iҗ%���Y��b��ӧO������/�kttT����&�7ޘ    �F�MU����eLVG+Hz�(�  lY�\��H$�d�`�� ^����L������s���q �s�=���/��  Ѕ.��}G�1  �IDAT5I?k�0A1    �.Ձm)Kz���X  �6�����޿�:�ϼ��}jj���9Ʈ����F"��I�� �H&��  ��QI���$���Y��+�:~���?��}�Ѩ���544�꾱�QQ>����     Z�\.�K�k��ճ�l���:�e^�u��  �#�H����3%����%�ܮ��KM��.I�t�5�^ߌcضT*���  ��%���C�������V��Q�   �&��4�����yy����O%M[�   �f���)���u�9�^399���g��%)����H��f��}?��l  �|S���4h��Y�bQ�bQsss��w+��������    ��YA�\e�b�h���$��   �6<<��L&�I��u���(��4e`sS&�KR:��\���:�-��T*�)�   =�ɪ^��6,�c6+��b�U�4�Q$�~    z�z�R��j�FS�k��9�Iz�u  �^133�D���s ��{����Ǜq���%)�NR�e�<&��y��zjj��9   z�s%�OmV uk�XL�D⬩���c���\S?�   `h�	�[�XT�\^UP_XXP��o@g�KI/�  �kfff>�{�u�OܑJ��Ԭ�E�u I*�˯�F��$i���p��H$r�u  ��I{%ݬ&)@�*�*��������hT�������@��xK&�J&�g=P2�l�   �O�P�ߖ���������jϗ���%��햖�����n�t�u  �^��s�	�Ƭ� =.罿��lzYcff�Z��ۚ}\ gx�_>55u�u  ��jIo� �'���q�b����׶i�&�F��GFF�p�
   t����R��b�x���b�x�T������|>�L&�r�l�V ��g%=Iߜ  h�t:�rI����kS��;�y��ܧ������������c���_J�R�w�y�,   }�m��� �V+����z9�V����������
�   ��4�΋Ţ���b��rz���Xd_XXP��o ��+��(�`  ��y������$��u�G��%�\�W^ye��mz�]�>��0h��~��Kz����}�Y   �Ȼ%��: t�x<�d2�d2���!%���Z)>�Lj``@�dR�DB�DBCCC���J$�u�d��<  ��R����e---iiiI���*���rZ^^���
�B}������
���Ţ�����.--�X,Z�% �Tߖ�XI�    �`vv�%}�{?h��1�A�����w�}���%ivvv�{?۪���9�����[�s   ��@�G$=�: �x<^�_�$�ŔH$���k��'��b1+���  �Wզ�7N;/���k�����޸_�9 ���Q��>o  �����WH��:�c&R�ԟ���-+�OOO��ß��V��O�s�����]眷�  Ї��>&�2�  ��i,��&ȯ7E~``@�H�>y>�ippP�hT�DB�dR�ht�z  ��h,���e
-//�\.+����/--�\.o8=�X,�P(�*� ��}�~K�1�    ��{�fgg?!��M��r&�y���tؒ��5�>��=����u�>p2�<����:  @�K����[ t�Zѽv�v�|�4�Ƣ��}�N���bP�o ��q�I�R�����q*�z�k�d2��e� ��K�͕{   ���9���W��,@�[(���馛Z��MK�433���Z�:@�{F*���u   (!鳪NY ���ɤ"�ȪR�����Ѩ��䪩���d�^�w�ippPAԏU+�מ'�I�	 ��
��*��
���0���Ҫ��|^�{---�T*�P(������B}2zc1�v,  �ਪ�)~�:  @�K��O����9�n�����[�-/�KR:��M�K��Z@zG*���:   �%�)���A  h����7>n�H��6����ݯV� t����k�����Y���N9�h������=^ZZR����  ��iIO���    ����}�����9�n䜻mrr��~�h�_@����5��ÿ*��x=��|#�OY�   �*YI�#�K�~�8  MQ+�r����f��J��488(�ܪ)���%ihhH��D�H$$�>�c �D�·$��yI�O$����eU*I�����ƥ3�Ͻ����Z2_{  v,#�2Qn  �(����L�W%��u��ܛ�d^Վj�wI:|��	��nI{���@����?rjj���A   ���$}Yҿ�  v�6U�9�n~``�R}�|߸>HZ]�_��_�p/UK�ιUy� �?����N��]S�T�pI�ޯ*�׶]�,�X&�M��kiiIҙ/�ݿq}c��{�J�R/� ��������  �����o�$�~K�� 6����T*�/�x���%iff�J���h��]�{�655�q�    8������:  �/�E���������U%�D"�H$R�v�}$���kje�����x�F�S�%����Z����&�o$�������^�X�>�B��0Ϲ�\.o����V��]�����Xk��a֋ݍ�X��1����k���s�(j�r  �6[��4I��  �����<�9w������gMMM��v�`�(����$������snzrr�O�s   `K~N�)L���   �}�2Um�   }�(�Y�n�  �����L;���:�ɜso���|u;_3�|���f�$��~]�[8�n���x�u   lُ$�����   �}�Ţr��9o��  �NI�D�  �k�R�?��W�9�N����_���~ݶܧ���J��\I������w�0|�s�o�)   :ȏ$=N��     �~U��BQ�  �*�9�U��oZg:пT*�g]y啕v��k�ּ��o�� �.i�U������R��X  �����/I:d      @�����  ��I��?#�$�o��'�0��n��/��	�5+o��%�2 ��9�w�]N�  ���P�c%�      �-(�  ���e���Y���{�U�]2,�KR*���s�Y�ʖ9 c%��3&''�n   M�CI�%w      ��Qn  �!�T�n��S%�� �*��799�U��wI��������9 #�{���ħ��   ��~�j��A�       Z�$�E��  �S�����bI�:`�{��T*�Q��wI�����{�z����LMM��:   Z��+J�      @����?h�   -�J�> �5�9�v�޿~jj�f���4J��o�t�u�������&�s   ��~A�%4�      `�(�  �t:�FI������R�ԫ�C�tT��{�fggo��
�,@+9��>99y�u   ���$�)�u       ;V�t��X  @{0���9������9�u���:@#真��|�s�6�,@�׉�����   �⻒� �u       ;R�v  ��399y���V�@�/�ɼ����R�ܥj���/��$��:���f��-   �M��~�:      �m)Kz�(�  ����r���N�,@���K.y���thd-g`#�{7;;�g����4�-����Pn  �{�"��ƭ�       ��v   �{���t�97a�h���r��+:��.up�]���g$MZgv�9����ɛ�s   �cPr      :�v   �233s�s���9�]���́u�sq��T*���:�,�y���)�  `�{%=Q�	�        �U�t�(�  �����[����Ա�``�K�R���r������ξ�{�.IQ�,�U$�"�J��    �XWu��~�        �j���n   �ivv���wK�Yg��✻frr�V� [�5wI���}��y��� ��y�������A   ��(�      �#�t��w[  @g���y�s�%��l� ���T�#�A���
�t���W�T>���l�����SSS_�  ���I�%w      �RIҋ��v   l��Ç��'%�o���iIOM�Rod;� �511���_��]�,�:���?�r;   ��ے#��       @�*Jz�(�  `&&&�Y�T%�n�,�:�T*��r�ԅ�kn��ᥥ��K��:���x���^{�u   t����I?c      �#Iϒ�q�    �N333C���{�u`ŧ���o��� ;ѵwI�޻t:�'ιת����wν5�ɼzzz:�  ��w��%�_�      􁼤+%�a   �m��z�s�?K
��9�ޞ�d���NkO��ggg��޿[��,�;�J�R�  ���_Ւ�í�       =,#驒��:   zG:��\�{%�ZgA�Ytνtrr���Av�'
��ַ��� �����:��s�[�J��n���Y   Г�I���GZ      zТ�'K��:   zϛ���K���_I�5�,�ߓtE*���u�f�K �p���f���{�u��;��=�v   ��iI����       @�9%�E�   -r�M7���G�m��l6��^)�K=4������s�s���;��N;���^�|   �FR��H��A      �pR���m�    ����Wx�ߩ�U��f����������4[O�%ivv�b���$=�:z��+��U7�x��A   �w�n��{�A      �.���'J����   ���������r�=�.�΂���H$��믿�G�AZ�g��w���/s����~�:�V�{?���f���C�0   �[QI�t�u      ��H�$��:   �S��*鰤!�<�Z���?��NkO�k>��0o����Y�]�s_.��/����?   :���IWY      ��wU��~�:   𖷼嗢��m��ߴ΂�� ^611�]� ��wi�7_ҒF�w{�#WY�a�y�lw4ݖh��J
H �!�"	�E�`P	��L��"d0 m�j�����e�ƽHJA�!����B�@����s^?̖�B-��3;�/��O�yv3�d��yO�ս7��v�����I�$5� �\�:D�$I�$Ij k�3�7R�H�$I��Coo��1�>��{T�Bo�y��3ft���WS������t���
��OC_Mݢ�B�]�R��9u�$I��7 פ��$I�$I���j�`g�I�$�}���N�1�c�z�է���j��ŋoJ�2��n�[WW��B����-�υ���啩C$I���t=p-M��N�$I�$I� ����C$I��������cS��n�B�~�\�e�
�RY�j�?�̙sKkk����@1u���c��X,����X�:F�$I�VS;}��K�$I�$I��� J"I�$�U�Vm8���>88�:07�M+��V��;w�hɒ%Oݓ�������M�7�,u��M��Z�^�hѢ�S�H�$I�ap3M�%fI�$I�$i�/�� 1q�$I��O�-[��B�p#p1������BW���SǤ���]����*���S4�	!,,��Ϥ�$I�F�%�π���$I�$IR
X,N"I�$�����c������N��wb{$�pU�\~:uH���>z{{O��|)0+u�Fݟ�<_|�UW=�:D�$Igw�S�H�$I�$I�(ݩC$I��Ѷ|��,[
���E���,��J��R���{���}
��OO���Bx<��e���H�"I�$�����O��$I�$I��� ppG�I�$i,�lZ�n��ٽi]�p�!����9p��)4��7��:;;M�"I�$�������C$I�$I��1�� x8u�$I�4^zzz����v�ow��Ú��/������<� ��{�v��ʲ��\.?�:F�$IJ�j��;&u�$I�$I�4^�6��[�I�$)������y� �pPLݣ4�̲��T*=�:�Q8p����ӆ��.!\��G��B�}xx�'�-z)u�$I�T�����$I�$I�F�������C$I��Ժ���B����G��B��.��/��i4��Coo�G�<� ��"�=S�����b�����J$I�$ՙ"p�Ӭ$I�$I��F�8x%u�$I�TOV�XQܵk��!�K��pӚB�ܚe�ݥR���A���(Y�|�Q�B�1�K�i�{���!�;B��J��R�H�$Iu���8u�$I�$I���B� ���$I��YOOϡy��Ͳ�{1��R�4�7��Y���T*�K38pe�M�6ͦ6�05q�D��}�q�ԩS�7o�P� I�$��� \�:B�$I�$I��.S�H�$I��R�dmmmsB���n�(Bo��1��u�9pC�J�#S�L9;�x�`J��&� ������ϟ�+u�$I�����B�I�$I�$i/�\
�C$I��F�bŊ����Y�o>p�ہCwm߾��J����A��qR�TZ���f�.���{�x(�xo�X|�Q�$I�4�����!�$I�$I�D�F���!�$I�D200Pشi���91�s��S7ձ��6�+ݴ��tuu�B8�p*�}��6�1���;;;��:H�$Ijg@[�I�$I�$�}T��"u�$I�4�uuu}�6�$NJi;�ݴ�MԌ�ׁJ��2y�䓀�B��Y�A���ҫ!���y��zƌO���WSGI�$IM����L���$I�$Ij<o��N"I�$5�����ƍON˲lv���'Sw�����1�'��;w�\S�T�SG5;�u���o����,�N�1|80u�>�
��1�!<U(����x!u�$I��w<��C�$I�$I����M"I�$������j�:;�xb��� �׀gB��<_����dGGǆ�Q�_�H__��CCC�gYvpp��u0)a��B�q}�e��y�>��lKK��lI�%I�$i�<�:D�$I�$IM�e�,`m�I�$I{���?mxx���qY�����!�#���zӺX<�����I�&����x%a�>�@�Riikk�B����4`za�[B |l���:��`ʻ~�v`�mvQ�f��#�7�m1�W��!��b�[����3gnnoo���)I�$ilM� �N"I�$I�����<�:D�$IҾ(lذaz�P�B�c<8(�p0�ݴN�G���M� �-���#�Wc�[��Y�m�1nޱc��J�2�� uG��\�    IEND�B`�PK
     ��d[���  �  /   images/a5640015-ff5c-4848-bb8b-6d4b42e5489b.png�PNG

   IHDR   d   ,   ��U   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  eIDATx�՜{��U�����nw�����n[����Db(����!J�Mj�$`$��	j�/�HH��"�JA+[JHw�ew�m�5�;3~?w~w��tvf��-z���������y�o��з�?��m���G�� 7Z0���,�HX2�������0s�k`�����gL��b1�f����㑑����6444�f�qM&��cL�7��Dr��vy�ZKK����Y}}��������'��sm����� �(q�	�@�N�b��z q>PH#�T�����q__������?�u��	��O��&��-�¿袋�q�TKK�1	fX�Rz`�Fzz,%��RB\+�Vs���ga�#i�C�ʈ��}P�C7�ߊ��=��`	>œ&M�z�~��u��z��s�9b�<�=z���L������Dr�x��R+M@ )	s������^�A����n#���֪�I�R}0�c�l�P��r��S����J�0�N��@��9Ӫg̰�E��a�76� b���p�4���O���������_�y�B\'��MҤ��->y�%Ĭ�Vw�V?�;&��9��2��i� �H��wX�=">t��4�'-Huu9�<�S�[�}�;���c�ſ�'�ZXQ�7�+�0��!i���n3W����N���&����jC�����[l�YgYV��0+��  �=�����G�3�/�o}b����s�lD L�D�|�����\&4�<@��Y.:��EHQ�P|S�A�8ٙ�c���o��2��>�Z���A��Д)6 �����>���H��ng�`K�);?"��-h>��
��O}�x���$-h��얦�459-�;�d�|�IϮ��a����Q�+*�E�-���Y}8rV$&#!�'$��r�PeK�Xϛoھ��[--�K��Z�T�='�O��0m���6�	�n�<;�3�i�
�1]2Yh^\��u�0@�͞]HC P�U�E����C�+
��dav�@���6[~�A����6._n��l�SW�����Fנ
 v�{�HpI	�J�̀��(�i��i�P��ò�������NZ��� Ǥ��ɣ� "�el� ].���e������4��T���g͝kS��q�B�u��G��S�G�Q�'?i�n�����oC��oq>C+��3���f������a]��u<��(-҄�{�؈�cQ0"=�Ƣ�Ծ"��"�� i_:�I7Y	���Y2U���r���@�*;팸V�k8o) � 14�A�(��ߨ�5��A��t qy ��,]Ӧ��BCF�8>���9>`�� �����|"�G �`B�	>DH|c��Z���1��@V�X�����6,�&���p�*g�d֪,L���߽��B�O=ՙ(2����Y�;DB��X�@�"�� �;Iya�e�D�:=Q�V��p�d��ciiW����O?�&�U��d�;}_���f�\�L >�4M�%= �)h(c,Ah�� '����Z�ż�je�Ah��� �B
�Ci�7�~��,sW�� ��*�Qڂ��g�~����8�|�����SOS���.���[�mVA��3����Ѐu)EM�.��������޴�!�iO�򓆏ܚ���<�'���=0�Lr+��g���6N=�D�7��_Jj}�U�*W]~�'l���g��Qѝ�h�RI%:r�t���$p�������euO���]�I��Y�0xH�*����KQji�����x�&]3Yf�Gt 5�i�\E�J�mmc��ʕ+[�j�U���$>W��1����K/ھ}��:�O�3=_��de����R7�U*�]I����-3C����P~��m�Bט�V|���u�F��b�sk)6R-�)��B����1Ν��޽{��r�9s�g/�䒃ZhI{o�:�ϋ�9�%u����t{�0LҚ5k�D��/��PEݣ�QNw!i���  ��LBP��@RҞ��Id�Z�Iq"(s�DP�|�r��瞳9k׎�'�@l�Q��o�V4֯�1��ء����~��2�oY���������2���+1(6|�+����}�'�
�g�����Kve<�Ջ��w�H���,%���.S��1�FM���_�+�H;b�2/cb<z~��EΌƂ�� 1��˗��/���XF P�P08�$�k �yk��U42R�J��g�e�m[N�EV�c����D��G>��d_.g��-�K/v�Tň�1��^{�R0�xo�] Yl" �bb
�Q�!�wA����Bo�A�s�Ǜ��@l89ߔgr�#��^V�/sc�̵��{����TN ��wK����S%4�
6�<az��\�U_�u	$f�>P�U4��b�	Y=Ŵd�sD3ʸ�V�@�ԡ7�d�?��")@I46�ayb�i���DdUDK�[�'�HT6����|��n׮]�lٲ�N��e��%i��֦o����U��͒3��o�!q9�r�(��b;vX���j
 0G�Z������R�(*1W=�����7���q*���EN�LJhU��e�y�66��{�Զ?��+� ({ �I��ͽ�Z��<"SdQ���/�}()A'�*�2ǃ��H� ���M�M��%�r yD|��h��I�s�9�7�|�o�k6m�d\pA��p�:_�c�z��R�B�4]�S�|�8܅�ҹe��\~yY������h��ڂl��~��kL-B3H�������>�쫷n�ZN��fϯ-�f�K� �
�*u+��+�D����k��?�p��ɵ�]g�Ѵk���e01��2x�%�F�DZ�(���=�i���g�7n̕��!%Bj�sؕ�b��������y���u_:��Γ@yiݺu��\s��I%��@F��o�����B�'���l/�7EV�|rɞO����$h��K����Ü�~�V����My8t˅����wu]��v��YR.�za��(�j�?,�Q�a��ʝ�ehE�D6Y�A/����-�A��4r6���ݮ۵t9�U+���c����z�Jd龺�-@��B�\�@J�5�_�
S�t��*��x VnB��z%�&�0�����&sqP~ �nݚ;nc��;gv\7#�p����T���Bh�pM�g�� �*2+D�l��j�p����a�#��+��;��i�v>��l���4c��EPhBF;�ۦ�D^5���ٮ�|��E#,r�-��r����m��	M�d�E@Q򨘢R��*"-V2N��cr�����ޯ�P�7s�jg��?|���`r�#�	�K,`�*��lL�������=�a����i0�����������$b�|>1�l��7bss�[��Z���7��d�Ιc�
�iX`˷���`��Q {-��^�����BX��}o�aIi���뭍����(�8�'�����/���g9γ2�l��Y"D�S��̟o�
����5b{�g��Wd���C_sN^��5��hM����|W!�n	SV����:��6�����G��H��l�+^��ɲ*!ПECB�݌!%_-�ۙ��cG^y����uM�԰X�'�\��#��a�V|�|KMk��+D}g�v�l�fS����~�1p�؊h�,��E(����Y�%hL/��#�z��L{٘���e�}J��D5�]k�2M��6[����C���fk^��E:߭듛7k�l����9GF!3c`,ɠ_��@n$��mQ
,j@v[�}�;��zI �n���Ӝ�p@��A	�[��0�ޜ�f�r�k���HؽA���@ �o�n2>�W��xj��/ �d�@��"��x?�4���s�&K]�� h��x�YǾI�s���3v�h��ӵt�Pv���]f)�c'I�\I�p�_槏r(��O�$�ڰKI�7y��aB�]�?, ��[�T �w�{�%�M�e�L�daR��"�=$a�g�#�� �3�\c�@��X!�ہ�Ycc@�+m�sh�hX��<ely>�l�ާ,J�@���E�)YX,�x��������l^����%ָt�h�@�:׃(	A��nE��������$AnłHilp�����'De����x�>c��O���q�z^^��+�~a)Y�I��\�g���ſDCz�!׽A%տME�W��;��"$ڄX�$w���R՚��1���;��(<�G#�9���1�Կj�{�/r�Q ��x�xi�~*�b�#���klx��Ɯ@�������?����z���|9�8����0ή�R��9��V��� d��-�h�'D��x�����{9t��r�1���x�Ȓ'����Ev���,'_@�g���1�����b>8 ��D    IEND�B`�PK
     ��d[�wp�&
  &
  /   images/1cdb40d8-22d5-4761-8204-85ee5f97d036.png�PNG

   IHDR  �      ��֗   gAMA  ���a   	pHYs  �  ��+   %tEXtdate:create 2023-04-18T17:15:54+00:00SMK�   %tEXtdate:modify 2023-04-18T17:15:54+00:00"�=  	fIDATx���!�Va���1�l�tW�&l&�f�=�Y��`uF NW܁#8�~��2s��<�N}�KߝB$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)�/8�{����a�$_�~^t�a^;'yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yHYN����qr�݋y>���y��r9�WC�ݫa?+����C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C�r���-��.����`�<�!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)�L��<�i���l�6�8�n������f��5IR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR����? bw.g�����9���<pM���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�H~���p���u��$���y:���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E��8�w�q·H~����-$yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)�#=Ng    IEND�B`�PK
     ��d[!��Ů  �  /   images/9ee875d8-7c7b-435c-a3d9-92ac29f03ab9.png�PNG

   IHDR   d   �   ����   gAMA  ���a   	pHYs  �  ��+   %tEXtdate:create 2023-04-18T17:15:54+00:00SMK�   %tEXtdate:modify 2023-04-18T17:15:54+00:00"�=  �IDATx���]N�@@�� !Q���5.ـTg,<;��r��%��z�N:6��0��Ch�1��Ch���ǲ<"�ؕG��U�Ǻ<o�&�3�?"eL��s�?G�G?9�i�1��Ch�1��Ch�1��Ch�1��Ch�1��Ch�1��Ch�1��Ch�1��Ch�1��C�?�-E�w8�%��>.{t��.	ǘ�;�k�2�2������#g�"�*����;�3�KJ��:����o���א.6�*}�v�zju}�.n�&�O�'�aDR���gxA�1��_�ԫr�|�����MK�2���b���:�C/k�u�Z�+���m�����t���.�ʧ��qV�޵�lخ��O;�w�/j�m����ȯ`�!GƮŚ�RC�Y�]Y�|w-��M܎�g{�Y��k5���9rd�}��}���y)����>�4#�/��1��Ch�1��Ch�1��Ch�yQ�K���Oz    IEND�B`�PK
     ��d[	��} } /   images/bbfae99c-8036-4c5e-89fd-a87441410720.png�PNG

   IHDR  �  �   ��ߊ   gAMA  ���a    cHRM  z&  ��  �   ��  u0  �`  :�  p��Q<   bKGD      �C�   	pHYs     ��   tIME�#Պ�  � IDATx���{�m[���Ƙs����8��GսU���袍�i�4��A�("�q�6'9�Dq��E�HEVd��HX�d���&�Н��g=��n�}����ךs��?Ɯs����{����f�J������k�5�x��p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8��}�𵂪 ʳwQʄRZ����k��{�Lǁ�%O�h	*T�J�`011@��#�QD
*B)�@ FI�"4"L�Db4��L[�>T	
4AU0����11��*��J���N�L� ��m��l@�(`\m.@aW��7W�G�|������%���<�Ç?���p8��h��@K�J���s�H��K���EFi��_j��R�kh�,A	P@	`   �jQb���!f(PA�U{�B8��W? � �FE}E��z�T�0b��P�t�>��1�yPr�P)[��7���I�����>P�+��T�hT ��ۻL���J��ui� ��5%Nd?#��z�vH
U�w�[��}��rV)R�""�%' ��f�v�U!�bs�!lJ���x�/.��Σ�~�S�����G����7 xD������%b~�]  A�=��~l�,!	"bz���
�*�E �
$S�
t�Nb�Z�L�WaEM����DՀ�Ĭ
�h�AU���!7�(���?��˯���1(��a��%�۽�����]���$���}i8���U�5�ժ��T�[T�GE�C-�J��eC�����	d�VE�RM��F���dQ�liO~M�?'0�w^d^�b�Op�x<��L�$����3x� T"��q���/@%B���w���w��ڄ����k��3o������k�q����:Eӯӳ� e�n|�Z��	U�M"�7h�Yr��((W���� D��@U�����y��䟽��� �6� ���X��D%"H�T�(�R��0+���	|KLO�x��8L����m.��>��m.@aa�]�%����P��/  �Sm/�J��eM�7h.�SD��J�$_+t�RM��
 ن^X�f��@�aJ��QS�t��k��纽o>c8y�l�BqĻx<������{MH��sF����J�v�������U�v�+��K�������]^\��^��������ԟ��|�^�/�-�p����; t�0�>]=����_.���FD�[%���P�)	R
b�K)PUÀq� ̦���2���_�+t�;������2{��W�~N�D�DF���k��q( �fB8�g���90��2�d�����q��o}a�X	�@�>�G�ᗍ�VU����n�./��'�����/%�n���Z�K*%��Pɦ�T d�ά��H��Du�Z�9��yeӕ�����}N�]�v�W-�~��;?��c|���	s)(���QJA�fB�C`036�`6q��F��,��j�@�.�q�}�_o��v�y�~���g��W~Ƌ��Ǉ��q�`ڿ�_�o~��-������<�Β�o�o��V�|����D2��\!���!F\]_#�(Q�W�Y7ƽ˧3]oqǕ�\`S���"ZM"�� J�jTM1+���y����M`��P���ϙ�gƟ��~�Ke�q�1^\!��1��,���;�������/b�]�����U��HI�Z2 ��"	���`^yۨ�j���l&��mH:��@��l�
^P]���u�{	@��9��s��{<��s�7��.���L@��i��%c��؍6���1b�<b�#��E�0�+l����U�_�������b|�_n���7^^���, "���~����g~�G_�2��W����O�����%�v��7�i��|8n��[���R@*��PJC��`�!9���E��^z�U쮯�(��RU����� p� )�z�5���5ki_2����&�5���5�Ye.1WEO�����9
�'����e~������3������1ݾ��}�������o����!����?��9�.��T��9���I�"')�
�慢�B{�g�Z{�^IU��mt�Y�8��ieٮ����$��qԮ�0Q���.~a�9|*���ÌL���9�((#cF�P��BDĆFly����.�<`Ѐ�p��Kx��|}��[����/�~���T�O@)������W�������~�ǿ��y��/a�yʘ��b�]���o�Ͼ��2r�~��p��3,����4�P) ./v�$ bLsƓ�^z��x�ʫ��
� "���ӅA<�t����<���])U��kH��Wy��P��]��� �r��G��C�U�/J?�!�(��#���,o�M���#���#��p}�����u�П���|�G�|���������e��_�|+��*�Z��BHU��(t�ͧg}	yK���*3
�U](y%@hM߯��@���a�y��`��s����N_�8�@IAA���`F �!�b�
��1�6<"P t�J@���p�勏��W�`xTv���8?I<��ƿ�H���4��.��C   �7��+��4�i�p�x�xx<D
�:�ߖ�߭i��A��8o���� � �3��Md�H���#��9g�./����g�N	�^~��������Č@=Q�z�I��;:_���LV6�^�l��H���_׾6	�<vQ q�P��@���Y���q�� �o�D7x�c����@�P���/�*��A_�����폐����_�^�����Ayz�� � �J�h�V���c��S�w�Vν~I5!�)t�j�/%]š� 뤸��P���x=@B"��%Ct��@Q2��j�H1�Z��JI#2fd8!% `@�� 	!d��������F��:��?����R/�t�{C�o���6=~��v��o�~�qw����AU�RP��Bd�p�:s)�ó�?V4��9�ߍi���p��·m)�I��{H:@JB �%�'H�(iF>�Q�H4(�>�@cA�	�M7�i��;()D �%oz����q�9t�:W�dg�o�;��#����u��I�%�X�a���|����(�߮y�#!���@o}���8~vs���[_�N
��~$�}�y��޲,� �Q*��9�%��kXӀ2A҄��4�z�P���oYY����aJ�E�*��j_�*�cYXk�PN��l-(/4;��.�S*7����S�����	��IZ
� H�H�.� K-��"
5�d0�6؅+\�x�W.���xix	�0"`Ѡa��4���g���e��2���x��p����-!����n��K�u����9��3 �����͗���o�*2��O�\~_��o���O�i��N��y"�3Ho�Z 2!�#JN`"��9!��r�0�nn )!��8D��r��E@q���5~�۰���FFV3#R0Yc���Q�.DW��ޛĉ�~��P3	j��6��*s{ͪ���O�u�y�T�����UM�0(�X
�'a:��C�i�ݏ�{|����Ȓp������/	_W��/}�!l>���(�Z��-��D'@Dg�(D$��I�\��%�-h�Ӿ_|�U�v7Zy��1o��B������״}��;��"�ܴMȋ�iT�b B$�j�,�JBT�[J�A�X���B� �غ �H ��`@)B�6(��3o��4��4 �	�kL�c�O��g���8�0��s�Ͱ�~i������w1lw��t-����@��m�$�9���M<|囯5��۫W?6�~�j���K���U��n�O!�-�dYfhI�r��-E��	I,^.9!oq�y
��0n�u����3�4�c��ͣ�-bܘ�#��a�K�J��J�S���$�U�ng9��޳�R_T�9�h�EƂ�@�����OՒ�J�I9D����)㯕0��D�ߺ�<�����~������������O|�ʬ����O�ւ�Z��!�㿡e�(�)G�r�j2[���T�<s��qن�R�T;�Ψ*t���F��9��z�Z&'銢jT�4*���-���9��ւ�Y�]D@PD
�H%�&����Q�VC��H*�b�#Ka�]"�Lϰ��pF��~ʀ(
�y�&��M��7s���Y���t��1�� ~!����g_�t�3�C ¸�Ї��43�3���/�ٳ=��
WWeh���u0����#��̀�rP@b-}�j%A���BH�L@mX����D���Iָ���Z�X�K���jZ����1�}��p�b��`@IJ�A��AT0� Ί�2f�vD���q����Q��0E�t�c���
����v���}����;�y�%��j`���A����o��I_�"��>z=ݾ��*�E�'E��Z�5D8���h�C��	�@��|DIGS� H.ȹ@0�	ДQ�#�t � C���05���uw��"_? �&[T$K||�7�ӄ@������u�{��KoΏ9\����%/D��=����f_tN��;EJ�֛R7J_#�@uF)�e��{�O�����~����~�w~�w�����V���u��o��|���W�|��K�H���"G�L�2�lJ�%ͫn��1F��Ϊ
��w�yL��M����E)��z�ž6^O�:��׾�aU �Z"@�lB��;��,O�@����z!�$(J��ށ ���l���p0R�Ť���3bQ\L��-�����A� ��RB�v������5���������3S��8��"z�oso!�o�?�O?���q(1��%��f�tv"�w��T�Բk�a � J�s�a�q���	L#�iF�G�M3�:Z2r���<�������}��ʟ���G�q���D��2LE��FG�b�c`��B���L��	, )�M��`bb��Y��I ��H�tr��7�>½�
�����_R�U�Fji����P��
U"����V!�K��R]
E� n�b#��:�Ah�t�����p!P �����^������ 8>y��h
n�S� xh+�Q
�60C�~a�.�J�s�JB��g�o��}�f�g��]4b��� )�����/�9^
�Hy@�!��H�q���7��oW�߂r|]U^*%_�f�P�W�Vb�%��@�y�e>"�(ǣy���-e���'@b��%c:� D�4�e����!�@nn��gL9B9X)Z) ��oN��%�T��G�ÛR&��!��Xe�$��nғ�A+��.R�m�e���Ξ-�K��%�i3 c)lT�D@��H��)�''�o.����nz���O��#���a_+|���f-�a�0o����5_)�R�Ũ'�H-+SA˃T]�oQ�a���g�8M�X�jU�X�6ֹ-���s��2�kѩ
Z)�wR��G�؅["D�Ь(�0A� 6A�(g(B��g��#B�dU*`Q����)^C�
�hA��43��A�!��A�^�^"���{�BxF����D�%����ox� �q����ՌF��� r�0��N����N3�W��z���y `_��"����.
D>����d�"ø9��IidC�qP�AJ� �1�C��n�	1��R؍X�S�4A ��(TsE��*7�\5s���C��L꒮oZP�7�7T�/IAbJ]�i*UΩ�Y�(DETUE��Q��q��THJ	�E��,Y@9�EU���PJ�&*��"���T�\��-�˂�-Ƃq,�~�_�9�B�R����٫Z��*���l��r�^�3=��C�<�������`�hH�޽P�E�#��HyՇy��\i�;���9�ΐ־Y�'ת
J� �(%[-�<��#��M	�fS�R ()4%d�ӌ4O��0#猔R�P#�b�R��0����f�� sg8툩9�M�5[���Kύ& ���K�{}��$ԭ����ԍ�ƪ��ηváv�_=]��p�b� �d�I�oU%��w�VDE�n��2��ܼ�i\����zV��*�ӻ�'{�q�M���/i�sH�G(gh��V�V2���>���@��L�QSƴl�N�t^~��۷}JQ{]/1��Q�&�v���^N� ���M^[�f��FR�`l8��#v�E�2CHl�Q��I�d���I�zp�`��DDe	 &&��Tn��u�b@s���\KE2�L��  03�Ja$#��� V�P�C��8&���(4�(QS&��L���U���(I��+���� ����k����v
�<;��T�i�����a���2���(��r�BsR��H�L��HDL̡*_��i`Bd!��͆i�/]1^}i
�U�K��q�u�V�����û��|Խ�6L+MD$���Ｔ}L_՚����R/n�7o+%Y6qVe) e0���([�DDC9BDTPP�([P�P	[`���P���VG��"�%�HI��R��Ǵ���V�!T�T�c֜7�������Z�̌�{5Z�v<UHUI�����V��b��*K� RX�0����b^}�P�*��g��S�Ħ�i�q	e>�oQ��d�Ϥ-�Rl��������
���cJ8���%��ْ�b b4�:M{H� �S�-iM�@cS���YS���3=]<4e�L��&��7��D]Q�2<f-��w�n.�~��G5�,"�mb%S� ����Cx5���k���n��4r�x��O��Z����~��C\~��雟�m�������'PI֛Xg@��=��F"�j��V��w~" O��~M��S4����z�}�,���歯�f͆��ڇ�d��fc5/{TƆ��BϬPeX�2��Q�D��p���� +#h@�!����!?E. �ƂѕD���huRTC��� �"�z��`G�� ��o�����Z�&�Qz�w��y��CUf�<eL���O�xrTd,�X2B����$b�:
�xf�<�3{�D*}K1�ĀAB���0!h��̀a�������D!�����жt����M޻��o�[}����F�,��'����ͻć��ď*A���Rt�-^V��$��%b�p��[HA<a�`� ���tܢ�K��щ�P��-!l*1AF��lbM����l�=Y���
{?�x�=Y��k�
h1o��Ĭυ4�C(�"E���T{OT�ԩf])tj��u{#I���|����) �֬�~��j��|D"R��<�8���8D���M�l"B$��ʼ� ��7S�(�i>�϶լ^�n�ﲹ�l]���{��*���F��* �:�et�볰<+2O�b芚���ĕ(�Q	Py���P��}������ȳ�O��)<x�[�aǇV��~����@���4���n��*�
��5Ͻy�B���4��*���{����z73׍ghq������K������������E1[���
2�P��  ���
��b,�F:� E�Rz�A+0p(��\`��y
(]Yk5����C#��jV��!�׃V�q���#�g*w�ξ(�/pW�j���1�$I @�3n�7�`�@����D�;WDP�@T0�	%[�b)&l+8�b76RT�	��U�h�\�	~'��}����N�25�6��~��	Z�"�	"]��l�
�{��)T��!@��t��i��#Xf��`�
@cy��4@C��-hs�v�n�p�{_�U=4�¼(��8�2�M�[S�XN?�m�(s�5	x.�5>�3��j�I�z�K���O�,=f�{���'��=@5�\�]q�P�#����JNV]R�0��V�V�3BP�t�����^_B&3��R�t ������ߢ��h��t%��2�O����T��^/�k �Tma��0�����?{�J�KM�CϷ��r�若�E�� ������������'���{�	�|�Sx��oy�g���R��޾�gሇ�UM���K:��G�̖"�f�Ve^�~	��!7�l�n[��%�ӂ�-J����ן�)z�+��O7�J�wLZ{Rj���5�X���ʜ �2�H
��N
S�\@�M�Aњ�7Ȥ"(�}ge5�t�@��r�1�A��`�8T��湒V:��}�*�%j�ΐ�E���m�"H���:��`�ύjڽ���D[̀�� �#O�,RD�l1gV�@��5r.�sF))���!R�e�0�-."a`���UjhדX�3���=(*x>V���-LY��u�� ��=�u4� pT&�NвM7
SX��0���vL3(O�<�'j���J�TD  <��:o �%�`�ov ���^rZ�U��Ր�5-mMZ�ЪL�p��Mq��g�n��[Bz��֥��m�h͏��_H}F�Xy�-��׽�O�}��)��a��$	��L77fP��
�����mă�s��2w�v�n��Q&���	6�U�!��o�N�Jj�u5��]�r���5[��ht�ʘj\���AlD���^�Q�2�~�*��~`�L3�j�Q���`���69W`{��$
�����O�G�+����`��e|X�S�
���ޔ|�'$�T�<hIF�kF��PG��r�V�V�̓v.+ֶ�Im���'V���wS�k�ܳ[�u�z�<��/[�]ey�)��ԪI�l���w&�v�@m��d0g(�*��%����6�%P�Q����4`�r�$3����л���ٵ��^&*�W�*ШUi��P�,lM�����Oj��w��(W�kJc�͆ ���Cf�"(U�81B��� �\��{�V0P�Zl��-×a��|Ļ���u��
H��O��T�C��]�rQ�͋�=����v��(��b�.�`���.��9�ƺrD��L��Ϫ	(
� �	�� %�����T "0,��T�2�)��!� V�._�� ���M�	b��GX6�+��:ٻ��5m�*��Z7�6���S�|��β(������h�Z={ċqQ=z�RKK�2��,Dl}�I��,N���9�!0(0r��b��#f�-V"I���`I��7�f���ۍ�<�?`:$�3dN����z��
�:٫��{�����5��x�M�wơ1w"+�[��`�G�����\�3���}4̌��OU�#֌�z�a	J�������9=���G���'�����q��gq�!m@�S�7��T���%����%�XӒ�e��l-=�]����+���f�����j��$��Ic�٬R:�컀&+D�F�¼��,����*�C5Fd@i�DA����2�b�'�f5+�Փ-( R$�FիoP��(2�5��Q��/#c/��2n�G�A���vo����Rf�;2\@� ���l�r�@�Ӣś����O�\ʲ2wj���k=1�B�l@R0b�u��	9<�f(P�le�2Z�p$F(&���d����Lur�Ֆ�R��
�12�����x0(X'�&�-���.���[����J	P�o�Jm�tU�띪�ꋵQz��-g�R�N_Dd���	:�V#���Wg��
��`L�,IrU�TD���*
���n!�-�b��PF 5�����B���O#�-�e	^�@lFT���<'�6N�5׵Z�ֈ��贌����3�L�Z�ZmHͣ�&�+����o�
o��vT((�e!OG�)a�8B�`�7�W�����O�<��֔��|�s�LG��"6q�V�K����YyY�nJ����^��:��*p���T���85�~�4�3�<�ET_������J *5�*˥�v3���k�$9�/!��O����ç�K/�>T
}z�H��'�|�Ki>|���:!�)	��lJڒF�4�Tzh���Bk1�"[�R��tE�uO��V+�����oS�M6,}�[}d}��x��
��!PH=�k%�����(��`�)�X��>6�	!��MHP��D	3� �z�,G� ݮ����,c�f-�|q�5�u*���m�cB��5���+/H� �������Ѽ��x-$R�9�T���9�Br�� 8��ԗ	`A���
)3�
���2z��@�R���RlT-�R0� S��`?r��y�]>�k���ݵߴ=q�e6�Z���<�~��{j��mˡV���Ȧ�+���6*����D���̥� %�L�3�c�j�V��?GS�f`�	 {!*��C@k¤�A��^I2&��0)jߘ�%le�w2�K�C<�<볳ؿ���[;�K<[����V���.��*!��m+��Y0�*aD
D[WHE)���h��!"�3?~�9M�\I�a`!������./���/DH�1����iF�%3�焠-n^�U(��Da��O7_Ջ���׶6'������ڴ��pL��idJ��.o��oK�]�����M��`�Ř��>��9zB� ��o�7_��v����[��/�>����Q誊��/!�Ã��͟+����<�J2�\l�o+�`�D¢Z�E� 5~��$�d�F�-�k�}+v]�D7VX2�W^�J�T����i{�	�槣�!U2�bk��Z'��`�[v��kw�~�%2� n�>�{�8ҌIf$(PM�#�f0pD�4� &�����܎$t��Q^)iՓ�5������Z�t�i�a=�R�P.��	�2$)����<!���JѶ��1FcD@�hID)�T��"P��{�Rޥ*-�K�=�z������(�^�VN��BJ�F�<�u��'5�AD�O���[�q[y{FEP������PB������ws�fԁ��B$���0K56YH� P��8��1�8�ᵕAB�~i��s^���^'���w��DO�ZU��_�.��B^����!��?tf�����0*~=DJ%�>���Ŝ��[�yBN	77Oq�&�֫���k��/�q��BDPR��`���'����'8�(s��4M� ��j�����@M�yW������BS��o���3�(���Bn����\������nșaѪs �_Z��%�ތ\�1�������O��;�����]|v�o5�&|(����������9������<�ђ[R�1b��%�Y\1KY-~�g�7ũ?���@��y��Q�%�ף�(zvh���3!��n�;�@�����7b�線�F���J�Lv�"@z�0{�v@Ĕe��$�P�g5�V"w(3&9b�	%�`W�}��j�����#@JFN�QJ�`��P��r �լ����h�"�(�F�׷�>k��F��Z%�2 �)f��~5\��@�i&���y�R�#�1 F�u����"�!�keA�sQ�T�Ů?FFL� �ϧ�q'˵�H盡��]��8`�ce���4�e��1&K�9��
϶΀e��ʘ��a�:im�|ʼP�T��R7��{U�x ��h� T�ʆ�5T�/D@f�<IP	�o�������c)��%~�i�n�/K��C��nG�V`(j������k�gM�=�S���I�Z:o�v�TK�<"BQ��������equ��d�>}�y*H�#R�8�v�ǓgO��l0������)%��<�\
�	����Gf��%l���7u�,,�%�ô$�َ'9K�@�r����:�җ�3Q��6�h5Z�:;-����)z�LY�u�2]�r=� ��2�������Q��|y���ǃ�+>,����"����]|�o��S����<}ea6��՚��I
�-~���Xr1�doz~d�z���������j-a�3�W��X��L�L��1*#��e���5_]p��aM�5�A{G&�L`����Q2a�#2f�Z
 B�� ;$��5�02�x��F��x����0F�U����W��r�%	���,KZ�v���߮�sk�c	�F�.��j��S�-	�Z7S��pn}�T�JAI�s.AB�H� �(IPf+�4`�ڎA�%F����m��J�5o�HWR��{�'�����e�`�t��S^�g���JʟP��fL'��d��`��ք�Z��e��["�P5LXZ�F��s�X�n{E������9ke+��u�v�1��Q^+�sZ:A��.9�gJ�mW��E�����]��wj���/	5����p���J�Q����R�tx�iNl//��G^�~������ FJO�1��r��a�ʌ�xDJ	Zex�)�sO}���a]���㥯�k�;"��Ȩ��\^c��V��$����z�S�W����I�z�^#3$��6B���?���/������}��O��cߌ>p��������7�v�돤��?U���J:�%�D!ɐ�{2��R��s��r�~��K&o#�j�2 �z-6Ӕ���9x�ڼ�x�h���z�,����|�r-be(b����q,��2n�P��0}��S��j�6���%aFƬ3�L�2c���l�!�pG�C�ц�l ��xF�R���,�z!��OX])t�$����x�,�{_�V��1w�J�
��� �1a@ҌP
B�Z��X )c.Y3rJ��>�gD�F���E)+R*`hQ�ڞ�4�*������S_���5��[h�y��������0+����e"��Q�EiA��iz�7&2Mlg�$��0��T#+t���Ĭ-�ь 5�Ό.!K�5�l�n.�����ڪ�_)�x�ٛAsj ��v��
���F��I�7���W�S_��("]�o���9\Փ�����QE�d�C q@*�<g�R.8'l6#�FpQ�qy}��|�u���x�����}�� �i�8L38D[����	i^�,����3��s���Qp�F��$c���oxnI���J�\�{j5�:+��8n=1L�����\�e ��L	N��
I>�����0=}��}o���x�o��T���%���ax���(��G�|T&�Z��6�	4Z��K?�Lړ��k��S�Qd�� K���Xka���Xv�2?��Kq��/8��V�t��=ʿ%C�6��"F���������ѫޓ�:oAT�X�M��Fւ$3�L]�[�j��z�bε�e�vW���8>@���:C9#�Yp�����S6���εRWt��}�L��n��lb1�w `�)،f�
��֖��c{(KY�KR��X�%�eA��`�C�hQxUkKlԟ�n�?m��
��;Վr���G-�g�hԽ�h�*���! %,^��>FcQ�GҌ[��5-�7�޲��%���q�8�&�ڡ�@�Pڹm
�Ң���[(Gc+Dj��T���E�:/����K�����װ��Y{R�H���3��(��#pzx{�W���2o�C7ԛ���3*�[�@ss@�qq�4g\]]���#���8N3�d#T_{�%�~�d)x��cd���T0�qs{���{�a
��rFN�ĠYd��lRks��t���8Y�;����K���:�������H#���ۺ�I�Z���~���B[�f	�"��A(vn�:m?rI b��t�^��/��>���;�>��ۿ|`
]U������_���{~����h>��2A$�g#����	�j<]!@� �Z��&&�-�D;�5i:��d�V�D�P������e��k���y�H�b:������;�[Љ
;�Ӈ:�KA1��0b[�Q��)����ژT�@�2*�n�aP����lY�(�R$HP䈩�"˄P�B	�C�Ad��$A�%=����!�xe�j�!<d�Bt���&a�1)���u��{+���E��qq���ŦTJ�BEj��"�pE�����焒	4bX:X��Ա�@$BΊTj�
� I	b`��`?�΄cV0�d=�j��P�h�0�e:��I��v% +ͣ�̖��R
��.���?ۗllPh	�U�	`LK)(Z :!ȡ6	1!�4����$"����JMk_]�F&k-j]�
��l����������4�����	����E�֑ �)YIT��ֹ'���ւ����v�m[v�,�Ѣc"]�-L�:�gevF~�>5�n�Y��+;��i�����w�l/����ݣ+l6�4�����f��^������	�b��<���,'�x8����r�m�{5M���#'
�}y���vΔ�q����L���g'���t9 �o�u]����C뫯'��Z~�U�؜�j�$��I~�������������߂����|�o�-�������=���I���t� 5���,Ѥ��-q2B�Y�u�A��ن�W]j��.�`��O(������W5��w�Z���|�$윾�Y��\� ���7}A���[�U-.W։)�M�b���,����f9X'�b���-CY��?:���@��:C���L��E��������� $�Z�o����,ٺ
�nNUa��ߝ%�����D�c�E���m$"d�q��fQ2�T�p HY�&�D"D��`���5z*�\�X7-����o=S<>�K대dzZ�*ζ:XNH�ԖF��=��c��Z9���a��\�Jw�)Ag��^"E! J1_�,fK����rWB����Lw��(�Evk76Hm?��[	(��a����e�`�|v�������a�Ӄ�&�E�5�Q��f��J. �}�j� h�H�S�f8�Q��q����z�-sga�Z�jkKZR��i\ (6�t6`ETPJF�'����#����a�-B���RJ��v��	2�9c�#a�ݠd`;��n�SB��)8��)M�P%�J�!�,,sKe��{�x>I�<Y�;G�����z���c��3���Fw�c/_���>
����:�	l���a.�24-�D"�%A�d��_���y�}+�>�<.}>0�>=~��똏��W��GJ:��Ɇ���#���T�]J��Z��5�^��K�.ٱ���ߟv�[���`
y�1�f�)�=v}rg_��(],����p
�u� m�.�bD`
��jrגd�(�H�ſ�P���EfZj�U�u���Z�EY��U�	a�#�	*���H�,�ea������DKM�Z���0Е!Ж��0�H(�\=j�GV@R��j�s�&��J�zܘ�$"g˼�LP@����Aр���@V�����L���18��ߺ�qCN�����CS>��;���@Kz����q��ǵ�U ���mF�V�3C�2їw_�Gv^�a}�hM;��Ty���"���d"Y�Bɦ���-=y���=�P��� ��"+O�5�i}�W�\=c�)�O�w�V���*I֝�t�m?\��f1�g��i��[_��&@5A���^�j� ˄i>b�#�`�MeZ.���߁����A�f3"��'X�RPJ�dWǨRs�Ob�f��f��}u�V�ק�)�ޟ��q�峽�����Ým��xr�r"_t]]�Ƽ
 *���=.�2�1���O�g���?|�����	�������UzH4g�o�B��$�w�:9M{)Z������dP9��E���U��Xj?������[��7�*rfMU���ݤ����sZ�Z2%���0%�Ɇ���&�B7Nl���i$��5��דs��SR˜O��:#�D��#����<�;ͳ5��d�&�N�������`j�nBAd�z��^/�s�B*�lXw[k�o����[���L�o�m��a� �%�Υ�Bd����T���U��CR׮������x��w��?���Q�]� �����s��vJe�X������֙��������J�+b�!��i��[+�:e��#v-���K^Rm���/�ql�^�:U�
ъ�4/{CZ��v����7BNAulks�AK|v	�-�	�>9�X��*��_���-�R\
3n��|#����)��A�@ ������vLs�������^sr��@���%��n�#�<M�ӌ� ��<�w��u��{KM}ϟ�����-���'��:z�*���V�ja=TÔ5�Xȥ�L�Kӌ m��@Hy�.�����|��o���>�m��'�s5�Z��+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs����|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�f:���E�s�.�L����)������@��w��{n�<��D�^K6�md�c�pcs��yN���I]�$�����i�!�����9�x��=���b��ko@�[��E�S��y�a1�F�bf���W|��	�64졻V�#���޵_���d���є\[���0�h��9N�	���N�!�2�}���2c��?�ߝ��
���{��HI��z$��W}����7S��o=�|ֶ�����]b4�3R. f$ʠ̠\@egJ��%�Ȼ=�T�4�h��]�8T7�1�j�{ȷ#�i���f^���=�d�w=ܲ
	�1Hg�|_��O�Zb#��cE-cm����>AXj��T M�Z�iF��3ي{o�GE�z�E�8c�v�7�n�6��e��I-����#qs��F{J��w`f,�y+ �׽S��=Ӵ���Í�����WV��H7h�!�kO��6վT�#��N�l�N�E��O�2��e9~-�����!�xS�U�׾�19��?W��NH�w�ȥ�"��x{a�p����Zĺn���|r�j������!,}��}cu��o�2�T�6�;�n���1tKY�&�!{��1��]�}zߺ�F��t�*���ER;�H�t����ǯ����z��d�a��x��iW��Hcx��-`�*c�&�b�ns�z$�o�g�{/E$\#>����ЅQ��HIM����+$'�4AZ2O~� ��yM]#�ߌxn���%���L�ځ��ہ�̣��c @�b^�l��1.��cch��}=��&4��ƒD+oB�#��G=t�b��O�Jid�m������>uʫ��C��i�&�T+n%+n圁��){4���g�$��J��kB����ͥ��V�ƃ;�:�J]]w��{�X�?�:�&���=��������O�m�j���*V�����*C�=,�!���*č{��UD��������ݣ��q�=M�\���58.ɚw�iY{���tG����U�-��~���7�O�o~�e���� �il0�C��Ъ��m-r�� {�sB*;P�~�S���� ����x��:П}�{���9 ���r~+��H�X��ԭ4���}�o�@j�#]�^�*$ [KR+�#��W���s�Ƭqtݱ��m�|�6�]�ݲ$�|zYh[=�=��{zQ���f`�{CX��]cX=
�եz�e��i* 5�¾Ag"$����LDA}L����vA��!�Vo��t�2vۤ�o����j���ĭ>�s�����Jk��\,fqO:5+�Y@�����`�083L��&1���e0+r��guU(ߚ=�/��N(d1���WG�1!� �wX��̽���z�ͷ�kߓ�XQ�d�:x����I�H#W޽Y#)���:M̢���t�܈+�$K�d�f�]��D&I^�h9��� M٢>�w-���ugQ��������[�˼`�ŵ��ͫ��}{{���F?n����%��m�4����>��	�s귕��WHպt K���S����TPe��Ċ�#�ہ�Z3!g��tlW}k�Մ,�c��xh^Dp��Hy�Ϙ�)\ER-Z'	@�>Q�ڣ5↳�BU��?��7�������a����^{3D��m#�2ڂ\�������$"�w��;��9�8A�
��r��\ (�N`ڻQ[@y��Ȼ?��?�7�����?�7Ձ �����_�9,K��n�JOr��ip��0���P��NԚ�x!ء�:*K{���G�������c����_���pc����YĲ	k�Yi�L��M�0i�>�O7�77������ɼ,�l{H�7�Q�L�F&��5ܷ�R��0�> �c}����5�%��� 6���m8�/�Nv�j�$~	��A]<a�:s#\WEU=������hJ��-R��y�x>�Ɋ���p�4N���*�f�kǆ��q�'�:G˩E⑏��5�QJ��E��k;������0<�/tv�ֲ�"�PuHޓ��i�l�����'���f�71�:�^��)!!�Y�F�i��^��̮�X.���R�.��*VX^�6�Zl�^X��t�Ϭ�$C}r�n�I-��g�����]��^�W����X�����ӫ\k`�f
p̌R\��>�4�h�v�UR��5ۏjkX*0�Z{V6�͕dG� �_�{���P�u9�I��E���5r3��#�Q���-b7�"]���=j�Q�d��^6��SF*djp�<d�X�4y�������t����w�Agq�����~��K���7~���NzE~�HY���h2�7���rZ=��a�]�o�2�����,k���m�cV9�߬�'76Y�hm.pϫ��Pݶ*�o`�y>���r��e%�y�͐t%� �V�:B�6�I|��9#�y���@N	3^T}x��i; ų�ÓD����5�{�!�l��彘,�^$�)2Ī�uV�M�M� r[<�A�J��`��ŕK������J������@�N	�^��
4��Sww��3�^[/���ӄ=�8��I���Z�:�����������>+�X�����:�^�u[���՝t�+�48�b�/��	>�N���SO�)�&9�5�~h+e0'��m��R�C1��ٌͨ0���z��A��g�y��������@"t��q���z�7�\\��Ū��Vḧ́�ך�_l{�=�$�ު���j\�J���r7������f`8@�V�	)OÐ�V��d3�ن�����u]�P<m)^i,zlp]��v��{Iלޮ�n�l��gA�m+���Kߺt��"������ϻ<��2��	x% R�(�<�ly#�I=�)!BJ�א��s����2�^���A��xS� P���o{���?��~�����|K%��M~W�̓���0��F�Эƞ�j��e{�����@�l��l����]e<�}'H.[�19{xh�gW�z_���
�0�y1��؄�Z�W�ZG����f.���X7��X3#b҂ H�$s�x�i&{���3k��!^?K�ٔi��@���u���:�6a��#^6�x[�sU y�V`n ��y�P������h��=�f���\�b���m��	˲@!�rBNdS����̣*��|�K��]$�W�����f׍y�z�c�S&�������خ_���[���ӱ��f=�����}� aW��e1/�<$��{�잒��!�Ecm�׾�\���@+�2��<	��$���,�v_�쨧��K�6�MX�/����ֵ�][�_;����@�/k�}���~��x�ǟ��vcٌ�_����o�=K e��6�~Y��� MpCI��n͢�Sbp���^Y,(@"F���ڈ��LP�H �)��M�3�،G�{(6?\1�q[�G�H��U�p��9ҿ�h�����8�8��=j�w����!�c��E� W��8O�#�8'(gP��T�<�R�0=��~2��+ǫ{�=���Q�y����~��﨟�9�����Ͽ��?�����"G4,X����C���IA ��۵J�ԇ���R�^/���O�6w��鮘�mB�:�D-�	�.�V>�sQ�Jzh+���R�2]�!�ILloߋglZP?_��IU��b��EO*�����t �4r��mU�g�{}�ȉ�h۞���?��26�5f�!Cү
�MR�Q�Rd�3��n��{���K2V�,��V\^6<)�L��Vۨ�ruh�S �U�d�3 ���խg�!e3D̨i,:��յ���޻�cܧ�g���ՙ��z�F�9��SztC��9z����~���M�A ͞̳�1r�������WkU�|4e@���zw�}-[�;�-���}
��]�2�Ț 9����ģX�0���y�\�|���q�����#i��n?-g��=6�k=��n�z��X��kU���4��"�%'L�	9%;�`�L
挤�T9	@�l�Fk�4r��CY��
z���M�B܈�\�H٣~�������zQ�p��������7�����zU�Yn����n���zU���{�*m�ל���@��(Д�����7�\��mJ{ ����ɟh��}���aqޤ�it"�~����Ư��q�����OO	��1�H��֦�^A����e�B�aH����#T�k�]M���C�7��ƚ�G��.[WF�yzŪ=�ݳ{�_�(Z��Z�V��Y�_���'Q�VJ�D��Z����3�0��t�6v�����"����)ﯕ֜��ٕ�n�9n����X�g�W�ۡ�s�.w+�:Q�M��s���e��+\���-S�n�qy!x��@� R=�n��j/SL)#1#�Aa�2RS�g��L4[;���抔3���L�\@<�6����h��q2���zR�b���M�j�7����Gd���{�CZe�EٚK6.b�֘�(2sF��BW[ߍ�
2�L�T��y���!����sF+tqt�.��y��@/�Z��wz�Q<�]O���zM����Y@���U6��d�{�Q�p��l�x3 s:o�!o����{�Z��li��~�4M`2�k��b�dbO�JV1�'�ͧ�l�*���*cؑ�v9EWEi���O���Q5�e��`|@�����ݯ�*�D7��X�vO��,cF�f�z=Ł�ߏܻ/w.�^�z:]�L}w6c���{p��yO{����0s��e������ `�(~���ެ�it CB�s�(�|]./~��<x����0��ݽ�q�k7�M!��湨����z��u������X���æ�lv�&44���%��t�9��#��4<�ѿO�屛��L�������y�Խi �40��v��`$O(��K��;�m�%v��IM>��=3*(�9�++	�������ٟ{� �:Q�W�JU���QEէn	�������Z�
hJ�1-G\��oy�Ɗ��ZQ[C�L���PB.�zf��y����&X��V@����ē`i���PJ��eƝ�~���W��&�9�f�mk�p�)*�zlN{t	MҪ7��w�Ev������aHٌoej���v;�a�r�l:�P�6��&���N;H���A@*;�i�@��'s�tq	=��.�8����Ji�n��a3�'7�ӣo�`$�\9��#���l���#2�kH�+���p�ѝ��Þ+��I�^���}�Wd��[=���m���b��n����N>��B�x��-��V/n�����G�9m���\�\zAl�
jd����å�>i�H�!��G��,����U~�������H�)Rqs�~�	�ŏk�EG�f��;@��kDJ��C��Ɣ����2퐦�T&�r���i�������S�����7���M�M}�w����s�(>����������K*�	Q����˧���9���e�ՕP��=r`�ʔ,TBCAZ�^�Yվ S?�W�����z�h-�R�ԳC
O���Gچ�\�]�F�����Ⱦ �(�a��B��@�)���j���[�	9�0Q�!gܚv��.pQ�8�=&-��9!��vJ�>'�Z��ۃ��d�ѣ��MW�z���am�{# *r�P�̌&�|D�'���l��{��	g���A����V.�Z��ǓU�i��3�
�Q���a���	mO(��e^���b��dnD*NMq���'2���t+cAc=�t1��}3|��^�E���t�Ve�*���E�x��;��}^wJ}F��NH��9���=\��&{b��кN�y<�i�`KM`�ВВ��!*�߃�'!w��g0JbdΞN�ϚR�y�<��7d��(�ի����U�&��[����Nڣ?�Ag uY0��=?SA��K��郡l*[�N�
�� M7��6�<��#�,H�L�`ڡ���&�,�V�'IR�tEj{��p<][$*O�i�z��CS,�tid�r;��?�z�9���"M�������[Ov�)�S�Z��E�v��6y�.��3aҸX#�}��+Fl_�}��
'���#�����-��:X��D�+�?��2A��\,���`���:�>ޖk��G����S�7�o��C�3�0n������^~��9ܯi��+𣤺K������|�%՞�@nM{ۅ􇗺����V����V�@�W��X���K��m����xo9a��Dmآ�E���ƿ�W;���	9��5�o]�@2#%�BJ�����[�`���T�����3i�e������%v(v%SvO P����=����U��>%�BA���H�_o�̬Tv�DBDJ�oӴS����'䴳��4�ݑ[���Z��¢�V�dJzJl=����`�k(�C��&�s<����&03��Ќ�)�J.���-|�Kh�Q���D6��� �	�+�d��'2�'�����б�������Ƴ�j����ѾǤ;����/xލa߽)����?�+T��n#]6�\lP���*H:���(B"�5���R&P�x�M�4�����m*����S�˧�r@&'�V��o&���5ZU��`���Ƭ AM�A�H9�%e&eb]�E[�*M�*n����������N|�����M�D���'�UIDIUHd�Jċܴ��}��.��0�X�R�)_�̱��� ��?y;��3)Ӕ��_@�p�X�()�	cވ�Z_����dެx�@�!���RaKM�}��M$��IU��u5�!d�(�5�;F��(���F��7������7�S'=`�=#��h��SA�%���r�;�:��ns�3���j�������\��|Ͽ�����?1�2: ����_�ٟ��˸������{�=��$���酪���k��+���q�����f�KI���ja\/"���zC8b�=4z��r{@������G����xiKtE'�zPTm85A�#�d�c����>)I�"��gMH�(^�iyfFJJ9`��\pk���t�|�|@!k� '$0)Zv�>�����������S#JU�-��DG"����> ½�t���!�'�{<pՓ�^K[qF������
9��*�*�T�lҞiwU���v��}-�:�'ngpR�Xt�@p�GiIN��2��e�t\x8N[D��v�D�����E#B*��pk���-­���.����yL��X r��k�ivD�2���MWA���vf����^�E���Y�U@�!��. d*����
��Ҿ��4%�\4��!�"������3v���O@�L��K��'�O�佧��̤��&�ĩ1s#BUEm�.�<SJs���r:��� >NJ�>щ���隠G �rﵓ��"h'-j�,`���W��(���p��C�])�n�����>�|	�U=�&��-mr)��փjۋ�I[+R[��L��$���"�T��HZPX�XG�\���).��)��@�KL��Φ�ժh�J��Ac�>TB����H��nl,��&P����=� �
�V�Aɮ��;�ױH����}���I5��u�g���)#�؝��*S�g���X�H��{��}�E)�K��7��v~��,�Q���w�9���G?���
~���=�f��˷ԁ ������+��q���_hy����m���<1��k�/Q�"%ki�&Hb�0i�N�:���*&X�ܛ��x=��hxI8������V7�U�C&`l �U`Q�PSA&��V�'�W ~�0)R�P�ȔL�L2�0�f1QA��r��i�;�ܙ�`���<!���VA[`�ښ��Y����T���<�Ӄ������5f�� }�2^d�<����h͉+���ݾ*s��n���ҔX.�����2��r��Sʍ�y.Rk���&�eB]
8=U�߯����wcW���������T�E�ITx�j���P�'n)�4/x���Ǚ�JΦ���	9eH3)K&����S�>+n���pkG�mFW"D���+����}��6̨��m�.o�J]ꛣ�^�lm�Ex���~��Z�.���. �Z�����	uf�(�H�V��݄S�q:	��)���gԚ���%��ٕJ�n/|�����S��#_3�Cb<,�����_�į xE��,*ߨN/��[.��[ޕ�)7�,�rc��D¹4"m��kd�e�&Mx7)�De�k�,�jEz�Qr��m�@��r}dL�y*iJ�K�Xu�mn	@Zj˵�,�%�9Km���V淋���R���|�H}mym~B��Vkˡ-ׅuIB�mAʌ�����q��i�����B�N��]ɸ�`\��КE2
d)�vB����hb:]��HPP]Еۈ H��u�Ż+]�����dE�"����Q�;��'�#u�BDS�;oM�{爌Z�q&�a>�@0{�>���>xe�R�#O{�2]q�-�������������R�9�-x�v���Ox���_�{��Oѯ�ҿ���A^�E�� -&�)&<Cb櫶il��R����D��dZ��\���lz�{��f����!���&N��@2AQA3�넂v���z�����+de
��M�1MH�=�N9{�3�JW�c���].pw�w����z*C9!��Ҥ�,Dt��&ί���Μ��S�\N�O	��*��9O'N��ʇ%]ޞ?�3?]�|��r��R3���֟Ih�J���n(������-���Vlr�js�L��'���������9\\�5��Y�q}��YQ�KD�[k���i>��c��[A*Y/��P8=��J��e��yλ]�23@���5��ä�ĉh_wD�/3������?����²]KοNە�9���D�`P���F�1Е�[�pV(�GE�B��:V��� �MՆt:i�_B�	����Δ���K�Zv;�ۇ��R�I��x�s�j��P%���y��SO�r��xI�o�i�Uʻ_W�/���
PK�%���VJie�qj<q�����7e��[,�"��y+��v��	�fc�T2���tЗ#�X��'kgj3P��5�S�L�z���Pv�L��Ί4�EZ�5H���P����"�a������u��Xj�3Z�2�_��m^^���h�۲�g��nk�����T��z(:CeA[ԥ�-���e9��#)���.�*{Bk��:5��m� ���־�D6��SS��' $Ӽ��l�J�#��vng�k)��0A��}��1 h����n<EYi7587"<%��Z,�;��R��xJ;K#��W����^*��J���.>��[�����-w��K���>���4�˸n����?$*���/u~{�si���fH�!��0���n۵b-�=�
�<�����L7��^ �ʱb���߱�l	�W�pya��������+�
����`E6jU��.�֐S�R2�2!sƄl����1+ Ta�
�|�C����%����gO�6����v�2	8w�_Ki����/�gSΟL)����IR�s޵��V=<�T��'>����z[3CiBK�' �g�y�o�z��W�
 �ZѤbYf���=�����^�ƽ|��5?|�Wi̜H[�Z+��L�-;�tGTo�����E�u߄wJ�������rI�3Cs��I�LXTY]S��'��Ki��T�%����z,,`�jR�["�*-��GA��L{�`�-�z/�C�T�R��fPv�RR�uG�}k=�ѓ�Px�&�U�[U�U����Y��ki���R[b�K[�R�)�:/u��~��ݾ�P3�ք_���|Yr������?�z�g����4?q[�p!�ť�|K ��}�SH�ۨ8y����l5����5���?���x~���  �IK���eF���!��m/����y��Nz���г�������;�����<�xWP��@��Y󤏧X�+d�RL�XeW��Rk*��tD=^��%��i����������R���f7�Y�t���A�0N��st���6C��P<r�3�X�\� `��X���/�6ʀ���ƞ���P&Fd��N6��],���H��i�������N����������Oķ� ���G��w��~	iaҧ����.˿�d����&�TZ;B<N*�y7��f�M���G�X��+?Yŧƞ]�.�^A�!�⣴�͏Tتe��ײ�ի������z}�Wu����
h"̲`>��Dؗɫ��r�dNإ	S*&/��g�j�(�w8L�qQ.q�p�������S�Ň��ʴ�r�ʧ	��=�_�����WN��i*{-��|���~���r�0��	���	w��^�w�RI8=8�x\p}\���}������Z�ڽ{�ݿ�w�S��,���=,�	��D��,hMH�uB�ɋM�D�o\1e��.�rb�2A�k�+Q����c�i��~�wW�ֻ���-�N��d�x޷$i�95��Ě�sK��wAV��&a�=0�o�{�M�7\!�*)TD�6�(�q�nr�n�r�ׯ<���8����^�_k�
�gk��.tw�6P��2��O��/t~�{��S�[O���3�[���ew@��HE��}�F��7z������~�+XN�X���f`>bz�I��5˼�\�$e��I�i�z�b�E}7P���4�ҔT�����j|k�C�j}�&�,G���ꅔq<U\_/&*����4pݴ��6�c�F}*�����T� �#&��Z�u��Zunqs[|C
ٍK�Q�H�����5�m��
ǽ��vS!T�^�m�ZJ�۾�T.>���.��?�����C�,���#o�R�'�[�@���/�P2�_��SU����j�ai�;[��&kaZ���R����pk5�9Ϗ�$x.�+m?��O���#޾����6�ի�{�+|���k�W���Ҁ�r�um�>�S�������*6PD�]���p�i��~qUP+ �q��;�{�$��}Wn_�zpk��������y7}\���~��_�}��اtwH�����l��t���^���Ջ#ꬸ���)�N`͠�P�x��5�EЈQ�RFk%��u�_b�9����6L��z���X��^~���p��C���ⷿ�{s�U��g>j��`��p�O?�=}j��km~?D_$�}����\?�;�F�|��x�,f8���"g�����Ԅ�i�i^��+�
���r��;>&�%&y\=�]�pm{��u-�+�P�yʜ���M�Ȥ/{�ڏ�o�~��P8%3+��J�B����bG)#s��8�\v���)���xˋ|���?5���Η>�1(	��5�O?��?�aY�����I����iE�I[��XߢV�0�}h�o�ӽ���X#U" �/���i�-��ke�"�
WU������#��W��'�bC)���QR���(�$L����!>�b`�&ȑӄ[��ؕ���jŔn#c�D	�/���~�ٯ=y��������n�����ҧ_���$4��sϾѷ4��B?�a���{
����an3Z[px�����{���%Ǉ/��J��K��Z�k���bAkC&��^�M	�
�B8͋�N'@��i3/W�Zsx�����F%\�I���+���'�9#%B���d����)���pLލB��Z�l#Y}��	 2��4ٰ�4������k9��J�WA����>���8��-��7�������@�/|�ؽ�i\��h�G�y�����^�N��wf�ߩ�h�����Ui{�Z �Td��^��G��7mܫ��#��f���a�
}������J׆������,*�#� jC|��I��WhRQ�u�K���%d6�f���i���U����\���w��;O�}�c��̻>��/}�ݓ�s����p���7�6A ��_�E �VA�3�y��镯���t�.>Ȍ�6ײ���{ҖI*�r�2� ���s�>m�P���ٔ7��@��xS����]�>�
U�b5�UKIu�����e�i�GǞ�2��qA�x��y+RE`���{ΩW��(/�r?O��r��/Q��H��r��;���/E����=�;��O���`y������SO�vz[m�gAx*ߣ��Է�ջ"� �C2IUXUX��h��d5�㒮��R���Ůq4%+a����{�}�EM`B\���� �����MLPb7MP.>�E-4�4�\�����������������O��,������e���[Z��?��O �^�����>�j~��[o� <xG=]�u��
�>��{���і;m^��T8^�Z5u����54��mmV5�&�'o
�v�k�z#�����3!�U���(q#2��ܵ!o(��p�˔�g��I�.�,̩��2_'N��k����?���?���^�� ��}��F���t~��[��?�ҳ��P��׸x�S}����[h�Ro�N"����P}Z���[*8a�������խ����c_q��
���7�.?IB�,�m��*����>�0��וf�����m���5-˂��Jɨb�1S.Z�W%O��������px�s���/�{�ٷ�-�<�����o�� �g�ԧ���x�|��� rxn�,�����6�<S8�J�U��o"z��o�N�Ts���(��yO
�jz6O���"������
�6C����ܭ-nk�$))aۤ>�i�2"��2%%NB����J�f%>�
����K�ӗ�����qY꧙���F�^|I_��R�L�Uo{���ѷﷄfw�/|�v�j5��@� /����#K]�&�h�Y[M�IRQ6�g"�邈n�-�iOL;UL
ͤH`Ndc���X��J�d�G�*T�`�FB��5���B}�+��De�8-3��#�*�2�~�'�V�J�����<����������O������/�u�4��|��ѷ"�JT�}�8�M����p��~�N��p:ͻZka���:�D�ۙ���������nI�Q�h�k�y^��T91133)"�b��f��@�Y�Z�\r΀���W��X))1	@ں�-�1QQc�
�
�3���9�gN���U��N���,���>+���S�S^��N������¯��'�
�����w?�Y�؏��}�� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��1�Ӓ������   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X    IEND�B`�PK
     ��d[d��   �   /   images/a262aa33-74c4-460b-b0ad-c746896f6744.png�PNG

   IHDR   d   d   p�T   gAMA  ���a   	pHYs     ��   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X  �IDATx��{y���u׹���Z�j��ez�����L�b'������2�eH$BaJ�@�dC��`�@��![G6NlϒqO{2��=��RU]{��ۿ�����1�'��n�u�{�[�=�s~�w��ʥ��1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�l�c@�a�z��Ti�R��)�|�H)����]ǧ0�Vg�¸K�F�Z���=:0��y��8L^a�&����4�"ϨH32ʐv4������>Y��6����=�n� ��w�H��)�~�����t�g��!�<T~V�Yz`�����j����ר�����Z�:@N�NF�ޢ���,S�ޠ��NY<�Zk��J��� m
& ̡T�nW���]����{}*f��>s���m�ݽ㯐[����u��)h~�����>�����R����h_�М�NݴC͠���ޘ�g>�?���g�~��P�R8葉ڤ+�T�O�8�,�`�UZ�	!�n�6�a���y6O"ǭVk��D o�D9~G��[�m���^�u�'^"�[^���O�N����+ DF�u
��v�����/M2�P���&���8\��
\��w�z��V�K3�K3���h㇟|������~ݟ����W���f�ȉCD�M"�!Y֕�.���n�Sf�	ch��G�&�q�H5���*o/��%�ݼIj��KI�Z����.J[�(�\ׇGk2�j�4���X:
A�tԿ�M?�Yg����K_����pkC通K�23�*0o�g3�$����0�v�g~�/+�W7��|��ּ�,un_����� I;���\��u��_},�~�n@"��-ob+b�v��X�I��f�L]�Һ^��U�8�E'?vV�x�C�k�;���M�}$�DLi�S����mQ�Ņ�:��(_Ug�����F�����	��ġ`VcrDqf*��q
4SU�NLm&U^�������G��i�8�3�.�۩.tؙ9|fp�[�D����W)�lSg}�����ѡ��0���%�]���pa�[���>PD���~󧢵�� �v���ԡ�����?�j�UZ��ε��@��_
��e���,�=McB�'�pt�&���.���
{^�K�zst���t��I��#���\N������r���4a�8&:��i�M����fS޻�0�*N�� ��%
V^��'B�%���w�1�@��Yuh$L�wQ&�0�3��	B8f��e�wA���Hi��%�?�p-,$|M^�0$ln���ÃN��'���S���;u���}���~g�| ��eP�>Gӧ>�����)3���I�+Q$d���򼴍�*ձ�aѣ�x�M�"D�ܤ,=E��Cdẝ��HKb�=~���kur��0!�-�)���!��D��)�px0D!�`����!��YҞ+sU9��x�T�J�,�OR@do6v�"�J��:������gB�K���E�����Ԡ?±��� ����s�Kh���+��7^mn����&]
wV�:{���i��u�Z�|�I��'��&��=�{��֠}m�r�<�r � ��c%ED��*�	���8k�0�Z��5�׃S�w����i@�g�ׅ�âz��w[�D'��I�Ar<��a�L*�އ\M����G�+�+��߰s[�����
��T�l1�z��=��.� �v+r�v��[�D�KO��c�	�K�N����[_|���S\�m#$ł��y��s��~)�oR�"�qm�ߵU�/�ԃpw��
"��U��2��Nڦ�<���w]B�^�X�U�F�ozZ�3d��(w�m����&�ҳɂ�d^J��)$��D� ]��X0�*\KIy,`Z�S�oا\G�څ��k�ԫ����G(4ED�+�i8���\r;Y_�Fa�bn���V�`���܉'�n��z �}G����#7��{�B���/ga�`:��v!{�%Z�A�q�P�w���~CYT�UM@u�C�D&�����m�O���KY`��Cs5�e@Q�f�\Z�m��-�%*$4�H`ٟ�i2WD�L]VCq�)�~�dQE�:�)IX˵喝
��O=E>U�)��:[[��Bβ�saȜF3�`H)E1��>>CN�?оs������=��;k�.�$�ҩ��x�~���p��_Α7�p�&q�@NTNu����	yф���ά�K���	]�WQ�6���p^S7����N�z��7e�WY��G�95�F��+�ÁBሚ�t�D�,UX�/��p $o�T(M{5�ր�2�gBrNa��r����
�7_׃s̟z���S��\!3X#߳�7��0��p�3��<��D4��Y���b4~�:��˝�7^�H,P��J�ܰ�K핛tv�y��'�w���y�����a2UNQ��8���/#z��!X�4Ee�w�.���9��� �ޙш���.U�5rI?��H�>��!���~�
S%6Y!
F��[ͪJ�亢�"PNтĚ�Ҿ��\�*Ȫ"�윬c�*#��%j��}���y�����﵌r+���Q����5��#w�<� o`Nٰ]M�꿞=��3������i#$�z,�Sm��}ݕ��}�{���ޑ(P���̄ZP^U<P��7�E�)s��p� �Jg�"L��s���8=�8�&Q&	�A@����d��U��Z%p@ e�w�C�� jT���xbn�[惟^��.�ӶxmhI�R�8��X[;��Dn�E~�^��WR# j.�5�RX�_�r�+��]�ʜ-��"���^�t늬դ^��G� x�s�⿸���ԉ?��Q���:�o��� j���g㝫���8��/�(���E�a���r��j�Tܻa/k8S�PY$����I:9s��;��1�M��0RE��<�Rھ��DR�y�2���D�*��$�ETdF�(�8*4�uD)1{6G�����@]-��=F���r��q����0��؜(y�s����@onm/;1�y�&�'����YH��.�KT]xP���SY2�A9qE���	r��������������έ����{>�����@S��/�c��eu��ʘ���	9%�Qڪ��x�"�4a�$ۡN�o��t���"��Z�m�O�ȉ�/SmΞ���%���b[�Ap�����29?gi�IH+�� p"��� xH_�\U�#�8 �=���� �Ʈ��Π�P|9�G�ex����)ݥT�$��5����)L��H��=�c-9Q��3�C���"��BS��4�=w9Z~j;�~����i�ě�}Ű"a��$�ڝ{<��X�1x;"g U.�*Y-���$�0��=��FG*��wi�f���zK�l^���~M��!t`����E�ޗ��5@���R�3�7(T�rl��<��T��;D5�PD��ѹ���d����\�p�!ё�I�#&��Hn=�Afa������[�M�����ox(�}��jߑ5*8�ҷ��D]�kduƵX���E��e��g���s5��w: +�KaS��q��0Y*rc�dZR��+J�*�G�Zc���"4A30��7���ޯ�Q�/�޸D���xs��D�p���.a����6�9%�3ա��XYn�"L[�˭"� �� 1��MR��(a�F��Pcs�6���w�UD#�ƴ�k�:&g�ɻ��P����]^[U��գ�W�s�%���@X���f�S�?��:	���.�B�r8�魐��57�ڛ'�G�͢�k�$�\.�Ӳ3�������|�R�|�|�܁�ڴ���P-���ץ�+Qhlo�)�^��˹!;�S��1C'�aT����Uz+�t�$½�;j�9�d(t��x����m�0H�Հ�"�Yi��BT������5���8R��/6�̽L�FKn�M_r;4��<�\�؊K�E~�%ut���ص;�2��e�@4�����*kY4S���X/���9������
�Y
p=���8�8,Xp��ͽʶ,�{F�>Q�H�Q�Ĩ�SCsnF���g���T���胁őX���}d�$PJR�_Ξ)�
���֠�hGh[���j����'M1��'�>�Hd�D5��8R��,
k"�Y!���C��\Ŕ�AqY�(7��=�b�H�Kr6���e�Nو+_2Kc�����]9ڪ�£���a�Y)@+[3N���?�u@Y�I��2�a^I
��a�|&R��e/Ki�Y����������<}8���$i��{{*2m��"��ZjF�R9\ c�YZ���V�#�j)y�*j�Pj�T))6�����Q�Ƥq��(؟���Z�K�כ�ό��bЃ�l%"w6�s9j�k^\	�m��J� ą�|�(�MҜ[_$9��.e�h5e��ؾ�eJ�F�M0>ߵ�����C���W��4n�&8A�{�^�U,|^x[]��~{�/ۓ��S���r�*��VM:�Ibh*,J2�{`PY��-s�&BU�S��!b%f6zx�"(���u��_NM��ϯ�]	p���[ِ�������C(A��ʚ�&V�%n��Ҳ��m��XZ)�77�lH>�~X���w>�ⴇ�P8Y��e�z��>�!,�S�}%�[��˕�P$+!g�0��Qd�F��-¬��X5�@�iPE�vٟa�T�r7����hޅme���-�a�����Ɣ��;GМ��`��?��{��~�ɿ��'�������C�r.r��Hf@�޾�ѹ���J�ƲЛ�J8����1��� B.N0���=6ۈ3ei��0����E+<÷�V�sI���ϋ{=)�[Q�����#�Ap$�r��q�a(�`�FQО�Y��jî1��X�~�ʍ����C��V!��e���z�3�r�[)W�`�'��?�%��_x���gg�~�Gk�7l>�UH��E�ǡ.J!�dv��:�Ք&�6N���&�1�Ri3צ��=#*�!>�
�mI��P�{�0$j����쵲�ABf�Y֒#����j�����K+GDA�iy_dv�Q��M��T�b���xm.��P�vű|����g�e�X:�JP�W�})B����qQ���H��=���t{��?;�U2�1�	���`���'�~?l.���!Q�w+gD��w��<F��8� ��#$�I�G^�Aa)�un��-O!
c�	����ԋ
�	i(6;��R��	�����|#M�RJd�sRa��
VO^'ANL��Y�k���PY��6��Z��<mMf7�4�t&{,E)�*v�t$F[��1!,�Y�y�s������}2;7YW�����c�q�u�x��T_,.y�}?}�y��,�Ӱc���Z��团�`����)&��|,Q�%�3�Z�T���OD�R����M�όy����|DJ�s�<���O(]��Yx�L�|��X�ǀ�ANY�ؘ 2��H0/n]��z�̍�s�B$+D���"Ys3�T�
Z9?�`NY�h$�(ͲQj�cIQe�_�)��T�~.�t�̳�z�U:�����!�����(��+/�����_s���n�E}��P�{o�����\P���r���J*@S)GG����Ae!ȋ�G\^���P4l�ݞO��+�;�,�}!<��F�R�L���=T`��v������[C�����8/QV�I��@�[�%���-s"� d����uH2��<�P1��:h��gI>�b��I�ѯ�Ch5�������7���st�]��\�v�~7-_x�K��c����YtH��O�-��:�F�"iK�\Ŀ�׏���4�ϐ�x��
�d���Y���Oi+���V���!���h�w�e
 Ң)�;�YِR;@nom��@O���#&���V��UBq���ͯE�.E��4�΂+�5YO�{�F��`d�mp_>��A�Q/���t���h�(��;�_�Ï�|���|����k����W�n�u�1��H꿡������H1��;�^�[��dQ!G��Ȇ2�@qN��A!)�k�ҶVE�V��u2��f�u�k$xn��(0p��]6�F�DSFF!^���+
��l��?W�yn��\Ԡ)v(�6�r�u$��k�
PEO!���$c��'�,]
�Q=�st�t�\���ׇ^�������yo����G����!�v@fg��k/����?���������S�ҡbЅ��e�~i+e%BVG��b�f�n��Cb,�N�w���Ƚ �T�k\�K��'���V��h���]�B�� ^�>]�����lM+�wJ�2u������5)Ly�2�MR�UI5�}��L��k1����k�	oN9Vy�߇�#Y1a;T�&�.����í�~��c������c��i���?0��e|�)�u�T���[itď��FC��'�Oūx��i�\�s����3Μ�-���'���*��jו�6$���-��4��"k����z��J�Z��sը�Pvo]B5��\Q�{߳5�[%g��ٽ)8�eC��0�,~F�_�J��@t�4U�*(�R��#��>�M-�hQ�3�܀�t�m�e�l�a=^s��������~�wx�̇�w�������K��|�vV.��}�?���?b��;����"�e��=�f/.��kT_���En��u:��!j֏H����V��|W;^�K���MD���*��4���AUy���Ss)�f������|��#;���.�u ɎHw���.!��#К��BZG�����8�%��N5O�zGSY�u'�}����O\B� ��Ȯ�H�N���a�'.j�.Ҝ�g)�#p+Ti-Qe��E����a{c��n.�������ճF��w6�S'�������:���H�}R�sn)���>���z�&�3�Uϣ�?M3�����Go�V�3����W_s+��&��N/�G�+���Q���Yz���k۝f�f�����@{��㙄�"����Ju��9�r�i�v������������X��� �:��LT��N{�/)<L����l߭;�f�y�5����ߗ{�<r����.��y/��^"�@�ZI=�F?s �<8^0��U�s���t�s;���H�}oJ��y�V_y�q�����d�����~�v>��n�%G GS+]A1��4��x*�������D�ۊW�=W��k�>��/]�򯷛G���	��P�_'�*�.kqgv{��RoQ7�d�*qR
}EQ��0�і���|�>9Bൕ�e2�-�i��,�bؕ=>'K�w6h8�KG��� `<PRvP<�)���y���?�ɠw��G%�:��=SSt�0Eu�婙�H�Z��S�z��M�yם��?[�N����s�<E5�X�����w3���}ȁG�CwΝ�J����is��*4������V��6}���ȼ���T+�����ڌ)	w�9�_����W~��W.�C��%ZlP-h������}/^�L?N/|�b`|P��֚l�nܜ��U�y�ؗ��ڇ2�[��}�[����<t9`@K���w:�W_���BՇ�{典H�o�4�f��2-��_���[�p�C��
��9.'u!\1���tz�5|�|��>t���W�9��D<����Auߙ'�~�s�"�?�7i��D�����G~��_{)�]D�D��.
ɵΦ��j[Mz��ץg�͆t����q����r�N<�m�W.~���CTi�݋�%�W�ƉluKu�P����FS��5����� ~i�~��wt�?�}�w�����O��O���wf��c�W�c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2f�D�{��w��    IEND�B`�PK
     ��d[�c��f  �f  /   images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png�PNG

   IHDR  �  �   ��ߊ  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  a�IDATx���|SU���M�M��ޣ {��Dq�����~�V*�~���(���(�"{�Q6-�-�M�{�'I�M������K��{onn���cU{�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!@��-[a츱�aC�5?�q8�^ݺ"���0�
�"���l�a���>C��p���Oo��vn����"��mE�9F�1\���?ۛ�����(:���c�X���_wlP(�ʔ{���=��|+��#}�Y��mo�w��k��]�o�������?�O�0�?���'�Q���W?s��3��"Sڶo�dՊ�}�I���i�f����gf^�t8Z������^d�g`���>�n�q�0K���k|=Ϗ���5�1��}���I0�p]�y��U��'3r��~'_{���G���ߢ��h������1o��v�#�����޵{�I��z�}Պ�ged��x0'""��!;;�߁�������t8�ADDDՎ��4���N����E�l4"""��L�����QQ���ԿTP�UK���	���sn������BDDDՓ}����{�������H/�=��|!'""�c�4a��sh׮ݔ�#F���u�}�?_+.q��p8PPP��o�O���m+�p���DDDG�}ǎ툯0;+k����C���PA܉��\��+z��I#<r䑓�\y���O5�Q�?�^D��R]�]R<�5k����q֦=11Q�s�*Yǖ�Ull,���0�C�Y6'"�`V|֠g�HKKS�o����T���Ύr���������GXd$���(T�:����=3+Y*��D�~2+3K��H�h#"���sx���_����`:͈�����O��;r��"""
f����6.��p�)�ggg��oDDD�����R�7Mgx�'�����"""
n�Cii����p:M{�'��]��QP3��SSѼE�8���,�3�:gOݟ�F��:�������y�
�DDD���";+;ơzI2�kff&���(��j����H�4�L��at""�`&��:���K@/3�^�a�Љ����nC����E��J膻��0���(���*w�^���(@VV���(���*����:��D^^>���(����p�Yo`� ��;w@/;�����FDDD�Mr�0��mPP�ϵЉ����iB��'ԭiՆ.������Q�V�%""�Qt/w���^J�&�΀NDD����m6È𶁴�{+�Qp�/^�T���t""��g߾m�*���6�Q𲧤�H������]��1�'���i��*w""��g����m*`��r���/��Ä�m�����NDD���3��G@g�;Q�S%�Æ����˝��(��3�����G����ΐNDD�Lس23��i�I��S��)U�ge���'{�3{NN�
����%�;Ճ������zdDD�i��K�DDDA�T=&&Ff��Н*�;Y�NDD�L{xD�t�S�:M�~Q��l6;|T�;�&L�Љ����=L��*w�Su"""
^v�a�ax�&�܉�����0�QN	�U�DDDA�T�\J�׉e���U�DDD��.K�|tV�3�|�i�̽t�U�DDDA��%���F��8tV��rK��U�DDDǀ�����t�K���˝��(���K�z���X���(��E�{	��7���t�,��ʝ��(�ٝO	�:��:űʝ��(hI����4�r��YB'""
fv��a�iz	�n?7�)���(�ٝ�sm��NDD��r���SQ�n��^�n��GDD�쐕�L��T07Љ����)U�J8|�r�Nq�DDDA�n+/�K�g@����<����@=?""�F��0;�*��乸ҵ033ii��k�.$'�@jj*>�����9	�QQ��S�ѨQC4k��6���\���1%>�|��%rpq��+�*3��?V�Y�?���Eb��-طo/<���<W�C=��,|��\`�!6&u��C�V�ЫWO0 }��A�&�f�1�Qȑ��i[�I@���p�{�W�܌���X�z5���;�:��V�ޯJ��(��Q�w�{�>)ͧ�Ė���/s0i�$t8�#�=�\|���ܹ��v��D$<�����pU���Ʉi7`��r��s�C��\�U�^�x1�����n�n٬��E�ۆ�)����`�E���Oq��W���GR���yv"��\�g.~��w|��g���;п_?�i`7нN��¹�}�\�-[�b����Gcǎ�p�W�����=轢������i�O��P\p���������O���u����拓�'�S��o�T!����>���2>�͘����3������_��p���T�Y���tf������ذq#��nԉ�cP'��'������ix뭷�|�2]�Y�^�z���'��2���V�{!�Pz^�0���*RS�µ��Gݷg��g'a��Mw���������{���#R�۟���#G���x䑇Ѡ~}u"
Zy���7o&��f͚���8��yHo���;�1��&��ޔ�y~&M�\�f��`�
���hܸZ�h�:�E˖z8Z�*UGGG#7'�z8ۆ�n�:lݲU�TU�[�Z�QV�a����HOKǨQ#� 1�A������K�,��߁�����Qi�tn��lC�C�����g�><����!??�oF׵kԸ1����3���&M��v�ڈ�{o���b�ʕ�a�:�~�:w���Gf ?/~�$��'�@LT�:�Ca�^��,���eʐ�0���or�gf��_�G*��`���9Q'>�>n��V=��v�Z�ϖ�|/C:�5i�H?�~n��L�<S>�\��S�5��s���[h׮n��z�~Y�(�2+&K�"��n�f9U��W\�Á�U	x���s���Űa�p�9�v\-�_+Ƴ�L�׭Kg�;��|2��֮�ù�J������ѱc�ؿ?K�DD!Nt�s����!�{Μ_���~�2�M�!����#г[7�_+O���/�	u�b��aX�l)�36�6��ѥK�� "�P�c�i7���*w]-̀^�n�ꫯb�d�z��L����p�Wb���hռy�Kƞ��u�@����~�H޶�����{�	�_xK�DD!ɕ�۝�i���q����0��)���_Q����p�����FTI0/N�}�Yg�����ǟ@���(�/3p�@*�y�m�4` ��cP'"
9�����rg��#���,F�9Y�.;ѵ[�G�M�VG%p��,2����/�L񲕁?���?���%]""
I�L�곛�k�Ԛ]B����i_c�jo��L������ރ^=z�R�'�N݃~�os�o�X��3��0s�L�{�DFDT��y�"X�X���x�����X]��:Ne��.��� ״������͞�}���[8�2{�u@|�ٸ��K�ɲ'8�w�{���O��������m=�c���xbP�p�ٟrss�����f��u&"B=�ߞ��y�v����y���Cn^���OV}���a+���N�[�8r��!�1�(ǲ��V�Nq�|����EFxȹʵ)p�>[u�rm��ץ���u}]�����OC��:����9�?���"��\}��ˌ���^��Пc�{�hU��)}>޶�R�5RT�y�s�C~J�@~�V�,�[9C�����57"��_@��U�?ϙ��+V�ۭ%cͯ��zԍ�?�7�/&:�^v	�M��C�0���-lطo�-_���Y"v���X�vV�Y��6`��]f��S�P�,�B�Z�ШQ#�n��:u�q�uD�����JZF233��]ۺ		:�*�>��)�f���X�x֩��s�N�I�##"�{hѲ:v�^�{����k�}^ŏ�r�*,Z�k�5۵k���t@����36o��{�@��]о];Ԋ�����u�8��W�3K��t�	�H��r��!���Q�X������u���lչ5m��}ջW/���u�9��a��5X�p�>Ύ;�q$C�����M�4E��ѭ[7$%��k U��{2��3-=[�l�K!�9n۶�))�����C��(�OL�3A��E�ΝѦMk�V���~�:��.�����MIJ�)���+T���6mB�>y��zK�D��f͛��,�u���㐘X��ZT��gVvv���}<p����_�X�����)�T��21g�(��t���k�8t�(���S_om�&���O<�R�>}�]}�������֊����m����ޭ{w�P��螛�J|���f̘����[�nEzz�����u^��t ���x�s�98��S�P%���w���x���٧��U8r%���5l�/��2ڵiS���C�o������
+T�g��>އ�";4h����õ�^�A�����8;U��n�����/�l�2���w/�k����(u�p�)����N>�$�R�ؑ^�/���<iR��r]d��_��*Hz����ᇙ��/�x�b��>>_�͎z�����5�\�s�g[O��J��`��F�ܰdrd�$���q�#T�T�9���u�	�$xUU��\�M���5�'���X�d����Hp�uT�.�6P�]O�ё"��*�W6�{�U�~1#G�ҁ�0��j�L�#�<Rbd�<������ս>Uw�MNNF���zoR����Z�.�1�sp��#�}{���� ���'��o��H׌2*��ґ��,X6�����?��v��#����.�С�)��^��C�`�l�R������;�ޱ�A.ǭ���*�4h�=z�K1�tP���>��U�ɫ3U[����{����z�g����t��.��c�JXd:ܛo�Y�ʮ'� ��%�ϕ�X��$�9[�
y���N��r��z�8�ޭ2�|��~��^v)U�gR�ve�]�b���ٳ����:���q�*w{�6|���0�Ǚ�Zɇ�J�͎��T%���_��u���<�+�ȿ����_�sGvv�_�+�lʾ��5�����y��ǟxݺv-���I�����B��Z�'_�.w�ځi_}�9?��ŗ\��{I����'g�k�|���z9ϕ+W�i���-�����nՏg�T���p�������KGb�*����?�{���K���Uk���̾R�����'[[��>'�dIAa����G��o֙)��L��M�����Z[j�֬^�u��T&��ge�ԯ���(g�pKU0߽[� �=�%~�q�I�������5�گ�GZ����[=�m؀�^{��9N;{$�6%������/�E]�r�Z����5�m��֩��,ǘz� ^U��7����}(���\�;=���}lٲ�����]J������7'��^��=�ܯ��5sm�?5o���ά���:v���)푆V*4u��p����N����|���f�?c�u�!�_L�[�n����|��"�>� /���]ŏ��VJx�n�\��cǢo�^��r&�9�UeXe�sU�-//��<{s][ɠIFsŊ�駟�裏�_����2��-�S�-��⟩��]x��gT@��&��̊ٵ�̮Z��?���H,���>��I����6��x���r�#����D�Х�2���>���:wB��m�Ӗ���[*J>�9*Q{z���믿�^�)��2�J(2���ч�R�J�H<�!C�v'T�%���'�x����d�k����~����@?���B����3�{5j��4dee��2?E�q80��oUf-�Ox�<�$�*�9
o��ffT�|ſ���Gzo�3�up��8���J�/�_R���>������O���$}�+S%57�F���Ƕ-��f�x��r��0��iذ~=�}�\tᅺ�_�SXO���/�£�<Zl�)��m[6]��������۶n�NjA@�����:lM.��t�t�2[�зO�׉�:�\jf���C����໻����m���WJ�Y��d��bX�w��_�h!��^�����_���*ڋ�	Z�1�w����a�B^���t|߁�'U
�4q�Q��-,���1a�J�=U�9�����NJ��= �r]���1��W0��	�ζʼ�������yx�����K/�Nco��^;i(��?��@���u�ȑ#�h�#!����F����9�[f��zH��������|���ū��s��z�
���zg㪫�
�gYڌ�3K�b�c���+�������Ǚ?⥗�cܸ�������eR:����ǝ�Tk��g��Ѝ�bz͹xť��`Ϟ�^����B�.]t5o(]!OR4��Y:t6o� ��ê ^�~��8ӻw4k�u���UT�h��]z���˖��]	��=gö����Ï�k{�E��T�ק�~��%���#"Ѵi3�B]Su���7';�R��Ҕ�n���VS�JЎ||�ɧ8���|�
_/�]	hLl��h��m�"11QG����uo�;v�;�Yg|�T�H��E_�.�W����=u�4LU%9W{y���D�=M�4Vץ�>o�$��RSS�a�l޴I��[_W�2L�:_r�
��0�L0w]���u�4G����u��n2�Jz��]�V]�dx_�X����(��N8�_�������ȑ��v� ���N��B��I��K�.�3�����Qڵ7oެ۶�'|��C�.Fq6=���=�;�^�I�$��t�2L�<����\ރ|O۴i�{�K�HG�C��r�򹦧�y9w��LӁ��}s���c��A>�G���}��/��\=�7mܨ�[�d��%�ף�t�S�֭[6+��)s���2>�����ak2�H!�ک��H 5��_�|9�?5��`�Db���T%�W^y��#פtu���ԗW��M�:����k�Nx�;�oÓO<�F�h�8Ce�Ru tu�+
�R��ۯ/���J�v�ih�����̈;)q�P�9����oM�R�1�f�Ϟ{n֫���]7�
�u0��3p�:N�޽Ѥq#=��s9���6�k\�����}{���#Ìf��:��^��"�>R�s�v.
�a*A�ޣ7�P���[�j�;W���W�dΤcۤI�����e�	�34t�x̘�طgRS���v":�N9�\}�U�qӦMu	�s]dH�֭��ݷ�����W`���"C�O���}zW����3�ǘ����yp'��o�駝����,���!�1�S��߅�����Y�,2K�s�{]VN����y"����}��ΕΠի� g�u&.��b=�q�ƺ7���zA~>RTfm��%�����H�Qِ�o�}�]�pB=����m곸��{p�-7���]���;u������gj��Q#1��u?�Lɐİ��?��kf@�R�+���D6Х�P������*p_Ub'�|*~�a�q�@Ĩ���'9��x��W�������6g�l��X��mX�z%�W	�۪�Ѩa�J't�P�\��T%���;q뭷��JPQ�L�p))�҅<������>V��t�Q%�����[���x��Gq�E��P��8R"�ݳ�w�'��?��*SeyUR��N�m\�а�8T`�*�G��"�*�ȃ�Եi�Jp�+c�\��-[��u-q�
�R��
�e��B�u��l�kޢ�=4LW97�_��K�jת���ҹ���N�ñ��?��IUb���{�͚4���^֬߀ѣ�ww����'�n��s�mh�2c��:��&������Izʿ8�E/�(ٰr�r�S�O|�Mԫ�P�{]�냅�Q������O�Ї���멈s�m�y2��|�q��aʔ)5r�:�����$C�j�9��nE�Bf��Gq��Յ���2����4��>A�I	��zg�'�q��ϬH�Zž�b���u���1}��qc�}˻C<��&g<�[��c�=�i_M��8B�)�|�ɧx���T�V�6j�Q�G��7�Ꜽ���R%����믿�vxz���T��^��K�DwZ�VaoǑ`0d�`]���۱g�.��lܸIWG׫�$.֊�K|ݺ��8����I����[Ǥ$<���X�n}���H&�ƽ8�{��1ͅ-���?U�1c���nƖ�-�c`��d=#�t���a�ĉX��[�թJ��1b�H]����ɞ�V_]O�II��V�	V��3f`�*9ߦ2��Q��J��u�_��T�3�9?o��!�Ho��]Z��~oSKK��|��:��^��X锸��Zzj|j^�9bz.w��멚�)N:rI��+�['P2�HL%&�6�i�ܵ��.2K5�u7p� =L+�]�#z�����J��t5���H{�|�ǨK/��\gW{�C���]����ݯl'��I�ᤷ�*wk�.=��`^ѡ���:^t�:�D�g=6X�z�J�+��;�w�q��ů"ץW������1F�t}��H�[O<�.8�����{��N��T`�>��C�aݺu8EmW���]���-��V�e��O>����+0��g���L{����t�{�+6��hˬ��z(��g֥〥)�|��a�葅����h*�I��K/�K�,յVs�H��c��	�N���Ց]���g��m�vM_d�p/SfVWs~��ŋ�[0�j��숃���V�ǞxLw[�'�([)�l~��ttx�� u��8��tӍ�ڸ��A�L�������mE��ύ7݄s�����9IIpР���O�x���1t�=iK'��֝�RʖL�ۓ�Fj�>x���J\~�e>k,���*�O�4��C("7JG+����S�#S�Ju�Ν�U���|�M�A�n+̋�Ƌ/�Pw}a����$C}��1�����Nt�p�Zb���W^#�j�G�)S�m�U��y�f�?p $k,��Ͱ�۳�&��KG���l[�V��P�i)��~��7�Y��~i�'�T.��SN�|;�����}�}�a���k�������s7�p�n���qM=%�u�]W���:w�&M���`��G'Z�l��.��2:$�~b}��f���A]�&"#�����)�Oj�V�Z�:�y�xm�>C�u�Ǒ���w�5)P����蒤�NS�*	����2��:wŭ�ݪ�D��.���o���f��.�+K��e:��^�\���0��$��a�k׮���B�{��]��Cꚻ:�ѱbJ��M&a.GMkC�_:Qe����B�+�ۄ�y���$\q���L��OI�.��=��?�:�X�b��5hr�9�<����uĀJ�엨J;�u@_�u�SO;�U��� �p��z���L��U-��V�[a���+���ؼE/S|��s��ǣg��*�JB����m�uQ��^�s��Uj+�2�aa�ͼC��z\�ަuk�{޹z� ��ҿ�.�M���[�5h�Hw@�L�kO@�*yw��	�M�n����̬��б�>k��]/�jb�db��[J�6�`�=D���3�:�[�
h��Kz��w�y�c�UU����0�!�^}UB)=g+P"UF�a��^����r�#��.N����72C��- �>=z�@�J���u��$��ye�лO�J��/���KH��uY�C:�z��(���3o�<����^v��F���,u��x�	i�8p &�5�G��ۇ*�"�Kf�c����(�;YAN'���*s��"1tL�v���u9�����M�>f��ܵL�*�W�L�b���:2ɔ���B�F�4i}�7\�c,XY�K�}9���B:]�t��{��_�׶BSO��1 �Ԇ���qb�>/A+�g��IV�mV�5�ef�U������U+Cw2S׿V-�m��zQ_v�ك��Vx}�k�nh߾j�Hr7M<����J&ϑ9�s�n��^r�ש�������"B���VMcNgH��Ւ����yU��n��sTt�ϭ$G*������٧�`)Î��z�Y���j��ڷw���n٪�l.=����� �+KWT��{�ԓ�4k��e�����H:�1u"ݮ]�J��}]t3���A�?�l��%ǩlgTڶ�ː@���;�`0���I����K[7o�|�y�w53+���m�Fe
7O�d�$3lU�.�Ռot4�_˫r����$ш�Yb1��4W�Ȕ���ɬ�i�u}TsV��]R�����<�b�0��;v�eJ��(qq�t'�ʒ�k�')=���y?�u*�픡��&ޛD\%t9Ve�U��쨌M�7##����=\��[Uj�_��d`�e|v�ڭgᓀ~dLDFE�q��Nz%�*ڼ-��b��/�$t���g���3�I�!���*s�I[]%�Ƃ��͝��Y��4C��I�oU�	��!+�Ig$�6:�t����W+N=j��IЊ�=�Z��k\�V2TU-Zer�t��*S)&	�nݢ�}�H&j��=���_�HaS��L�*�Y��?x�S�W�8��A�@L:TD������YCg&~U���JJ2��M�����۷O�U�w��`���4�eɼ޲�CU/BӴi]��(�8��;��[��.�?G��X�(U:�N�H���Q��H�������܇�}޷G��YO�����Ǐ�믿T�o��ѽ��z�����d�1�F��(8I	�^4o�L��]KJ����MWz]=��i�suj);�7�����/�yJ�99e�2�:Oα2w�T�JG��&�;F5J�$�v42 R"=��M��R�&��x#�k2��q6e�&5��؏�d����j�k�#�\m�5�m�Q�ƈ�]���:�i{�w��`&��[�M�*>
U��1���Idsr+7,�nS�+�����]M��W���e<���X�����z�Uѩ��jH	���n����dLm�zu�o���.;�Ɂ������O���V��G��*@Ib���C���l5s��J.�J�*��<�f"W]HG���e��@u�*��d�;Y����r{��jh@o�X퓒�F�3^�kv$Y6P��7o�3e5o��u�`>?��>�P`��+\��U���Q�*��SNUC�1G9��qk%�Nӽ�0���pk���a��򎥚�gϞ�V�;���˗/׳N�`��ʒ�F^}�5|��7�бz��޽{��%�KOfo3_IU��`)�hf��0HR��g=9�!c��5>�'
��L���C�v�\�3G�f3u���@T1�Yn���5��^*�K`?�a=fu��eض-�:f��#%g�/%EO��c�6����l��ZĐ�3z��K/����)�N�p"	��(�H�`)�W5�s����OT͝Oǎs��
M�?��$&�?f��:U0��8ӟznC�u:N�n[`��(�mHNކ�9�]�]��7�B<�*=Ʒmݬ���ڷo�zi����A�p~PzȘ*�gdT}�_��Z+�و���Ы��`^+�{'O�0J�\h�8��TT�Mu�H�ʽRU}'�zY����?���_�e��]	؇���%����t򓕮�ԫ[O�Ѷ��(��Ν;u�۪v�59���v��1̍f63�٤������Y����mT�:1������]޵Ls������U���v���_�d�R8�rF[�nÌ߫�J�̭>RS�v*���� Q�������*K:ffe!.6�J����]�N�L*Svq9������m�2��Uږ����۷��~�]���R����ft���;�-^��k���Æ�;vbʔ/зO�c6C��gb����|�z���#q֠Az-i�O�^�zhּ6m�^�e�Mz�}\_s-������6��u2;�$x�����BNN�I�d�����K.�Z�%yd^�#��n�Ն^3'��%k�r�U)}���^��u��]vN9i�Q�b��yr2>��s���d6�����mZ���O�܇gq����1��_,�"��u�֣e��
[�n�ƍ��mXY�֭u��(ڨ�^�nv�*��|#d	S�z������H���.���R� 'AIa�������������t�m6\~�e��/�q�:��ٰ=y^z�%t萄���G�)�L@1y��X��?�7��s���0{;�������`�1�Х��Qe
N+LtE�i�쟱{��>���٫�^~��ߊ �y���T@�a񬁕+WaŊ�8픓z\��������s�~��*cQ6@�&MФqc�h���:�����N~3u�	[yU�5��]�}�Νqɥ�`��qz&'+�&M������ȣ�e�i�l���{((��L&�hּ��'A��9���[q۱}�f�*���]wމvm����ٻ3�NG>���ckšO�����}'R �=$�����s����>uON�2����.\�_���Ԕ�أ�d/:��]�>�p�'�se6s����巽BL��:/l�
�W]}��6�[��e����+HHH��s"�ë얔m�*�?�̳ػ�[�z"��.��{�*w�R��ۯ�;��f����0u�T64`S�����|K/���ŤI��úw>ё����3�w��S8�����^ݗ�^���k ��r�ÙY���U0���;��2�UI=�S]�h�����z�I�YN�l2����~�m�a�S��p���؟��}N_��o����W�|�^�/��,^���dNt��7�|�.e�:ݎ^��?�|UZ����&m�'N���N9�J�/9�e+V���^Cf�� ({+JO�s�=͛5�B
$��ڧo�4�GX�1�=9/�8mޜ����W|e�Q���o�nW;g�uV��i��ЭÏ4�y�d����Ə:sJ"\݀7� ��*O��+/��6]���O�^<p?ڵi��	D ����3Ĩ��x��`����E�.]�>�Yg���y�υU_��[6���c�L%rmZ�:���j߇^��*�[�V�hѪ.��|]�
���O��UW_�y��!+Ӻs܌�CR�x��'sd�Lxz��^�cǎՙ~o��N���5ADd�^��j1���<�Kܒ%�ωe@p�v�����ª���n�{�X6d��a�oa��ŸM��SZ������6�I]6mقw�yWW��L���NJ�W_}���
�۞eY
��oT���*�;�����J4�0t�0�ya:�kW�DN��c�.<��p|�ŗ��l�$,,�^{-�w��`NU��s��_���V�z~~�|��G������n|���ҫ�ɧ��?{�j�v��|��hP�~���ccbi�?��}���3rM����t�SB7ٖQ��XRU7��0l�CؽSz�Z}A}����O=���'�����y��'�u�V��c^r9��,lܸ�~����5V�Ҭ����X�W<s }����}���~��3>��S��e%��_���}��GqҀ�^�&��Zi..Z�J*���7��/�p��	'���E�������{J��}��WGw��.:s�����q�
�����"G%_��Q����g��Y::{�ٺ�����w����<k�̾t�����z�T��n_���N�e�U�Zn	ݕ蒇L6q�嗫l�	��jއ��Ds~�	���;Z�j�~���G�����84i�1��:�K)\������{�`ٲ�X�d�.�oS9��Y�|��LO��1ϣm����}݄x�Y�իWc��%�J䤏��ٳ�f�\}�5�����!)Ig ��N:mڼ	ӿ��>�[6m.�WYN�l��?��^�`NUi����{���#��]z���eMM����q���~-[�@���}f��`��ǧ�->��l\���8ѵ{<��Cz\zM����j�ɢ֭�z���];q�}`��i�ԩ���9����ߥ�q�1��+�ak�r���6`�ZD����_�uz���F`�~�+odC��v�����٧vĨĠN|��)�H@�ǲT@Vw�����}�߳|�I'�ŗơO�^���ӫWO�5��s�^��[-Į�;0�����T/5+��e<�L#����g��)Y�p!�'o��᫆����`��0���@T��b-*(�y�ر};�y�/C@��z���xRe�'O���w��4j�	ut'���=m�r����زe�*I�.��{�F���SO���WMIg�}Ʃz+U��s�^�ru2���4���as��2q�i������G��T@/�#�蚢*\����$��z��c\r�˗-��Jg�[��d!�Çӽl��J���0���{�y1�Yt��9 7�9C�F���裏b��M�ԥ��k�v��~�=�UxD�c����<��Ư��M�5�SÇ��T����hеR*0H&2?� ���C�v�m�#遽i�z���˯��uהφ������3#��y�&x��q�X���d������u2
���X|�\������{�a���HP����z�Q^���ß�Rsx��e�^�6mZc��Q�q��ɖ��\+o�:W�L�ÿ��[q��w�I�FKdH��a�����ß��E���^)z����I���ʕ[�ҵ�J܆�63���&%ntlɽ�X}wF??J��ߞ�6�I/k�Mi�W��*�+�[^F���mݦ-�����
�\�����G��X����f
�))ػo��Ŧj�
��k����={b�ĉ��������H�|=�ze��W��SO;��s7�W���$��;g�^Fv�8���-2����U�9�s��:�	���K����ݺu�Čp�3���^��:�=��Ӻ���W^����aZ� X�E�ʻ���=22��q�}�����DU�]N_�#�=���{?v�H��A����HNN>f+\)���ˣ�����?��ުґCf�[�j5������G���!O�[OO[y�5W��s��OH�۽kL��:��x������,l.�H�M���O���O9�]w�^�F&�����^!N����5Z��W�������@�S�Z4���q��^��z�Ksp�	�>����*�e���G~y]lt4n��z=c�dοV���7��~?3��C���
�Q1�ر��Tw���6jРR���Ɏ�{��^�Z���bu<��qD��Is�|��F��}\(oi���9nӦ��=Opv�A�Н�����Ti����õ�K�L���m.���lݲUw�������HH�G�vmq�	'b��A�ӻ7��M�[�*Ty_҃]ޓ�������3�`�?ر}������К�fG�
�mU�\f�2dN:i �={+}��^�[�e�v:�zᜰ��Wmʾ���t�ֽ�LWr��I�V�!5r���֭[�kWu���Ǒ��S�Jur��=�d�%�v��!`��ʔ��{�,�w9���� ̋.׿Es�믎Ӷm�A�Hy�:��2r�sz����9?��ʕ+�����ɽe\
Oa���Eb�D����w.NS%r����Vi�٣�
n9% ��e��/=���tb릮yZڡ��/Sjk���W�\i^�fK��|���i�Oزy3���c��B��Zj3dTP||�����K����]],�J���մNG�s��gC�t�8�3t�;v"y{�^&TƖ������Y���HH�ڵ�PO���5k�\y�W]�fw���[�9��&w���ur�v�Y�F�N�e��Y%#=]�Ws�$*�j��^f��ر:w�W��#d����׫�	Z2���$�뮻���V"""W��+�I���>����QQQ~�ŕ��qϊ]�#>@���S�/�r�p��}e�#������-7�d��|b��+}lԵ�N����6m�ڵk�z��}�����lnn���bս.�=˒��ڵC'��v�{�Z�Z�
��s;��S��w�-kO�\�����S�|��/-�%� _��C�:�����Sqݮ

�����~%'�:u�ѨQC4i�T��1�2�S�
Ԭr�"�W݌�*ˣg����ِ\���5���@$��A)J%J2�Qj�����_��%�o��>�]� C��2w�zߒ ��� ��Ë����}�u�Dӓp�:�ʪ���qU{�o�VD�=��������"�LU}��qq�Q��)�/�I���&=ⳳ���ס�}��$�(:yHf˰�O�H/����r�;P�7��aUu<O�Tc��Q�9��k������΀^)f�K)C�\����b?�w,��#��L�im/��;�hݥ��8��|��8ގ)�ňp�z�����<��58��0K���0�~L��6�@;�\{u�yy�PM����Ni��f7����YB'""
f�S\�[y:�Q�ѝ8�)������^����3�-ӯ6�|v�#""
b���������(�ٝN��ֈ���7=S\�[�,HN�Љ������W~	]�9:����T:v���3M�r'"":�����,�Tn�7+�O"""
�K�ݯ8-%tFt""��d��m�::QPR1����DDDAKW��UBg�8""��e��˝Et""��U�:#:QP���U��8t""�`&U�~lU�?"""
F��ΈNDD�̊��3�)݆ι܉���;��~e/w""�����,�NDD�L��YB'""
jXm�m�DDD��"���������r�z�DDD՞S�r�5""����U*�}�k�r'""
ZR���VN�f,'""
fz�5?7eX'""
V�ߋ�0�'��,�U{�˧2�5?�r�܉�����m�r'""
b��U��DDDA��Nq�����(��~W�Q�b�;Q�Ǚ∈�B g�#""
~�C�˧2�+��^��DDDA���2DDD�ʏ�\�L��NDD���ΨNDD�����*w""���*w""�`�ʝ��(p�8""����kb=S+'�܉��B ;�U\m������K�p.w""�����\�DDD���X�U�DDDA��Q��LqDDD!����,DDD�*�˝m�DDDA�ɉe�������CgX'""
R�
T�Q�͉e���B��m�&�܉������6t"""
F�U��Gk��DDD����܉����
t�#""�`���WЉ����Dh�m��(񃈈���aT$��UBw8�HKK�!�p���� �`PS
Q���c�=�l����j���둓��ז�n��0l�C��Wæ�5�������]8
�������p����*�&6���e��-�8\yS~U��^�t1����h2�g�.��6��sDDDt�I��f4��&��� ""��JJ�:�烈���+UB7��͖n:�� ""��Hfsأ��ege�U;6�-3:::�^�n��������{�g��0=""�I&������K���;w$�Өqӻ<�t^^^/�4cTD��u�ƪ�3*8���c:1ϑ��g�#|���g��OF��x���$�����jժ�y�����W�<l��k�ŧ�O����;v����LP�F��]mn�G���E��l6�&m�v��0�æ�`ap�4�����rd��ϫXf��Ta���
�+����ſ�F�_JoWl����l�	�Q�k1׉x����󇢿B�8*�g�J����b{/���}����(:f��Qxn(���.u��{�`[�~���0T�.b�ҥ�{v�
/���G���NC�&M�T�^n7TWr�֬Y����[f�������=��ILl�o�Nɟ�f��MX�<[Q��}y�~����1�\4%�Y�wϮ�����,�{������vW��3K���yxv�c?%�l�Kb�R��\��W���)|q9��,q%��[����ĮK��}���n�a���{��_�]�r)�'�z_/)���N�l�b+��(�-6-�Y�b����J�-��ڨ�9��G�}{ΧԖ����t��pJ�e���%���-:�b�G�J�JM����.rџ�ݠ��:IϹ��\�������0̘�hg|BvIIs�����Saw���ʇ���G4�΅�Ϡ ?W?j"�gY"P������Ӑ@�p��ÐB�l�S�t8W pr�����T$u:�Õ��p?����w���&���\]$�b��$�o�^ܙ���kѾ����m6�����u�]o�ٽ�ً\t�Ÿ��[Bnn�;z��͸�λt"Q���N���on���'�<�������OOL�<O�EyUw�g��&�%�f�L������õ�Y�I�?\���u����hY<u���	S�,�;u):/��s�]6
ӛb�r�����
_��G���R�����̰�^����kc��4�ͦs�6Wy��-5�0�\�����6�]^cs[�e�._�CA��o��0RB�zHٿo��>�S?�� O�l٪UH��7�

���Vtx�is8t��4��J4�m�j��m�w��/�(5�_�O!_ega2�J%J��#��X�]<�g�إ{�i�'6�^�٧�Lexb�Y��Z�;�'���|��������Jl��2y�.�-�܌Ȉ��Zu#WD ��x���\���j�ژ��~̯s~Y߿}���E���[_a��p�2�mW|�ҥ�R��(�P�F�s+��(��/��(]�*��2�M��x�k�9��?ós�t�<�t�B�{��#�?=�Og^�{Tx6�k��F��'�����ܙ��r����w��=��M\�C���x�y0e[��|�}������vU��2��pU"R��Ɂ�
��c8�Զ��r���گ�S������r�Jt�ܹ�ug����e�,���o��� ����W;����"�#

�eF���e���سgZ6o�/S�T婌���o�c��-]:�mҬ�ks�u���'`��u���+AD,Щ���T<�$$$����J��ʬWr[�l���kt@�`.�;���*CS���f�^��?�>��t��6��{�Q0a@�2ڷh�ǞxR�����v��V&����a�?�`��A�>������_<��sػG��R���Jn߱ø���vh�] "
F�d�q�&�ݧw�_|�^�ڵ����������:��m;����x�駱j�
������f͚���/s�~y��6�w�� "
6�d)-��p|n���V���]*�J[�j5�nۊݺ�:ҝ���1f��y�l�i80ԫW��O>��/��Lꐄ�cǂ�(1���N�#:&f�
�y*�G��¦;�-Y��������λ����(�	N����h׾ݘO?�$%'�0���:Y�6�6m�ʔ���#���5*�M^n6����\s"��Q����{���K���@��0�=�Q��o��}�'�?�fM��;�"�`ŀN�.��b\{��6�#""|Wf��Ȫ/���K����^�jӎ.�bي�1b$��މ��\�����g��w�;��>�Y'>�G<"�`ƀN^����۴9�����U��Uv[�n����t@�$������ѣ�d�b�	�JtTTr��-�L�655/;DD�:y����`r�ڴi�Ff�*;ͫ��b�e8���Q���㭉1��o`5���W��k�.���� �n��O?"�`ǀN^}�~.����j���s�yyQ��q8�p�"���"*22��g��oLx��ٰ*�׊��ѭG��Np�����޻o���:`@'��M�ݺ�@TT�&e~^nS�v�U+Wb_J
Z4k�`�i75r����`��y���ϛ�����C��޻Љ��`@'��z�\vŕ��Ď�QQ۳27-���m۶bÆ�A�u��~w��b�vs�ݞݰA��+W,[8��G�Գ;n��jU��S߾}p�ק�<{�Z〭�%�:tK�.����`$����˒�����|�)�ߓ���mxi� "�N�ɧ����
���e�Ͷ��뻗�t`ѢE��ɑ�AՎ.'+��'�h7���]ٮ}����-c��� "���ɧ_�͚�D�:�W���g��^�j;iG߻oZ�h�`�״����p���n7���hܴ�����)_}��K�aԨ "�n�ɧ��.B�=l˚ի����Xt��۱~���	��SRS1z��^Ǜ6�,����\�պ�k0�|���K "��Щ\	uиq�ݪ�%=-�M�-����y��y�5�fϓv�I����v��:uz��/�ʱ���)�����b@�ru��I��9�U�a�Q�c�t`������Flt�1oG�v�7&L���[��#���7o�r�/?��y���ؽsN?�tUW�T.w�8�{�^�򚣠� �j�U+Wa�޽hӪ��x�#Gc��vsy6���s�͜�����O��3O���:c@�r͚5]��@|B����������e���ؾ�֭?f��<�`�E���_{�����/���w'OQuǀN�:��q�7�t:��/]�+++�n٭����v��:��(���y�EtL̎�mڌ�����0 ��Qv;"����_�z����/��?x�`�mLӡ�S���BlL�QoG�����7����`n���7i������3#����`ND!���Ҹi�rӍ��:���l��]y�e���ػwڴnu��MB�Ju\�j߻w,�����P��'�<��AC�1۶m��oL Q�`@'�<��Ø��iG_�J�9y+�Ihݹs'�o�p��������`���n��]�v�g�������q��_3�QHa@'�HǸ�I���Y����J,�v�e˖��AgU�9I0�/(��＋iS�I�?����#�7i����[2���ѳ[Q#��ÀN~��q=��t"۵�߅�2�3,�V3��ѳ��sƣ�4�g���k��΄U����s/�`J��]�v�Z<x߽ "
5���m����n94��S��`5��X�z��KA�U3�g��u6�y�w��˪vUX��]��Ν;��釙Y���� "
E����Cҹ�ٳW��av�� ?�2��x�M7VY@��JO�ر�������n�ڢeˑsf��)�a��_����Q(b@'�=8t(>��+ԩS{UDDxFA~^�	f��Ұt�2�y��*9��~�?|���0M'���e6���Mz��W�r�x���0⹧AD���o���Z�i���M��ѻ�23�Xm�׽*�G����ܹxy����̀uU���s���Mxz�3�5�[��ND!���ֿ�?^Ƥ����/������m�5�Wc_J
Z6o��K0߲u+F��m[7���m�ڷ����{�r���_���?Q(c@�
9����1))�s�n+m6���Hޖ�M�6,�K0����K/��彩�-�����4m�t��?��9���дi\q� "
u�T!��ɨ];			K#""rsrr"�n�jG_�l�vj@��0M|��g���>���U��a��~�ĩ���K/3���1�Y��Q���N2��3q�"22r}dT�����&V������%K�������J������k>^�"2��[���ۻ��*�<��?�����n4$kBGMk׭�bv�r�s'k7��f�v�Y�j^Rlk�Uh3#l[��dE!0�&"��*'8��e7��s�[�<|?3g8����w��9���L����ܶ�3� ���~�>*J���k������%��8m�F�Y�Dz򃴘מ���5k��\���G�|}[Ǎ�� ���T�|~�3y��' ���~�6�f��ҥm�3�t��_`�Kjj���ٳ
����Z:;e}F��������zWxDĎ�~����
� ?_�n� �pB��oK�zJ[`ƞp�m%��e����A�%-�-RRR"���;�jQ��y_v��]v�����	:���cGW@@���1��v:��Ç%.>ABCCK||}�m6k�����V)*:!]6�x�}:��W���Xa��MY+��f�����	�����Z�N��M*{��:�m������gŠ7T;v��J{{���_�|%M�&�w����74HRR��*+�^Q���ᆌ=|��W^����አc@�B�d��Sr?ʭ���0�Ӹ��*����	z_h1���ƍ�$���<��
�?w�?����/�k� W29�$��ϲ.%��*�~���p3J�su^ZZ*�Ϝ��s�ݷW�l�"6�U<͛�Un���o�ަ��RXX(��� �pE�1 ?��DG��M�'����X-���q6[�?^$֧�b4��禥�Dq�$'�H���t�����=>�Ճ���; �.\���x�ጠc@���f�~��������k�X:�=]Mk����-�q];��,)�k�d�	����N'QQQ{�WO�?c��v����+ �;��������L1u�
�k/{�$?w��������&[�n�?�#�}��Z!�!E3�e���hjn�m��  A� ����c�>bޙ�uZ���{ڨ���(��e2c�t���ҝ��'37HW�7ڢ�r�K�Z~:yrʮ���t�3R[^..  A� DDE�,0��_�Sl��~�����(/���EEb�Q����{W���%yM����Iϭv7��Fo׍��;�צ~x�;��Ȋ�� �_6w�,���Hxxx�ȑ#-�W�~�o�����XZ��亠����F6��Jj�:���/�Ӽ���ZdT�;�ߙ�>����%9�� �w:L�"uz\����-��dn�����R[S��o����)ٻ����i��%A����3��^{�g5���*� �C�1`�G����>Ѿ^��Ω����t��_� {��S�Iz}O���]��.�X����s����s�bc7�d��ߕ�P�1���y� ��:eF|��
h	)3��6���8m]��۷K��Y2g�,�8wN��$u_�WK/��i���_�Т7W�|�.�,~H  �"���ks��y��t����ߔNj��%=-]���$c}�=rD<=��]�GFF��=gv�ƍ�N����
 �cP^߲E��#gΜ)�;엺�����򤪲J*����Ԗ�u?o8j��֙�fnX���g�!�>yR  �t��%�n�Nʻ�|\z��t~�)�'��MR�e���i�L�]���훶lq���ɯ�<)  �:�d2ɒ����������ں��tz�~���w'L�X}Ͻ��ݺu���ݻD�d;A��tZ��J�:m��/>q����ā��%�GZܽ s�����j��u�̝@t�'��˧G���;�x�iʦ���X�V����`0J\|\ުU�v,8䊈���� �aC��?��{\Ǝ���?���b}�.�K��`4��W�Ǜ��j����pF�1$��^��:f츎�G������q���>��K:�n[xT��i�ؤ���[� �Cf�Ν��ޮm�r�������T����C�i�+��<�����-�  ����2˖,��/���s�J�ط���w���-���*<!!��]wߕ|������� }G�1���ِ������l�X��m�I=��������3>m�^9��ŕ���*/���  ���cH͙3Gv��-oeeɁ��"_�$�ݑ�]�Qn���z�;f�y��g�9��ӈ9 Aǐ[�x��d2���D����t:&8�UN���|�����`4�1��Eǋ���ʤ��V  C��8UZ*:�QBCB�'LL375�X::��lA:�����'wtp��u��wZ,�z�j1M�$ ��!���86ih��^��������dn�:V: `�:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
�O��Ր���    IEND�B`�PK
     ��d[��EM  M  /   images/d3694a2e-5bba-40c3-8069-8db85c4c9209.png�PNG

   IHDR   d   d   p�T  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  cIDATx��]	xLW~��d�(%�J"��}�%(�Z���B��_[y~R�R[u�E[[����J����ҿZ��j��B)��'s��;��Ĉ����>���=��s�s��-�37:�PTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��AW÷&��z\I���7�)I*�Ev�Z�:d;iJ�3mtRɲ�������V�$IY6��"a[�d��$}/����~�l���99��t.��$u0Z��d�M��(��5D��a�}0�*�
��?���h��dY~�`ȫq+��L��yY���@���[���������ƍ����0��`�Aк�C��"�|<B&�������r����t�PQ:�;w'N�{˧����a)y���3�t>���ʂ
E@fB\yyP� �f�3b�1�(p�3!�<ÃY=��䫄(�d���?0��&1A3vH�JIi�	�YCd��c,�p?��0���g�Ж���lqtws���%b�G��ɒ�2d'jaxR�v�Zl߈s��S�����_C���2Js;�i���8�f�ɒM>�Q.]�����С�x�g/�5J<����зO̚=�g����f6.:6lX�t]������B��5�D��;ѽ[7���s�p�0g�,�n�=_x��(���E��~/���u{���F�m�6�2�h��!����v����;����dX�i5�7�}�����ٿ�2~޳?��#n������1p�@xV�$��u˖�Ѳe��H�zi��|��u��,�Ν'�����ԩ3�/�5PP��7o���,�_���C�޽ѵK���ǚ5k�t�:>�,^|q 4�XȺ����7!&&�+{�_�~��d��ǎ	SԥkW�o؀������A��n��B�p2�7n����Na��>$3��ARLN�G��&����~�� �����QQ��wq�������Тe+xU�ºu_ lQ������͐�լ�K�.����ԙK�.��9����(�QN4|���X�p&M|�����5�OLLDu��x�"�.Y�9o��&�l7ww7�b�rD�c�)��?��޽E��jO����[���a�0�?B��ۿr6n����o�Y�}��E�E�:uh@lAZZ*�i`5]�ر�u�9Ǻ��<s�4�V���ի۽��1�Q�n�:AƢ����D�?O�F�g:b����a� i4puuÑ�#������W��u� ̜�iL8^<H�Ȏ��ʕ+Bui������®�v�u�zS����u>l�ФΝ�P�U�@.��+��������^M�5c�L�L��S��nW",�Y��e��'""#�|���'B�B�FMТœ8���	�R��ӓC��w��t�b�_G�R׿ƛG߭~=L�6U��?���קў��ݻ[��Z���\�rLd0�q�	��o@Ey.D<kI��
2^U��~�zB�!C^65V�E�6m�W���$!-^�j� ��溃��������͂�٤������m׮j׮����{��l"��e����G�fg�AQ�%{ΫbM�6��F�흚6m"�.\@�ƍD���]P��	��g�ΕG���e?h�V��\��ӊ�����ٳq"m���`1i.�[8c:fd��Y����<P��6���׻�2�sq�{dDG2kd'j	h�͛��)2;U�jW��%�=z|j���)�b~b����!JcӁ�L��+$3�i��ߪ[�Fc�8����2�F����~~���dG��?��%\�9���ɡ���3lw[wGDD���Ç�6�V�Z8AQ?��6U_"���YԢq�0��$��_M�i������W[P��@�nns+�F*Z��@'����!����ǤI��`�<a�CI�>��p������<*T�[�Cɩ�1K�,>�>}�/�h�M�vhD�*��89�-�aq�֭�M0m�t�jQt������5k?C��M�ۻ�Mk5���Z�e����ZSVY'�����L���������'����F����g(4�Ŷ��P�^G�>|<(��p������_�R�VUDK</`9rr��WhI�6��E^��9��~��΁�ʧ(��K�c��K�^���}Ѭis<���b�s���J�efp �e
���,���5��<�5o۶oD��h���%.�sab��F��%a�ȑ4I܍��u�Ȗ-�!00�==̤?�9@���������A��"���K�T����J��2
�������r�̋h���C�Шn+���\�t	�i~`�'t�dA�����Ӄ|�'���GEDCQ��z�5{zP�gA`�@��?�h����\�h*��5���]�r^^^pbb(��1��[ޒbo�ػ^8�s4�叽|�4�@����4}�#0(h�my
?A�#����Mg�<��7��?�il���_ �2Eto�����"����j�37-N^��4g��)�8����&��'�*JBCLQ�JH�C���=d��,���}X5D�2`�����0��g窆(&Q#,���!�.o���e�TF��[���9ʲIQ�[�<l�M�V��|/="D�xOR���vG�_G�3˚��7��aj�gE��s�6��ˋk�Q'I����܊�GBEiB���j���QCG�h4Z�D�$ݢY�-R��By%�V+i�T���I|3����4����ĉؙ}���2r����)���Om�fk\]�zH�|�R�iO�l�Mۗ�I6_dْϜf4G��Fk-匷�ݥe�k�\𛍶���V���_�3���X:�-�b(ڴ#ݾ���KĤ����h$�v!VI~}��+s�^����xg��p�h4"�E@�Ӈ$^N������1���	�����ǁ=j��������o��qbZW�?��i�1��wI�t�G��v��e��^3�x޹���k+�t�w��`-;q<3��rJ�r�##���Κr$55G��޶;�a�±c_�ٿΜ�V�{J9�Ԕd��=�(B���}�\�.1�7����׭w�^v�.\�[��"{x<����̣������{�"o���]�|ҵ�"#��[v��n�ٻoޚ>�Mۢ�̛;[�A���(Ks�#�����@�V�s��I������׸��������gn�fV��8\��@�*e	%F��#�n�����8v� �2�Ǎƙ3�2+yV{<6���ܜ����#d9�¡��ȏ ""�z�ז-_�M���^nzjJ�QNk��i�܇��#��~_�Z(_��?���&��2�G9��ɡ�=�gge|�yx�fY$�Q�/R~�'������ll���<����� ~�N�z�����t
s�PVQ��<^�q�s��mOrrJ@�=�t-���K		粲24x6�;�;�%JHJJ
*�|D��-KKMN!p5�olI�x��ݺ�Ge�F��kǏ�H�"A�ռ!i\�xzz�/_�<�R�u�7�u�����U�F��K0��N�rx����̬L�(B���^b���x:y9��}���E������k��%u����QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB����Blg���    IEND�B`�PK
     ��d[ZR�y�Z �Z /   images/f51f6ed9-d8f0-454d-af8a-e11415a94f15.png�PNG

   IHDR  �  '   js1   	pHYs  P�  P���Dm   tEXtSoftware www.inkscape.org��<  ��IDATx���U��Ϧ��酄H� AJDz��D�P�@T���J�RB	%�^ ����Fz��o��ܝ̼u�}gv��y&��}wf�̝;�ι��ټy�(��(��(��(�R^�H©���m�lg��f��l��Vo���lx*DQEQEQEQ����l̶�l+�����6��͛7ϗ��8�n9��`�fke��[��EQEQEQE)��f[h��r�u��>3��f{����<�Dtsa�0_.0[_�u2[{Q�<�ٳ�t��1��̞=[f͚˾[�n-�{��:u�},/^,ӦM�6D�����K߾}�Y�f'�W���ӧ����#߷���ԡC���?�\���X���@;�f��޽شiS��nԨ��L4m�T�d�ʕ^������M�ӧ��m�V���>�/��2�}w��Y�w�.q��W_Ɍ3$��wM�4���*N�c׬Y��k׮��E��<s�Ϗ'�ԭ[7�ڵ���ܹs��O?�e�-Z���'�{q�t�R�?�[�.�}׭[��O-[��8Y�~�7�b�A�=�S�N7qڀmڴ�^�z�n.Z�Ȼq؀)���:n�`w�k�9��=�|}�l7��Q<7=e��=̗�e���%[�䊒7����V�Z�ntA�.]�^�z��2J0���Eq�k׮�aÆ�|�4����~�g)�mòe�"�'bj���Ҹq㒴����������{�=q�3����GE*ҹ��c�Ҹ����;�,���'֣��?x�`π/Eb,�U��gDF	�!�37�v�A>��HE:�{��������.2v�Xϙ�s�5�U�m�Y��?^�͛�q� �4h q�c��L�4)���8�i����#�v�g������w�СCe�ƍ��'Λ���F.�q0 nK1�22�O�:5��b��޽�i'qـ����nh�c̘����f��G�3:��DI1�a���l;�Fʕ"� ��Q�E�J�[q�aG2D/�hw�-��R`���D��D��̇����D:��S
qn�}8*�n�9�oQ� ��)*�n�y�v�"u"e;���G%�1H��~��r�a�J�[q�����}�cF%ҭ8��d�)��A�y��J���DPő]}��V��*U�w����Ü;��(U�ƉZ�ӗ�S����n;�kT"ݵ� j���~�~=ӌ����W���8Z2�n���r��v�-���(�8/Q�tw`.5QЮ8/5Q�tW����Dz9Ĺ%*���R�Hw�y9�J�[q^��8/5Q�tW���(E��� *���R�Hw�y��R�[q^�����Ap�zm��7c������caL�dt�l�<�E��r�sK�"���������R�H/�8�+��)�-Ŋ�r�sK�"����R�H/�8�+��)�-Ŋ�r�sK"����R�H/�8�+��)�-Q��r�sK�"�:؀5�n[�������z�S"Mϊm�1'̾j�S��C%"� �-���$̖B�$�sK�"=)��R�HO�8�*ғ �-��t�g�C�Ź�P��qn)T�'A�[
�I�bDzĹ�P��qn)T�'A�[��I�BEzu���9��#�5c��Q�8��Ɯ�`��f�AD�ֺ��$�-���$̖|�$�sK�"=i�ܒ�HO�8��+ғ$�-�����sK�"=I�ܒ�H��?�.	�ܒ�HO�8�"ғ$�-���$�s����\�t$I�[
�I�|Ezu��*p#���3Fo���m��6��~l���l]DQ"$�����%� �āْ� �Dqn�U�'U�[r�I�\E:���RE���HO�8��*ғ(�-���$�sK�"=��ܒ�HO�8��*ғ(�-��m�$ғ(�-���=�M�'��U�WP	���F��]3N�jƕw��Yd#�9���Ͷ���]�V�q$y`�d��<0[��I�l"=��܂H�p�9sf��,�-�Dz�Ź%�H�yf�y)�9/�l"=��ܒM�'Y�[���$�sK."=��ܒM�'Y�[���$�s���D�ڀ�AEz$M��'�0�ʯ
�I$��9�6��3fۙoEQ"$�%l�N��l	�� �-a"=-��b\�HO�8����4�sK�HO�8����4�sK�HO�8����4�s��<���ϯ�4�sK�HO�8����4�sK&��6`iQ�	,��8��|%��w�ܢGs���˿�6X%b�40[�t�f��N�8��Ez�Ĺ�/��$�-~��&qn����s�_��I�[�"=M����i��b��\)��$�-~��&qn��4�sK�HW�<�H�����֌��3c˚|������5ͩX�W%b�80[� �hѢ��h�����{mH�8�X�N�.]��N�[���!�6qn�F
F�$M��bE:��gϞ��+�#i�+�q\џ�$�-V�ӟxߥI�[\���-m��bE�ܹs�q*M��bE:��D�Ĺ�錯j����� ��׌���wn���<��3_5[oQ��I�8�0@ӆ4�)K���e��vK��ł��ђ�� ��4��>bĈT�'D����%������o"��|in"=����w���Hǉ��{�H�u�]=��V8w�aE�ǧ�`�@"}Æ��^f{��r]/� �n������\�	��N;�/ɐfc�R�ThJ��>T�3���3Q]��"���R��Sb P��'��k���4ۓ[#��}8o�nvL���6PEQEQEQE	�+�=([�g$/�n�9;��ن��(��(��(��(�@wf����7o�2�����*���T�#�����ߺ����(��(��(�R,��/5����G+�u)��|��r��l����鯅}(g�nvt�l	�דҀ�c�/�6�lo��}�-1!X<��ٚ�qNT7��4��:���(��(��(��(���\�})[����e�f[a�U�E�#�ъ����l;���lY���l)�Vj:��OF[�4"}I�r�f�%C�����q.�Gf����f�H��m�ƛ��s�̑?_�܌^���(��(��(��(�Q>M�+���Y>����̧f{����Dt�(��b6V&#�[ʪ~�w�R��2����Z�x9&�'�ùT�ˆ����s�5_.�-Q���JBi\S��o6۪�ɮ�Z��&���׷z]�lڜ�ʡ�?���z3�ې�{�����?��4q��$�A�A�MR;�)�^W��'I,uko�zu2�����?%���eN�a���D�S�z�M[2ߋU�?mNt�d�S�Ϭ]_!6%�?�L�lgb�c�nHvjd��lE��ޟ꛱�N��'��������m��iG��6��uje�I���s��i�ˌƛ]���>��S��A�[��W��l��R�����g�s���Y��ÃdKi�8`Q�O�v�9��tn����˦-��כ�6T��<(5�����3h���^�����J�6�2~���[ɬE����?�;��.���Of7�'6���Ȉ�l�i�y���Z�����D:�X��3��Z�-K´�`v�JF�Y��3�|�Dޚ�D�J�F䔑3~f��:���6�d��P�7��_��me���.�{�e�v_g�̫��ʇ�7��ҡ�:9f�⌟�bq=���V�dN��$����v�~crE�>��ˀN�3~��OZ��$��h�V�4�g�}�@���Y�9؀�~����d�Tz�ͼ������k sV���Eq`k��eF'^m��\�L��.�������J2
t�Xe�6[�8�HI��9�R�q�5m�S�D�d�>�(��(��(��$�Q�;��q�8�9޴+�Vd�5����"M��6����0[�Z���Dp�r�O1�)1��vs��و�W+W��(��(��(J
a��Cf��ȶMRb�1)<��/2_/�-�����c����P�n>H��{��Rl���َ1'�Jʈ9�\�ƽ��d�cE�iSEQEQE)3���8�>�9�[�V|I�s㡘[q�l��I|��hÑ6���N.�7$�����6�����EQEQEQ�����	LI��`��c��7��a0,�C5��o�7�o�� )�Dϣ���rh���%	Ĝ�զ�Lο�l-EQEQEQE)��v��dS$a��U�St|��C���v8߄E�)��?��~�lgK�1�&s�8�-��~EQEQEQ���vbŹŜ�R�1�}�l��t�]�1��c}&Џ��枿c��gK4�/5��li�\DPQEQEQ%���%IJkck�����1�v1���.3�ۈps`����@����R-�'˖��vEQEQEQ%jȲ��щ���`�u���t#=��#��+��䗚�MXn����̖a�w��.ߗ-ޑN�(��(��(��D�f�����d��A濣b�}/���"�Q�e]�(x�4��B�y�3��y�g���+��(��(��Dk��8eY�.>g.zTY疦f��?�>�l�#������ӏ��
(%�O�k��3��ż�Y�0gc��,XU��x�bq���b��d�a����mذ)�E0��M�A���i�ڒd�ϯo�1�^�u]I2+���ڟ�mL�}�W�4�:�2���j]����_6��K3�?�Wԓ$�xUݬ�i������'4�Z��mL�8���������e���-���?�X���Tl���5�If��Ăɶ�^6�|��s��+**�f��s��n�e{�O�h���0'>KR�9�U��?*[.|�� JV(Q8����v�,I�a��V�6[����Mբ?}�(��i��u�-ͬ�P�Z��Oԗ��`E]oK3��U��i���v��=oY����5f|Z���Tml���go�@�%�~��~��E��NA�b��lWH��" ǚm�(��(��(��(��4�9�rL�WTT�C���(�HZU
ts v�-��~���ek���D��(��(��(J1,6۵R}�I�� �+ʝ�t��\��֚�n�^�,[�Eo+��(��(��(J!Lۼy�x�&��|]QQ1Ib軛�q��c��'�a.�tsᧉ
tEQEQEQ�ByQ�w�m�EV8��;G��OS\.?xzvEQEQEQ%_Ho��T?^0�l�p�5W���`�K��!��d�F���e˖I�V�D)?�7o�F�����%9hR%����D�ڵke͚5Q��K�?�J5ôi�y�b�Ū�%f��TO�2�<���$|��G2dȐT��E�ɒ%K�w�Ȟג�n�:�2e�0@��I�RVS�N��;J�fQ�"Y���+Y�z�t��]�
/�3fx��V�t�^��;q�D�>4n\쬰�1g���\���+WʬY�d��O� ٸq�ןxO4l��e����vQ�z���y��I߾}S۟6l� �&M�~��I�z�]���D˖-�,3؀���'�#����x�;���w���R�͐j�V�i*�KFK�E:3�i�&Ϡ�ӧ���c���_�	áC��R�c�̞=[���K6lX*E:���O>���Q�#��O�%^�<�i�\��?�X�ϟ/.��w�9�"q�s��S�N�6������{�v�!u�ʾ�/^,K�.��SE�̙3eڴi��<xp*E:���>�.�'b���Nhˊ+���F�N_�Oծ][m�2�ڀ2W�/c�vvT;s��b��Ŭ'՗Ţ����tw`^4���?0[�%M"�F:��'�64o�\҂_�c�@�D�+��>#i�8���M�[qn���I���xF M"��`����t+��>#i�8�H�Hw�9���)M"݊sP�|�$��]���o��R|��ó�� ��[��}-���2QJN�h��lI� 60�I��Ź�1i�~qnI�H��sK�D�_�[�BfF�&M$���9�g� ���ܒ&��疴�tW�[�&���ܒ&��疴�tW�[�,=1�s�j��Z �K���T�F�!�	
	���/��e��-i���i�a�ܒ�&�-i�a�ܒ�&�-v�^�Ez�8��E���sKDz�8��E��sKZDz�8��A���sKZDz�8��X:b�@��R}Yi��V2�6VE��uR�Y"J�H� �m`�$y��u`N�H�&�-I��Ĺ%�"=�8�$Y��<s�Ĺ%�"=�8�$]�g�$��l�ܒt��I�[�.ҳ�sK�Ez6qnI�H�$�-j�O���;�l��3�m4cDdZ�Z׈�dYF�c�(e%�t��%����I鹊sKREz��ܒD���8�$Q��*�-I鹈sKREz��ܒD���8�$U��"�-I鹊sKE����|yn�K�*�s����TG�A��u}�޴��$m��w`�$i���#80rlѵ�u�M�)�|Ź%i"=_qnI�H�W�[�$��疤��|Ĺ%i"=_qnI�H�W�[�&��疤��|Ź%I"=_qnI�H�G�[����s@'���f\�p����R���B�����Ѕ̖$Ѕ�s���酊sKRDz��܂������C�E��ܒ�^�8�$E�"�-�̈́	�kѥK),ŵ�W�[� �疤��BĹ%)"���>��üŹ%	"�PqnI�H/D�[����sh [j�UWx�G�����?�Kuo_�(� ]��la��x�۷���bŹ��"�Xqn)�H/V�[�O��}-�HG�ӟ
�r��bŹ��"�q�b�J/�H/V�[�)ҋ�r��bĹ��"�Xqn)�H/V�[�-ҋ��dB9Dz��9` 2ۛR=�&: ��-�`U���^�\�
� ]ʗLT�e֬Y��R���Ĺ��"*qnqEz)��Ĺ�"=*qnqEz��yF@,X� ���"��D%�-V��o�^JET����R�8��"��D!�-�Ho�,���r"*qnqEz��J�[\�^J���b�#PSqn���)���"<�
t��2�d�f�x��м(K��E����l�"�gϞ7\�(ŹŊ�Ry���+����_r���)K)E�5��k���[��
��ĹŊt�S)23x�L�y�c^�n�$n֮]�/*qn�"�c,�?Jqn�"�_�~R
�������ܹ��d��ɑ�s��c�fQ�s���Q�s��cKaR� N���kV&q�?��c�(w�@��TC�.[.zQ	��%y	��XQ��ٳg������łA�"��d��"0�J՟�6]�QCA��L җ,Y����H'C�^��8��ƌ7q�'D:N�4���t�S)��՟�����S�J��ٟ����KuB��7.�c,�e|e������T_"��F�>�f�Q�Ǜ��(��3N�T��+%e�#�������O�a����@����)hJ�***���mjN�1mb�E�·�z/s�u̅O�SR��M\SEQEQE�^0]�4�])Ջ�$����:��7�?��PQQ����$HEQEQEQ���>R�8W"^�;j��"��K5�K�V�򵊢(��(��(Տ>7o�<A��-�ȗt�Z�Î�d��������ӣ(��(��(�RJZ��Z�%Ճ�Ȗ�H�C�w2�uf;Y��4�(��(��(��ToFTTTtڼys�k喘��pm��Q�;�{1w�\�Y�R��,P�=�(��(��(�R�b�ߙ�8I7L��ǎ�蔚��lߑ�r��0�@)��-[V����3-MQ�~}i��U�֯_/+W��_����n�U������|�e�y4�A�I۶m�I�&�l�2o]�iӦyk'Ѹqc�W�^��,-�t��m>W�Niڴi����N-�}��^��[c7j׮-͚5��k�ʪU��X�7o^emV�O��`:u�$ݺu�֭[{�6�|�h��Ki�wa��biذ�w�-�\c�ܵkW�-�Λ6��1}7��u�z}ȥ����y����~��Kн��O�t�����;v���:�\�+V~�?Vd��׃����\�p�l�۷��3m��㏫<����k��������t�\ؘ��;w�l�kG��o��.���&���Σ��޸ҪU+��>|���}���ܻwo���-��{���FPxo���`����l��3>��r.}�]�v�s�}�8w�!�r���^�.���h�O;8ۆL�=���g�g�%�͑	�u�>}�M�6ҢE��6̜93ﱎw<�z�Ĺ�������l1�E�9���~�ok;�����4ƀ���俶.Ŏ�A�������N�XA�s�Y���)�}͹�46Λ�B̹S��T�Օ�K�î��6�1I/0_F���(��^�aÆU~��ʣ�>��[o�U�9�������_.;����?�Cqq���E]${��6/~���o�C=$��ߪ���{�}��U>?r�Hy뭷��l�=���^z���|PN:������^3��ŋ=��wޑ�����A�;� ~�a��0���������ߗ���a<X?�p�e�]���q�Q���/�.]�������^n��@Êk���;o�s^´cƌ������-�<�L�����)��"Ç�ڀQ��?��O���ۃ:H�<�L�k��<�����k��v�z�}�����������%�0}��w����"�#Fȡ�Zy0�-8\�I60�C�[��v�a��?�\_�6,Z��k��s������o/�\r���>ңG�m~�@z�'��.���y�'��rK����;��sϭ������-�m7n�������ac}�6�p����c�y�X�u �5�\#�w�6�4ƕ��{��0�,g�q������
3��'����C��o?������+��\ǣ��>E����/����޳��:49mx�7�699���2dH�X��|���e���^��C�>�`���|�=ό+~��.��w���^{Mx��Pa�������W4Yx�}�Y��'O��;����o߾��g<��O~�9����h�+��i��/����~肃�G�Ƒ �����SOy��駟n������������V�?��m>kE�_|��{��9�	Ldܧ������'���\
�w/ϯ�/ǎ�م��Ƙd���ַ����ĉ+��~2�Ў�~X9����g���w�yn���v��gK�d���X��s�=�#��D�6���wq��iv�]�`g昹�;���d���������sj��ߠ1���5�ﶊ�4.�����k�q
�f��\��̅�#)��/���%�����%�
�O<1Tl"�F/�r�x���,'�pB��q�o���gD�����_������ֳgOO0c$�����'j���;���g�ctc�1�� c.0~��9 n��O����6^h׳�:K�L��	� ��q�|�Zy䑡��\z饞���k�q�ֽ{wO_}��r�m�y�`��c'C���?�F��m}c��I���]��~z�p�a|��
2���>W�z��#�8B~��_zۯ��m>{�G�~�q��'{�`��wt���N���;�,f�m.Qj�&6��*cN����w�d� �\���8��LaΊ(!rd�@$g'�aw��o�y"r<�a ��<��������9:�e��vZq�kώ9����=c�/��6��1�I�q�y��K�(׉��t��~h��Q����<����|���8�x�/��ϙ�'!�*��#m�s����j����1���!�oa�<�^�<�a�h���]�4*Ιg�f�162ކ���?.��h5}�W������	,�����`��O��\�;��p`��T8��2޳R�{���g�}&	��6��/)���3%�"�q
t���C�!���wa�@��f�Q�Ă���5,(R���B �B$�F:RO?�t��2���A�7�����
"
�+�t<�� c<���x�����a�!�0f0�â%@t�֟��	D�����d ���ц(� <��B��'zH���R:"�A��L ��(� @ `<c(Y�A�\�/)�>�|dJ�%uԦ���>�'0P���*�O"v��$�q̘1�F��ם҂��5��%�HW<���vAS0�dӐ5����[8���~�
�_"��8g?D[�Z�w��L�\@q��Apo����y�>����]%�C���B�B9�#��l�� ���`���A��YHM��+<��q@�q�0���]��++^��g���	�O���g���Gy}��ǽ'���x�0L��%�J��c��1�kXLb8��8���]���6p�8W�c�MAM9���=OF��7߼�ﹿ\�	&xm@#"�,��d�������aQ�����1H�d\�o��w8U\这�F�~���+��ɤ��n�(Γh��c�.��`��`���n�?��(xR������,��:!�C�2}�y�|<))��+sί�-��؈[��æA�l.��S"�92��������$�:D�"�~�ɍR`���M�`�ϭv�p��FH�҅���=��8��E����GX�'�A�4�\��h��ს@�.`�3il�"����a�z�����HÓ��,��{��h#|1`Ĺ!CA�y�Q-W�#��	t����|A^�xɭQ�0!�a�z�1��#F0����ta?s<�D���o2p<��<���ԩSe�]w��	D��я~T%���F�a�����F�~���  �=�_�����Iڀ ���]s�;��;,<��#�H��'������
|� cA�v�"�"#&�1d-px����\ѧ,��u�~r>D�0��Gn���F��~�����	J�&}>��W�����'���N���ӟ�T�3
������qA���l����w��M�(�hO=�T��C�mp� �h�;E�-Qd7����3��?�A���0��Z��A�f��c�s��D�x��$���d���Sѽއ�8��e��2\x��Y���Ls҉�s����6p�.[8��xQ}2O��\���f���� ��Tp��pt�^gludpp�Yp,����ta�FT2���p��@��;�"�[�A�{�>���� ��wQ�R�>����Ac:�?ׁ�s�/��3��c�)��̢���æ�$���^	����g��9�o�'	Ɯ#�J�n���U
��1� xs�+	�\��/�����x��@��_�c,��+"#�B:��yn�5^����@�cW�`Pqp"?T��ƙ?E��'���\���4�I�}��1m�C �Z^֤��ii�9gؼS^�v?�U�0�a��6Н�Y�g=�D�������N��F�sCT0��=B�q_]G
�.(�4���x�W���`����������5pj`p�)�nVI� 6@*=}=_���,�I�5����E��4�����}C���K�0�VB ��rAY;.d'�6 �������0�}{<�w�qG`�_���s��{�c��i�S-� �v�6� ��u�1݀��4W�uPF��W�g�����ﶁ��60�ȝ��p���br8a���g�1���OX}���Vl�9��8u�7��&7�s�q�:�Sa���p��de!������p�$��lpl"b�dX��~�v�
t�+���<�m�
���E��� ������l��v��yo������>q]���ڎM�s��A���� %ڊo�	���%(��&c��;׹օ���3n�>L�$�0iҤ*���:��?<�8.݂��Q	t�^(��2M�K<<s�m��I ��ЇL;H	(�@,�M�ȓ<#i�ts^�'��6��^�Ƕ���xح�@��,�F6�:;QL�%v"ሇ0C�ȟ[�2�%|.[D��M���0+�ʯ"c��m=��� m J��`�p�
+E	�z7 !J�C!`�ᤱ��)B�xCZ&����x���}<�6E�HN�B����h>:aΨ|�O��OZ��M����\G�\�9p��`�u! ����8�SG�&ڹ������y���%c�ی��\C2f���\11I(*f��D������mC����a����y����Ϙ^h�Y����`���]�F>�@(�EJX�� 8������8�x���6�f�D�3��﯇�oC>��V���:�]�� ��g�t���S����0��ę���;���IP(<�Dѹ���l��y�����%����!��_ԯXx��r�q�sW�3f����	����)8�p��f��mp�k������p<<{�M��a,rz�5��@`�[d��s�pH ��{nk��� �9��a�j�Q*���۠�i�q����O������8��梤'v�����)�=_���B!��Q���}�R���M�anA;��Os+���1��v#��,Dj0V��|"��t�~Q��/@<G��y���#՞��V@ �0��-��	R�]ㅨ0F}�E�n�p�f�At���kr?��8�lj;"1�!Ftg���A�́��A�ב�e�c@
�����
Ak������7,���H�';ß��0�q��/J!�^K$ڝ�B�@�D��'��h�1�2'G_�ř�B��&h�_�c�S|�~�� '���!b���`!��Z��@|Z��U	��dB�����/�q�b�x�y0������|�u�|}�n���q�afZ���@���Υ���;�)Mٞ!5w�; �y?U�g�BHLq�ʢ����#d� �xo�|���3��V��9cz��y���,�$��:���Ȝ�$�'�/���
�1mˮbkn�Y��w�_�s]�#q�N{�z�;���q�+DY����L
�a�� ��;��i
�E)����a����~�W�9^>��,�qK)��9��n�e��u���%¯�a����j:��-X��.6u�Ц/c�˃dZ�ſdVPZ)��]�͂��G\0&|1C0��~!�)�z?��`Z����lQ�lU��P�K�c$�vS%�Ґn_(�����,�8��¨���l!m�Xq�hD�3br��*�@�mpz.��;����}�x@�<��&��_�(Wh�+�s�d�c�dPA�\��=�0�}�� ��
��6 �b�当)ڌ�MC��a^y��]��
��6 �ڀh!��5��{XH�.�0��X�>Am`:GP8oR�q���D�=�hv� `y�g�K�1��=�ԭ�`�!A=���d`������Ԥ�&�i�|�bo�f�6}x^2M,��a�9j1��� z{.m��3���d
�[$���f�aW	"�H=�6R��2!�N����������晎���9V��{J�)�@�r<5Ϛ��c����޷��'��(���+����xi)n��֍m��
��{��ޟ�i��Ej=�.OA�����9�b�W��b������BR1�_���j���c�s�U׏�e8���p��R���CD�^[�U�P+�|�χ+)|ǔ����]0n�,�:Da��ې��&��l��Dt�_�-��>��1����;���6d��{�n
��%h�@"@D	�Z�s�X�8?�|���+*P�݆ �[���e�o1&�)��\�'�ȷ/�p_����6�ˬ���F�}����"ҋ��6p.�@����~'8�qv3%gs{���w����p*�aUL_b\�ɀ���u��������]�Q�@'��f.�,ȵ�Rw���'����Q�*� �u����$����r�� ��r�%��]����5r�[�fK�	�CH�aƨ���3IJ�9&�ǈ!�W��rt�^�ԇ�q���������?R�q�gW>J��Eb�����^��4D�\��?w3Ӳh�舛*k�K$�TJ7�3HO��nۈ�E�8*��B�+��+�5Cy�����0���C-(�0���q�C��5$�~3���L��Q�?�D��%D�,5��Ka��ZA�����u�u�s;��Bq�(ȵ\S�����!h�s�.�/�?��8'옅Q_��ߗ��@�g�[�aJ=������0}�V1���Bz.m��G���j�����6s�i���₸�/�LE�ɀ��$8I�/$��y��$����D߈�r�d��t{�Do���y���u2s�����|A��������kF�@��c��q���.A����f~.�V7�M_*D��Dx��%�kۀXdUo���)*�1�1Kf�-2KA�\W)dU�Z\O;Wޭo�3�����qg����ডG�f��C�sg*�I��2�A�+8ly����S!]�K����ɸ�ɜ�bq.x�Y����P��h�2�s���-S�K5w)�@�,"4�(��Y�Ѩ�̾yk��Hu��'�(e�yL���$�ϩ�N�Kݮ�[(~�Q�`ϥʺ�� �!��D�~�2�%A�Iq�/�U(r���B�^~��%���V`ǰ�خ��(+T���;@�9��\U�c�s��gL�v�s<�}��Rr?��S9p2����&��F��=�O�� ��%��8�ܔUo�i����_�h���=��צj�$1�����0�1�H�\C���s}�@t��o?F���&�A�&������N6WH�B��G�
�L�N�"l��ՊU"�̑���w�;�@�Za�5b�h!SW�~�Rgjc�ʹ*��=�=�\��4ԩp�8�8v�Xܚ.��AE�f��i�V�������g�n?.�/�wS�駙
s�j�`��G�Y��+�AZ��d)�������y˼��h�xAT��.`�����ªdYa��g��<g�6�]��mSl1F4�jpD����7su"��;G�]�GP�`R��e��s�y.H_��y6�I�l�Ў7���5/��*�@�paXC��+ͅb���f��P�n��;��+,$HсX�W�i<���
���߹D='ےk���yZ��/Q=^xQE1�H���(�F�q�z����6��� pp` ��K#��6A$�%�B7��ؐ;��( �����
X��]ـ�[K!
���͝��U����I�=`(��$ǧ�;Ǜ�V�l�~�0�֝�B�|�s?�8\\�#Ͽ\cF2B�BĊ��L�Y��Ž�A?�_eZ+"���b5��B�П]g�
gS&e�I~��=�u�ZBt�� %����r1�I}F����B�!Ӻ�SI����#r�����
tڇ����*�Ԅ(�4�YE���ϵ���A���q�w.��/�l��8[Z͏��5g��;�x��U���󖃦��v�耰v�c�<�.�F_#rn����P�mpS�� q�L}ȵ�9��|��&�Y,	G��[�2����M�f=;�W��<��Gg�����.��1w7[nk���t�3;lݎ0�s��č ����í47d��T�=��	���-��1�ƻ���4�@w Ƙ.��uT0/	ϥ[��Q%�k`��y��ai��� �׍�QD͙S�/\��5SJ��k����a�Sۅ��G����d+�Zr)�FT��" 1��º/z��B��
1I8"&�Q�Ӆyd�g~�)�� ���V;&�Žu�_[�*.r��=u�ĸ� Ÿ���m�\Qww*"2�:d��m`,�Dʡ��ՙ]�M� ���j���H���E��"�n�$��Uٮ��l�L˭!h?���&ϔu�X.��*K<r�����z8�������������t#�@AN��S��ܶ�Tb撒*�fv�L1����	��%��m�N9 ��h5s������<�l�q�P��#p�q'��=Ν�)W�r�qb��ׂ���w��``� c�-�J��SX���6�2��6���I�v�3�uw�Ǒ�_W�kaӿ-D�]a�S�w"Bş�Øλ�%[_b,�8��d�uk?p��Tkq������9_�Y�p���;��vW!�J�=�Q��d\�>�=iߟ�����7Q�T����ϥ��$N~��T#:oݘ>ڌex�����q���P]ʲ���t�&[���
t��E�󳺒@�&�]�m��ߖ-���$6�N�D��Fw�Ź�TBT����`�8���S�z�鶤��a8�"$�/��r�`�g[�7"��"G�}�0�B����o� K�E��)�\'k�Ͷ�>~�y08�	�X�0�g3AԖ�߈b��kh�#�n��1sS�Q��p�84s��� �2ER�f�'A�1��j��s�9�Q3�-����a`�R��½ɶf2s�����蟓I��?���.�:3�����/]��>��\�\��p�K@ҷ]q��v�p� ��Y��5� D�o��6O��}fs2�T���c��n&���X�g�X�>�9#��H�f��&�3�Qבɳ���f����NĴ�,E4���K���_C���;��$ך�C�1.q�{�n�A�my:�5[����w�D<������0�Y��?��:�pd�W(AT�=����T)�������`<�G5�zN�.�Zh�qo��Cf����	@�	��g' ό���Y���?�Ʌ}��B@�P ��甍6� ���	�@�d�VCX4�l�^���q�p�����[�����:G�5�٠�<v���³�i��쟊�Sp(���Txtٺ�������������NݭFejV�J�@���z��
�h���!�e��@�5"y.
a�G�|�\��<Q�B�2A��h �Ǌዱ�y��͔�
Š���=F'[��B-v�;�8�� �/�Lm�0v���1Q(d�	�O+�p~����.�� N�*��a�`8�B��|ٜS���#��z�-;DOÌ��~��(&mq�#��
���P�I�<83�I��9F<e��AaϠ��a˰��@ց���"��BR�-��l06�A�d�3���n*%\C�T&3���`N}�*��d�-w8ɩ�P�j/L- C��U��,�0pN���P�0H��p�aU(�(8�ê�G	�� ����Z4iЧ)��<� B<�5|�@����\B2�6�x�п� rS�]ш'��]P�l~on���$�CЦ�R�ȟꊈ$J@�H��X�<��
Zփ��n������ങv��@<`l`h`|�E�����h/B�"}T�'ښ)m�c�+ט%�AT��Q�&�`��B���s>�?6׌��ϋ���h���˵��9��̈́�~���-��z�YC�O+"
�R�����G�����o��&[���j:����|�AP� �ɽ�8�r�A����\+�+ڀ��V�/�g!�D�x�pJ2�����D��"H��@��Г�M�>,�9�6�}��r">�C��3QH[��q4W9�؜'�m ����05(ly$�'�=���s�����`��do�X B��E�>@�OP��C�Οc��#S �F����n�:�7�ݶ��#�O�l��9�̄�/dj��k�5D,�\K��G�F�]��D�7D�y�2�?.���yK�w�,�3�g���>\xF�9c	�������8�(�ǳ��*���&W'mw�-׊�B�xg�3��9���U��Eݟ����$��f�;��es�𿳊-К��wx&�~�N�j�����ff%iY8e[T�+�����F��+^L����+�$���s	�F/*0gZF����e���1��^A`�G��@d���zDw�w�9Y)��
��6&�^"`n��|�XOT��te�(!�8�(ڀ�Xl��~!�3ǔ�XHGg+����L�F�s����@�<l��3�6�<saɜ;�ڙ�i�=D��6���dl�=�h�!Sԛ�<l���Cδ$cR��L}�bI?{h���P���$�p drrg��t[A��v�f�W�?����ӆLEq������~[�q�m�?�X��I'C�6П�����@�?�q?�4�\����9�s�	���\pW�(
���s8�������R&�~9ɵZ������(߀!�z���]��\إɂ֝�F�h��I��R(vy�B�@Đi��_�	������lT�+��(��(��(JP��(��(��(��(	@��(��(��(��$ 芢(��(��(�� T�+��(��(��(J�D������0�4i"�����˗��s�����(��(��(�R��D���p��^���[:� �ΰl���?��g5j$��(��(��(��)(�R�5k&u��-z?���|k�ޕ�?��x���1��߮k+�ݯ���θW֮ݐ�8}{��__����7m�,Ǟz��5�_\u�б��}O��G���=\��j[�=�]a�ع�\v���/Y�Jμ�����q�,�Z.?�䑌s�'H�֍+����/ɛo��X��iڤ~��������Q��ף,�?aD����~%W���Y�s����qG��~��9��	�|ݺ��{N���o~v�O��Og.���2XN9��s�4e�����	�|������.u�Ԫ���~��L�<7c[��#=��ϲ����Y�~o����$g����߀��_��T��ϯ�~�M�&�/_�gg���x���ӥs��ƣ�����U�ׅ��� Çu���ɧ>��~G����ˎ�:W~��?ߗǞ� ���$�^yH����o��O�'�qvީ�\qɁ��/_�FN;���s�GI�.-+���ݯˋ�L�z�?��8i߮i�����W�����~~�}��yg|����g/��F�3�q9p��~�n��O��@F_�9��!�����r��O���_���
tEQE)�����K��Y�ڣO��_�Zo�p�����ШaC�o�@�֭�n�wݺ������!���ߛ�S�����]*��8�+y��i��:d�*�6����ӥs�*��⒫�%�7;��?Wh>��ͱ�d=��]{J��d�=��D?����>�W�skԨ~Nm�գ]���ء��x�K����������u�2g�п�]�*��٣���7ᙂ��6����W�gm�43�Y,��y��s��L�Ϟ����ʯ��t����P��j׮-w��v��w��ܚ4ih��̎�͛l�w�{��)����A��v��~��y9�i�A]̱�q�}1g����	�ߡk�s[�f}N�i߮E����iѢ��^�>�ox��5mP����M��X#v�^eLyc�g����Y���ҳʹ����8�>ޯO{#���<���T��ۮmss�E�(��@��8��%ڶm+��$�^��_=��S��}��ҵkW)7'N���zJ%i�9�ے��ٳ�G��7F��Z�j���.��zj$b�֮]+��s���G?�M�6�������J��9s��~����k�I�پ�̿����0��+L�-�ܱE4���>�yd�}�ԯ_Gzl�J>�lT��ٶ�8/���w���h�b�Q�z��(�]��ͥy��l��؎�����'g�}���֌��""~��:}Hd�s���	�G��}�Nͫ��b�v���8�Z�l$�����8�D$!x�G�����z=�/_.����c9�;��3��~�3����EQ��~��'W_}�$��}��5�\�~G�%�s�$�w�<��s���Gn���D�s�޽���/�>}�H��ޭ��6���yw�6��]��s�N�넣��˯M��1G�L��[/Oh��bۈ+�����8ᘝ�W�y.�wG��8�;���7� +Vn+j{vo-#vέ�n6xG�,<26���G�&�3���������Y������eÆM��n���<'J Ȉ�>�ҶE~��9T��~E�z�$�Ջ�8;�,������~6�+�;lG���*У��?@Z�j,�o;��c�f��ь�8k�:�ǿ�N<&�6)�Mq��%;��%I�|��*�%G��k�X�۫W/I���vn={���R��I�kGɨc��MD�'?�WzE����q��Cv�=�I��#�.�ᾑx�u�ˉg�'��}�I����k�,g���<��$y��w�CN9~xd�!���"�~�JJ}�u����9S�b���c>���Wupu��ߗz^(���ޘ.S�W�r�@�m/Q������~[5��>@���k���|0�Y�pe���{�H�q��L8��]�Gޫ�s�_yɷ#;����'�S%���_=�;Үm�Ȏ��e}�e��.r�i�e�Ἰ����e���̘��_�9������%/�o�6��Q� �*Ы)̥��Q�4h�A�(��­�!a�^aq���xNi�������w�.�̓�-zQ����P���{��2t;y��	�v�z�`����Ky���G���<r��q�2㳅^�����	�(�W��<|��8o�+���O�w��F���͉�r�����ޖ/�-�>���yg�y�,�c�z����d��{��9�QF�����GΖߛcP��^�:�ȩ'����>��oI��m��G�z)�L���{V��];��g�y�w�>?G��>}��;����4[n��0#�;ɓO}"�V��a;u����W�.J���Y���9^��ڵi��#�bA �w�Ir�}oɋ�L���v�%矵���������3���g/�2P�>uw�%Mח':�WǼ��7 �O;iW�Y�(q����W_yk����͛K�֭EQ����/3f̨�~��ѱ�]�}���ꫯV~��ϖ��Y�`�\p�%=���ǜ�����M�~�i)�\t�E�V+���w%n���v�o��A�w��o:Z�(�����mq��n=�-n�DI��~�O���fa�7�I��781p�E��+2�z�7X�)lq���n�7M�4�+.9@��T+��f��2e�|���2w�\O��[�Λ#߸qci׮�W0���ҴiS�i�����OJ���K�7���(J��4i�|��7��U�VI�x���+�_�~��������Ǽ��s�ܸq�Jznd4�Y�+��(��~R/�1.��N�]*�#�)�Ct�^�z޶a��3g�g���%s���FQ7EQEQEQE)'��+W��'�x�[�Neb*1:4�\g��ӧO�D�/� ������rdD�kM�D;�	X6�Q@EQ�a��]�[ߊ>=�[���bk�{�4n�H�䣏>��^zYEQEQ�@*��/�(��{��X��_y�r��g��ŋ����L�0A.\�x�夳7j�Hڴi�E�Y��9�l�u{�]wy�؈|�G��Zu������I������(��N���/G�\�[o��h�~�a�F���;"m���<�mq����ҹ�Ϥz��%9����m�`Јx�P�s�^�8���7�-n֯�X�>w�5�񶸡0[��t����8/�:�dm�}�[Jr���7��%	�J���~�m��[o��	�V�Zy��>���2{�l/"�k��cǎ^z�1�#�]w����e�]&m�F����(��(��(���Bj:�����^8
�5k֬�wD˟y晼�G��~X}�Q/���/�|P��N���K�t�=�]�EQEQEQEQ�(Z��>N�t[��[�n�G��_~�̟?�Ko�r=mR.I�3f�\u�Ur�9�x�ީ���_�Rz��%QB�=��-T�W��"6�v�k���ܹ_��(��(��(��h�ީS'Y�t������?��d�}��� ��ȹ礴������͓SN9�[Z�k���n�Iڷo�q���k̍W���?�TF��Ujd�{t�k�*��(����~��I�Z�
��%K�x�CQ\��=��C���v��_�B&O�,q�����Kk�S�[X�9��m�����-�v�7xky׭[7�c"�݈z��~��,��(��(�����\`� ����"�YC���|���9��|�Mo�y�i�ٸ���=o�{��M?��Sc9�|�9ıD��(��(��(�R>[$�����s�W��-W
�N���[o��#GʓO>��c~��(��������REQ�C��k�JR!���R���իW K�@�'�u�[�n]����r�Ay� Dѯ��
Q�f�2�d�ā�;S�a����N8Av�}��2�EQ�h�F����婧���ӧK��hw�v�DI.�f���>�I�@Ǜ���O{^�rz~(PG
?���~[����»�(՟c�l+��2Dn2ۊx���Xޛ�Bޟ�R%�����	tEQ%9 �ɲ�@6"��ߍ7��C�}�С�<ja�СC�'��ox�bmI��ޜ�/� ��~zQ�"]�]��
�U�%��>����Ұ$Ǻ���U�+�� ~��eȐ!�(��$���
9��<��-����V�B)Z�s�1^Ty���x��W��uI�7A�s�N;�4�!,�lc�rVo�k�G���(�f���^�̨)fܴ��O���EIӦ��q�/�G��F�/Z��K�۴i�(��(�}бc�*S���{oo(
]+J�$.ŝb�&M�q]T�`�w�|��Q.�z���{"�o�k�+�RzH�[�p�$��K�yD��A��dI���
"r�I��(�RS��&���B���_~Y��J�$N��&�������S�:tEQ%�|��߮R���*�EQ��ӱc�J˖-�G���(�ַo_O�(J!$N����-��ѷ���^�B>�x��4t�����>}�T�^�=EQ�d��l:��1[)��	t��sГ�4w�\Qj��.X0_j���EQ��r�,QEQ��O�ҥ0�bH�
��St!���T�X�x��X�[	F����Ϩ(���TGKI���Kj��X�]�9�1AU�FRVPPEQEQ��D�:� �K����b͂�3�4MV��R@?3f�(��(��(�R:'�5j�	a�$F�9?��вU+iа��4��(��(��(�'q�u��Dѓ6���;t� ��(��(��(I�i���׼B��dРA��'q�K�.�����'J��6;N�Ν;�Rs�~� iѢ��4t�5EQEQ��vaSJC��߉�� �U��'4HNj�,��@M��8��gPQEQEQ�Ғ8�޸qc�ٳ�̜9S�Ě5k<�ֻwoQjS�M��JMcÆ��(��(��(JiI�@����K�O��E������� ��F�=͚5�aÆKMc��PEQEQ�rS�@'����v}�u�J�:��v�=����O����Dt΃�u����b?\3�NQEQEQEQ���\s�L�0����;N��g���ٲeKO?��s^q�b1=���������?2n����۵k'w�}�(��(��(��(5�D���QG%/���,_�\Z�jU��X�b�'�O:�$QEQEQEQ��H�@'�|�1��<क़S<��������[��+��(��(��(��X�Gy�����2y�don{)�oܸы޷n�Z�:�,QEQEQ�rѬY3/�ŪB,E��p1v,�W�Z%,��K�zu�EI>��<�^z�\|������t�zܐҾd�o��ѣGK�&MDQEQEQJI�Z��k׮ҫW���I����(��ϼ�(JrI�@�6m�ȵ�^�	eDs�"�A�����+���}���(��(�g�ȑ�-w��zuf%�4o�\�I������gϞ��G����EQ�dRE��
��K�9�6��z���%jz��!�]w�W1~ѢEҴi�X���e˖y�'r?bĈȏ�aA���kW� �uPEQ���%*�^�b%�:u�!C�D��-��Ç��'ʧ�~*��$�*o���z���C��qһwooy�n��P��(.R��S�9�_~��x.���V~�<�B���(�������e�ԩ2o�<ρM�-"�ЧO�{EQ��m۶��N;��|1����ؿ3g�EQ�E���:t���>(O>��,\�P6l�E��L�`��{��}��:�\QE�ѐ���SOy�ZY�$2����w3�����0��#>��X6l��v�:���M;lذ��UD:*��T�d�*��??��Se�}��`{��w=��ϙ_C�/a�����r���gN��'�,�EQE���N����sW�����W_�1c��QG%{�g����/d�=�v�,��~�w=�xi���8#�4}��Z�;� �KQp<X^{��/EQJK��e�����Jf͚彀\��q^^֋�Ƌ�qn "����~*�EQ���{�GƎ���!��l���/��c�u�+���jѢ�7���d-��)����r�Jρ�]D�!+� K>�����G�?*�s���S�)(Ӆ�Թsg��/DQ�d�Z�nA��y�r��{KG�?^fϞ�
��xI!�y��"� �w�9�Q�PEQ����#��-�]^y���?��CE)lD�
k^����bl�=�;�s
�Ι3G���+]f+�`��|��Ş(竻JA�n�2W��$��t/$ֈdSEQ%w�y�/�XH�'��������($���:�	���<��?��+���S����p��I��K���?(J2�6]QEQ��A�Qx5
�N��c��O�SMu�j����ڵk�kFEf��_�E�m�<���s	R ��� ���'O-����f"*AD�V���SEQʏ
tEQE�����{��L3�0aBY� `��5��%D5�Ť��E�Y���t�/Y�$k�>"�T��G}T9��?�g �z��C�S�G穗"�a��!�S7s����N�;SO�&��(J2P��(��(5�?�0�}"�!�I��:5n��Ht�@:ԋZ��)�D��R�
t�`�O��%J�O���.�
�βz��\Ȥ���D�6m���}F�g+&���E)-*�EQ�3eʔ��9i�$I�$�O��C��&�������=GB�HyD�).g��;�W@�O�8Q�N��U�&���;��ùB�^)-Ů{N����s��₊�$�J"�EQ�vm�`^6������>��4֬-�F��e��բ(J�0�9���Dr��^�y�N"�vM�N��u��ׅh9N�b��݅�_V�[�.ӦM���OT݂�`�w�O>�������,�ǆ��{IT�� ��P���E)�H:�.� ��ⱽ袋�:Ë��o�����T0^�2|e�B#	Q0a�xQ�Ccl�:W��D=���׊ �ҥ����^7
�`�}�VR�Yf������b��3ŀs��޹�D���@��k��N;UF���w��������͛{�Iu_�����Že��Ȝ`*��(�&��o}���r��R��1�뱾��$C�����y"]��l0.�ㄴ=}f%:�r3~g*zU,̳&M�0�v.."����{�K��/�IG�@_�6���e\�L�	�������.��/6�̙3E)/�s��@�:S�J!A��i�6� ynT�+J���
/kR�e_���,ҳ���TE�4�皞W��}�Q����s�-z�w�4l��(VM��g+j��(��v�J><�1����n2~�xo�w�@8���x����~g��
m��qPd+6��`̘12l�0/{�B�8~7w�\Q�����:S����⋢(J�@z�;z�����C���W��'�.X J͂��V�[k�BZ�?җz��^�(��$3+%�hR���}���8`L1b�'<� $�t��e� ��!��$�UZy&��s��	G�Ǖ�@w�ɥ<�m�ر^u��;z?�I��Z%�,�� A���}���B ���oP��D"�ǍW�jh&� zꩧJu'WA�ڳ�����^��5h�Jua��Үm�{��RJ�Qt�0��#W�#rI�f�O��Q����ӧ�����+�Ě���EDڮ�TڎS��_��q�k�7΋��u�]+#�O;�x�X"�52;(��_����C��mZ{�Y/8[2Մ����{��o�-�Ԟ���H:/6EQEQ��z����}�~�K���tJi�O?��g�G��Q�P��1ɺ��e�1c���=r���y�""�QD��߿х�b�y�5UHwF`ٶf*}�H��{�Y��@;����Y��?����B��B�h�Vr��""��q�T%;��(��(5��|�<��Ñ���#��*8
��F�g͚�s�7�1��mK��Ca8���>(Y�K��[g�o�2�I$�f��i��ٳ#s��t�M�8�2K�{�sBA9j	ϷQ��w�]�|�M�Q�B��ٕ!��Q��(��(5�����[R��i1�vEp����|��/��1���<)��������ñ�l��^/D>��z��bwDW��`Z(SK��r�2F�� ��`�"=�U���7d)��]QEQJ���ɝ�K��SN��B����O����.v@\�[�n]��Q�\�����v�w�;[4q�h+dy9Λ9�6՝v�>��X8D�������8����E�B��|%�����`"]k(J�Q��(��(%��������A�?j�1jGc0ǳY!��~��#�<"���z������Q�FŶ����f��\a�7��R��b�0w8�C�Bʞ�k��V����ګ���e�lf��������8oΟ"qڧ�0���s�����';��q���-,ga�B�� QO�G�g(�R:T�+��(J�X�|����Lo{��	r�:u��R��D��O>��L�<9T�#�w�a9��ý��qC�3
Uɡk׮^�?עkݻw��?��B"��@`���T(��D�9���,O���/"�@��o.K�)���5|���W�Aܳ��"n�
�b �c|��g�(JiP��(��(e���'˽�-g���$�,�t"��|�'��?�?"�r�9���L�:�K�"�,�6a����s�?���X�{&܅
������ܫB*ss���3��B;�^����R����<g�S+�+JiH�@ǳX� �w�? ٗ�Ҷ2��Q ÿ^$/s�+��(Q��K�)�-��MO
̱}饗�NF����˕��U���$�Θ3g���ܭ[���P������_��*�sGIϞ=c=F6�^���҉Z PQJC��~��'�>�lA����F.���*?cN�c�=��gIo�#�w;���r�M7U�����?o��(Jue��M���E���m����X�.�(nu�q�?nH#��Ԁ��r�
*W�À���6C� �+ee�4��_
���ر�����S%^'�K^૯�ګZ[�h���{#��'��EQ��<�mIdԨ�Juc��F�j�#:L���9������i�j)�s�s�-_~�����5�Qo�Q1�7����@��ݭ�_D�����vzJ���� '��(�Pc:P��o�q��IM�宻�"�����u���IRH�夐J*)�( pP�"�}�^i�\���p���*
���
HIH��;	�����|��?Ι�ev�������g>9�g��ٙ��+�OQ���ƾs��&�q_�[�j�*k�;"��Bf�x>��������!B�,n����w�����B�$������?$P�Y �^�NF���M�6��pT�@�D�ӟ��>�����!�H&G�hb|q�]���I�O�����C�]ٳ�8e�e޼y��D���t<n�s̋n'Н�_�Yo^�ˍ��$Dj�3�����*����@���N:)��|z��Q9rd�_��
�]w�]|�ű=v�=
:WQwڶmk�gώ�1�x���+��/���.���pۏ?og�� kղ���u ��o��9���
h���㳂���"(���7��r�-�����7���q�����v��eB��P2��B�:�����p�	Vn� �/G�aŤ��oB��gwȐ!�D�w��*ez�he�[a"R��Ҳ����jJ�9�ad�y���t�L߻woo|\T��$eU*�^����-��fƗ#|%Ѕ(%#У�L;'k'^�?�x;��S��g��r��m�24q���.�I};�ᡱ<֧��q 7�\q�)i��2�d��e����;��._����1W�{��W#+u���CR:����οu�c<��-v�}R�� �6 �Kl�m��}�ҥ:>�Ha�D����&�P ��Ϛ5��=����Ȣ?���e�L���Q�q3B�J�����u�Y�
��>��z�g�g?���EL�X��/�~���`7�p�%�GyD��ĩ�Ae���w�{�-[敠��S�[�lٜry;$i�IY����7h$]Hgʗ+|6M�4�q��\<��WT����>���(��"���@�Y_x�Zn�~�%˥��G?���}���'�ؗ��%{��G�\�&Eم(>�ׯ��Ç{��"0n��!�7n��]��l�/�J�}�Z�b�0����c�f��z;RCɺ\�s	F�8�:DY�uh�
&IiDO�j���y�W�uI���L�Jǃ�f�u�z�%Ѕ(%sd�v����eժU�����בUz����,��=�\�*����O~��˅p�B��zn��K����?{[9���k�B����\3-����xu!�@�3�իW�� �]��u���+Ѓ�#	���+зm�f�;w���~D�L=}d%[�,t�;��K/����>+G�V��.��B�|	�e�*h�����Q��b
.:�.[�>�`eˁ2i,�Vh��Z��S%�JRڤ�(G*Z�oݺ�&L�`�^{m�u7�t�=��CV	��5�!�-�"j�9'����ik�.,�y�Q�]�{I*G�2�'���|Z)��L���NЗ �00z��H�<��kH!�?(�Ny6&/�ȷgs��.��z�'�#.��r+wC3��&����x��ߛ"��0��O�yn$y�WL?���|��&�"����Fl��9�X�;���Đ(*�B�.�,X����#���.�lʯ�y����ri	,u)�'��t�c�=��%t�z\���H���+Wڼy�"�_�8��.��������BQn�~��v��כ��3g��JEr�?�oǌ�0����6�]�6��,��?GJ�Ìq3fL�ƍ�l�`���`ٶ��SWK�'� \0��@��ר ��S2���������Yu!�(7z��i"�W��1�O��̻�P��/d��#b��[�?�<,����~���s��?��ݏ��K/�d]�v�N�:E:y 
4qB�� �~Nn�2�?��:�
!D�qH�F/&�W",������;^�uoN���k���|�	�hѢ���;O� (E曖�իW{���/S�;m�܆ϫ�fn��*D��@�_��^����W�GM!ʝiӦ��X�0znذa&JD%�~�@��2sL�p�.��)�؟ɮ�Sz��ر��@�8oŊ�?e����e@Ԧ���cl�@��@�Dtd�W]��P2�2�l�5k�佸�@�"�w���	!D��`y��M�]}��&��P�>�h�g��-ZT�;�G�>}�r�t�E�:�d���9'`1e��\�T> �Y9S�V�ZD�#��p�����,	І0�|/p3dȐ�����/D�(��\��e<���@8p�	!D�P��.�_�k��}d�-���7�eCe���/_��2S)@t�)v�/^\������:o�,0�|&\Q��oX��/#�׭[g��� �2U�Z���������x��۷�HN���~ń}d�������8�;�? D�(��pn��F{ꩧLQ�����k�s�ڕoY1itP���UY%�[�n�x2�ݺm��3�d�����Q�J���$���&�>`� O�DY����X����s(sw0�]�~}d�߼y�n�d퓒!N*���s?�ۆZ��
�.!�C=�ĉ��L"�B��e�����í^������|������wl���c���t��[kL�~�2D2�Y���^t��d�Д���޲eKd��4��+�G���G�����@���x(ehy�
�ٺ��;�m۶y�n?͗|��	!8�>g�;�����T�8_y�Z���u��/L9�(̬U!Dyp�]�z��s�7l���y�G<��TB�%�����]��8^��mzÆ�(q�ԅY�y��~xz��2�.��s (��6#�������6T�?��@���0u���ߏ�
�(B��$N�}�r�,'�\���R�BT���T[�d�����ƍ��5���D�/_�]�g�(g�������vbD}��sLu)>��CQ�����'��(��x=~^{�5y$��
�(zԐA��
�E��Q8'�E|P]5:`!Dj�i�M�����]ۣ쮛�`c��0���ڑ�����k�z���w8��5���7�I�9%��o�@D?��
c�^�zy}������rP�^W�N��R}��Q��;TT���r�Y� ��o�UPQX$�+������sРA&�"3[�����=�������M����?�z�����Z�i��/,�0��0�ҥKu�cǎ�P#kYH(�����cW��z���9��#_���@��`I��{8�J��5�@B!���~l��v�M���L��R�Y�fy����v��\&�Λ7�PO��_�j���ׯ�:ƷN�<����Ɋ"	 ���T��~gf#�
1?��a_H�@�w�ߟB���@]!�(k�6�Z���~�嗽tĨ_Df��2��l��?�C�;���M�z�)�?��c=#�tlڴ�:�4��������N��@=��۽�����]9B+E]]ӹ�5k�Ժ�J�Q��ѭ[���֧zB�h�@B!�D���L���˖-�+Vx}�q1����j�x1�"�G	x\�f<}���:��<�Td>AW�t�A�ݵ  ��������^˂4��0����
f�ق�o߾�@�w�} :w	\:�.��]��#�.�B�C�g_�d���A�"H�(Id��:��Yz���pB/�-�p�Z��-k���{��q�����p�3���!(&!
��B3͛5��r���D�B���G�	_�ru2�;��;�Nƶe˖���ɜ�9�?��H�7a��c��A D<H�!�10rxW:������N=��5i�)�A/wT}�����H��9��]�v��1"�q��^|�f]�@D�����:��}������ �p������9lذč]�K�.5!D<H�!�1p�wO��c�L�ϸq�j��օ�S�dz�����;�I?���E�ͬr�� �����̑ǭ=8��ӽF�E�+�={��R�}�}!�9�"Z$ЅB!
"!�i����y��@�e6��`׮]��)��= @0`� O��af��E�$�ī��ꍿk۶��T�ȃ@�x�@B��{���c��1_BTd�1�b�;c��� �FC�1Nm�ڵu�~���;��|tJ��%�fv# Ea!XC`�y��d�`,�"^JJ�c�B��E��b�䆓�g2qGB�� �$D���۰)�R�J˹?,�q�g{ˍ����7�3��H,\��O'�Mz�0�����E�;cܸo�{�M��Ο?_&`1�����ٳm�ȑ5��$�8O7PQX/����g��r��1�FYX*����-��+{��"��BT���8q��Ey���UN,ra��%}ֹf�����W�`k��#S��_��}���S�L;p\;��S���v�c/��͜9ӎ;�D�t��ڕ9�x$V��5�.���4Ȩ#�پ����ĉ���K�|T!D2y�WL�L5���Tb3����!D9;�d���9�A�+dÝ@����37�Eq�3�6m�g�GB�P*���ٳ���9s���A�l���N	.!�K�:}QW\q�7��.p�;묳��N��������{�gB�Xe�و�y�H�[eB}d���Ej�#ɚ4i�e�Î)kڴi��*&�ꓱ���S�N���"��<�TP9@�;n�Iy*>��s�z-��J2���j�F�ŬY������$J��{�v��WG6BȪ�k_��N:ɮ��J۰a�	!��.}��$������v�-3!�B'�)�g;L���G]���Qd%̳a�Hg����_�|���GaB'��j
|r�Q��A�s!�A":��������;�`�AT���n�A%�B�j�~�i��K�QGI���_��&��	"�s��՗����Ƃ!z�N�p�o$'8���^��~�{���o@^�S,Y�Ąɦ����/�K���0o������G���B �;6!D�ٶm�����݁W��p�l&��r�'s޸q�����Ѽ�ش�r����(+T�������8Ĺ���M7��E�.]jBQI�@�4����H�)=8?�� ��'�5��O�w>��Ts�SA�R<i��!�"=E�g�y��w78����?��.�(���B�#'B!��N�������M$��g̘a���I��h�s�B$��l��5���B$��	tf�_����'��Τ�߭\��39�̂3e[�j��cJ�O?���ѢE��l����M!*�}"z��"}���^?zǎ3Α�,�u���,Dq�s�{���x�T�/�(>E��8O�O�X�L�!pa�;��Y�n]ڿ�G-->|�W^?}�tB�J���1cLd��(9�ӽ�Sǣ���G��������;"�
9~�����o�m���3!��s�gJAP�㭀�_.кLZ����Gyd��)x%Dr(�@4h��p�	���>s�LE�(a�t�b��~�WI#j¢���ϻ�X�x�no�����O2av���W/Z�ݍz�7��x;�*����\��b<׹�B$	'��:�u���Í�9�G��$��(6����CЌ \���$��WUU�g?�Y{��gMQ�<��C^��H�B�V~饗��s���7��Mf'�x�q�&�qC�-�m۶�&�̝�P?��
QL�UH�3|�!ЙG�GZl���/H�Q1�Dfh��t!J2,Aw�`�� K0в{��X�z��D2��:t�~����ٳ�8L; ���2�B$���)����ȭX���J�qB�&I;�$�+>[��9���?\�����:8u����� L�B��1�"�lܸ��[��^�zE>Þ�LS=�"9�.ЇfI��+��o��	!J��'z*����y��=��#ּy�з�������X�ӟ�$��)'���N����?�5���u���.<w������4�N�v�����#�17fR�ҥK#�Ib�ѐ!Cj��}�ݜ�����;�]�����?Zh�4
���rowྊkԏ�}fz��?ޖ/_nņ� �YL�<+D~<����G�d�:물z�ƍ�-,�EFm��/TR��ܣ>ׄe݆]v˝��s/��G{�2�B�j�-[�IY3F�q�dҷoߞ�P���Oi{�o���2J"a�?(�0�-	�+�\r����رc�s��.ԁS!ʐ�6گ�g�}���L�cҤI�ZZ���"nذ��uTKQ
���{6o�<�[�}�I�&^�wkz��=A�LkC2�l�o��� @�^�,�6]��� �����GyĦL�R0�!��a����9��1.A.J��;w����~qW�Nh�,x>��\�b�|�H(�	�h��]��\p�w��@"w�8�t;��sCߞ�;v�$@�M׮]B����.�}���+���	Ȗc��)�+dߩ�$/�H&��{"P�"�������'*��$>��Cv��9����e/�@ӦG����Փ�X�q⸞&�Cѕ�{煏>�����D�ٳg�M�<ٛLУGo>z� �׭[gk׮��!Dr��[����Z�ψww?��]ֈ#Qh~x��	D�@\oܰ��*�)ʏ��u��.m"<���g�K~��І)�m۶m��R��Z�h�	�t���T`����f���<��6L<ia�0GA�!D2�Q���-ר���($�կo�۴6Qyp��ڭ�m޴�>V�K���׳��-�������]��:���ְaCo�b&�i�&O�3�
ڴi��FW]�o����	!ʛHz�%�E��w�n�>SQ�t���v�|Û�*D�����8��Dy�P�KFq��KwU�:&���"�(�"ZЄaL=ˍ����)�I\��މ{	�pt��-��<��OEv_���v1!�eˣ��k���&D)ҼY#��Av�����s�ze������q;�j!%��&����&T�LL��$]�%��w�{ ���0a�M�>���Cd�[oق�[&b_��y=������/���z#sa�9����bp�w�ͺ��y����'���*IB��~��'xV�3ƛx���>�4^!�H%)��E¾�S�|�a�{�y�?�7I(�fq��kX�fm�^C�6m�~��U���|��ެh��;u��]��=z����T�ߗޡC�TK����:�(��66>cZ��0�9���y��7m���
�
!J������BQ��u�����e������y7v~}���Σ�TC�w��ŘTCEVӦM������A%&~-Z���y�1��ќ�m߾�wߣ]�v����m۶mi[�"iH��|��B��c��uE�Vѳf�{���Qj�v�w�G�m� ��s�NɠI�&^@�y	D�*������D0|ǎ
�	!��B!J�L�fdJ�N�jC��J�Ӂ8[�x�'�Eq���k׮ֲe˂>���F�k��f�7oVE�H$ЅBQ�˝)F��	wB�R�)S�x��-h������5^��P�NK%�q�{����{��W�!�H�B!�(	�N�#��������[�PgC�S��F�4%�d���A���@1`�6l��S����!DR�@B!DI��w�U�kLV�f�:Yr���=1��b��B��az�Lǎ�^p��|�3����l�bBQl$ЅBQ,\��Z�j��ts�ɬw����ȸ�]G�#���A���={z�g8��V��M�6Y�@�{챉Ț���g���^�=-�MB	t!�B�[�n�6�ի�'�3A��~g��L�ˬ3z���B��9r�7�-.L�b�c.Y�Ē s�)#O�3c�`cd�|�]O����c!�13�-��m0{�l�
!�F^���;8rr� �fzsR����6�c!�B��	��3gzB��:�<U֚Y���fC�]/����!�?�裂�8��r�����ݻ��IG,��oi?�� 
^O�`
kO���F�>ג��͛ۨQ�l֬Y����lx�G���~S�*-��$'�N4��0�y"�<�8	q`�DH$RB=y�9=��Ñ��e�MQ�<��Sָq�зg!|�@a���B���G}��>J������2��k�z��T7Z��Z�ܡC��˘խ\���eӬ�(�&8UUUE`��#F��Y��d�������`}�3;Az�Ɍ�a�"}����|hۈ��B$��aNS.�[uN�D#i�"r��=��cB�����7Q~w��6���Yo�w����I�+�$X�`��I[\���4�����:,X`'�t��؈QʾY��B2Wq�0g6���j���֭[��/A�"p��!���rw!D�����A�$��oz'�8LRDeAI_�Q����Y8���y��O>)���b�#QJ4n���:2�8�� $!��sɘF	�l#��u�3��y�-������И�RS��q�FϿ /2�.��	2�C���'4B�EV��ɥ��=���s���NB�^z��3&�����P'���:��ի���C�b_|�M�<�+�+�5��5Ѥ��O>�8��ݪUK��}7�k�뮻L�׷\�c�(�ƍ�z>�]�vy&qd��_�Ž�/� ���j�d�I��u��m�%�LI���-]�Ԓks_>A�*U���&��!D�OT��T𻨢�(ȶ�}� ��q�Ξ��{ݎ3�<��ϥI�d��M�G�y�}�nݽ��b
t�#�?�u�6+m>����qA��W^	}{�:��$@Yf.��0��|f�� ���W_m�&��Pɂ �ː�=��z��׫g�ʹ��	�e��q^��q��$��=��?<�0w��&�T0��27���'�lB�Ҡ>:��qP�hu6p�d��I9)=��|�sP�'JŢ����Y3���C�j'N,�8��֭_�����x%�^{-os��{�k/�4i���"�<���w��&�q�1�Dz���y{�ŕ֧W;㴃b�(e�r���l���.NPk�QI0	k`�9oٲeE�R!=c��iޙ�e�v�&M*��B�� '��QXʕ���I��{���a��'��ؼ��;y��|�A��YY����^����Q%QӨR%��j���x�v��[�|�n��t;��L�F�Q��s7%ӅtL5�\:p��P�]�z��X��Ʃ!ҩ&��1�ד�nB�7�e"=IY�8��DeC9�!C��I���4Y�CQ�$?�s�λ����{�ڵmj#�w1�8�S��F�{��UWݻw��A�Z�Ĺ�`��U�����6ڦ��B	�2��?�~�9�ؓO>����z�wT_fA5���E������hؽ{�F˼�+��}����
��<�ch;)$��z�������?6Pj��[�d�.v�֭�r�{������fH�������rZ�>��_�!���Τc>�5I����ٳm�رY���2u�TB�B!�.J��u�m��J1������
��}�C�U�Y��ز�x��RdM�I�Z0"E\q\"����Q��5!{�m�.��y��%��*��)w��r��(B�B �.J��6mL�E�=�bC��]�vy�m1{�1KJ:f���'�y=�lٲ�D��^�j�r�cx���>�)U�X&�p�`*������K�.YoG�U���Klڴ�+e�DUUU�:�+��0Q�H�W(���ӟ��~����O�WF�:�rHB���yO(b�!uxޔ�F�W\��{��P<����#����qcC�v���$A��ag0���^x��ŧ>U߾���&r�є�fd��9Nq�֫W/o$�ʕ+m�ڵ&�N۶m�f����O>�k#�N������ՍM�`Ѓ�[*�/��Le�"�H�W(,Z�9��C��(y����K߽ ��šy����fM��	c�����y+]�t�~������>�H��SO=emڴQ=,�r��{�5�X���C��ꫯ�}����	�k��v[�۳h-�@�ҩ���ֳ��mL�F�N�<q���!��}�����_���S�F@��@��6�m$%�<�@G��Z>� B�����{�V�|�����#&%��G	ʻ�;�m1Ӻ��+M�Uʌ�$s���lԈ֧W��w=(R�SBಝJ��g��s�s�'�N�{0ˎ�ܳgOQ��>���+��*c�%�qҰaC��c��LJ�c��ȔE��"N�.���s"+�q��P����K��<���B���ү���c�L�s���2Fn޼9m�������J�dG������"L^)gl	|�dr�'�C[��yN3B�tԧ�+ݼ`"�Q�'QZ�K`T�#�I�q��&��<��o�!�������ܱÒ�f�җ�oݺ%�~H!ↀu�-�/#�w����>�)S���ѣ��\s_|�v$�{�T�	t*�J��%�m��c�� ���g�A����D�um�|;w�u��yn�B�dS����.�,�/�<���?�zq�
�9��3&�ue��A��[��E�'�����%�sϿ��>�������l�A"D�BB�_NKKX�+Z�0�:�㪯#��C=/���T𾖺�8m�_��;�eDoж�k�+�'���6��A�c���{/��Y!J��&q���o�w��E��Q��/}I���A���E���Ӽh!�(֮Ú5U%W�p��ʅ`?t1[Ȗ,Y�rM�;= ����O��0�!ۤ�����#�@wq@���'��`�&�G&�O��aÆ��/��	|!D2���N&k������'���:�+o�D��BQY\{�9��5	��\�Aïb��*�$;�4�Ø-	�J�l��9\̅3�z'3�~��QPxG��<�p�S��U�V�"����H���k���\C����w\p�<؄B!�^_ʦ�0G�l۶-����ݻ-i�G�R��'�(��]6�N;ARF/�f�g��K����79d��e5��0N�* �{��U}=�$ЅH.��sb8����㏷iӦ�ܹs��]�A�L���=��Ç��!j~饗ֺ�����&�H��+������ʤs��_�&>�r��7�� [��k��.��~!p�և��2���/Ȁ���b�xg��o�\���k�ԢIeC���?� ���A��U` ƙ��+��"ل��ܧ�r��q�#2G���8D����{J;�����_�H��w�iFg%���I6o�ܼ���O�a`s�wد��?���>xߊſ_����0ˇ���ͮ��0���Ki����W1K^���;�d|�V��Q0Y��[g�>�`���׵kWo���̯N��Ǟ��*/��_?��$��:�d���T��g[w�So3�1�L� h\�0���A�q_� �
'�+}�(Dҩ�7�FǎMD]�h;4=j��9���3��8w�.�^��{��R��Fz�y������z��K�������(������v�\�i;.�� ��8�;s�ٳ��	Sz](���8���$)��	V�R}�lV���g� N�D�Z�BF��c��%Xb%D�/�c���D*��3٬y���6o6!Dip�1�x�<�3�&Tĵ;�����ӱ�L��8`t�Q��2w��;���!8�� I�c�dHr0Z!�.�� :u�h'�tr��L�6�.\hI�gU�u�>���K/��4��>�=���Б#G���� �D��B���q�F��<̡�4�W�j�?��w�^��`x��H�!ʞ�+_�q�>1��g̚�hq�׬�֭ۥ���_�"=�ʑ�v̘1#��g6Șo޼ٖ/_�#�fϞm����!�d8s+Zylݺ��8��S��~�O���WR�E�44V4$Ѕe�wmڶM��z��6O�p���ʭ�S�TP���:A��\��9b
7�`_9�˓&M�J�Y�R���ʅ�r��v��e��{���5��E%m���&�%���^���\n�^BQ��u� ���謷����H�رc��2B��|�z�q�7�l���r	sL, ��\�T��arp����3eЅH6�%�իW�B���+���c���������B@�7����:��X�<y��jpA��iǢ�e˖^E	��<���<ձ#i���@B!DI���7m�d۶m�Ԓ�Ĺ��?ڇ�(_$ЅBQP޾}��#���o߾��YuzqU.����@B!b`��m֥sk߶�կ_|��Rd͚5�Fi/Bì��)zs��ֿoLY�L���B�� �.�(+p;nݦ�}��?�{`����H�7�.ޫ����ի^��>���5|r��[o�e���e"Y���g��;�nGq��{��v���~�Cy�U���޶m[O�7iҤ��pjoݺ��	Q�0*�Y�f�������	!��z����SN9���,ę�*���8���;�^u�'v��/_���5�f�S(�����e���«Q�ƶ���]v���	j@ �r.�w~��b�T�~g�����<u�M|�2��:�>���\�e�\�.�@2��$ЅH.�%��Ν;׺�l��&�Ʒ�~���*�=o�����|��m&��5;m��_����&��/�	�1��~��
�!�($ЅB�"1s��
\�ٖ-[�SO�;<(V�B�		t!��0�%�}���7�xÄYӦMc/��ԧt.4T���k?�%杧�~����.n��J�$����t�x��o߾��ke �D�=j�PvdEmx�
���3!�Ȇ3ELŉ'�h�5�~fjA*o��N;�;��Tv��a{��5!�.��ܬ�ӦM�������߾z�p�E]< �?�V��!�"$Ѕ��X�n�����Dv֮]�}�nu�����.��;��>�r�/N>�doZPƻ`��P��]�v�^�zU_ްa��X�� ��>��98�������������#��5B��%��V�\Y�zp�",[�n�z�b����/�-E(iw}�dy�����}fl/����?�1,Yb7n��w�ׯ�L��iưqN-D���7߬���#8@`��`|7`���kfŋ���s����	"�"�pOգ.�H�%�W^yń"
�0y�׼����{ѭ[�������3-��z��x:����#Gz��4c
H�;j�}�]oƴk'�ׯ�u������o�Q���f���`?�߿�-_��3ܢ7�B�"z�>�h�zhȐ!�gLÆ����*�fΜi�'O��>��D� �.�B���{����=]v�Rxʾ4h�]F�B���ŋm�����]<V\��TSY�޽�q�N�:y=�{;�ɇ��o|���/�F �1x�`;묳l���v�-�؜9sL��B!�(9��]��a۶m����tB�xw���S�N���<�8�ymdΩ�A\e�iӦ�S'R�s�M�L>��;��N8ᄬ��eg���v�M7�s�=g���@BQ͝w�aGuT��?��_���$P��!^6!,|�]~��?���֪e��V�*��ڰaê�����3�-Z䍛��m�q��b޼y����2`Q���{A�{9��"2]B�ƍ�
�E@����F���z��y睊2��u���$x6���E2!sF�;V�x��~�z�j���B�j���c͛7}���淶o�>K,��X��}�,^��HS�*Jf�f��zn)�D�q�g۷o�6��s��5�6�y��g����ٶl�����a>�V2Żv�������y0��{������ċ.���u����Ӿ�9�c�=��Kw���������2Q�H��|YT�z����	!��T�d�9��ݻZ�0�>�,{�ڎ;L$�#�<���k�.�j�uǠ�@^�`eE��8G�3�����*�$���wPR��g�Q�=��g���n�-�d���~�7��?�x/�U��y� �^"�;|��Z�s��@BQ�P���Q���	�W_}51��;�O;��B@�/}�l�_��ܲeKY�z�]-�X?QXh�q̝;��-OWBP����=��#��'�>t�P����f�t�@B!DY@I�I��Lzǎk��"���mn�(<��Ӓ�KKM���"�gϞ�t�R���������X�j��҆c���ڞ���_|�N=�T�k����B!J��Ntc�
Jz�e4=̈��9������
Y>(x��n�\��LD�/[�,e�p)@U A  %�^������wN��b�*���B!JJ��B6�Գ���V� r�]�PZ����*I�D���ZP��*	t!�BQP()g+f�<�l����/���]$,]U�oaZrZ�jU���J	t!�B�,��"�[�n�m۶�Hr�A9��|!��j|X������Z�={vE�Qɂj�÷0����^�6�%}E����T!��R�V��d4�af�9cٔ)-,��#(!��=d1��s��ئc֬Y�z��#����
v��ǌc3g��	5]2j���/�O<��h��������H���(m$�KF�=��c&���W�.�m�j��axb���7�<����m옪�����ƌ��Jf���^9r&�{͖��S��|�h�sb\F}�@�-��d��m�>w�{��g���@��]�v���~d�G�eӦM�Ɩ	'�w/�����K�,I{��c�zU0y�d����B�����<N�CVדּ�I���O��V�7�ʗ���;vd�-����b�E�S�@2a�+d�q�g�9B�O�>�����#Gzb��I*�v���G��������kC�����7Q^H�!ʊbD��}�ⴿc��X�#ɋI!D�3p���U��7�qR���/��!`�i�&ϛ�r`f��1�#�I����;��Y�B��B�B�dEoX�$МU!DB 
���.����l�\��Ea�ԩ�u��1�m���oF ��۾}{�qo�3}���Xb,�Q"�^� ������~'L�`B!j��=a}�t�cz��/�5�:wln"(�ElQ������<(���S�\���s��da�������\��IIw�g4T���Cݖ�nL�����L��eǛ7��=����7ߴ-[��B	��(o�֭k]�I���B�d�f��y�;�܋+l����W}־���M�2阊B*i&��>7hР�2F�8�gk�AD4�Z�3N.��t�o�t&� �U��Jf̘�e�۶m�����HQh$�KH?���׺�2��'�B��ᣏ���xֺvin����D�@����*��0x�֭�wa_�~��:4�NI5/���$]*�͛gC��*�i�b���&��D]!�(?:W�A�S^�h�L��ׯ__-��L�G���[Ҡj�W�^YoG�õ�����эc{�r����{��\K�B	t!��#,���T"�D��7�|�DeB����3�t�͈ZW���,�8�ѣG�9�.[]̲�t���Ν�͓�6��w��6u�T+e��H6!���B��a���I��֭Ï�E���{_Expw���RpJ����S}����! �sD��Lz�1^)'���������X�re�=s��Lz&8��J����h?�B���`�B$	t!��#d����b���s���w.;�Dx����J��P~���ي	���Q�FU�:mٲ�'���3��&M�T_.�xԺB�y��9���k�Z�A��e80K=��j.f��W@ 1���*.!J	t!��#,~p\Nǁ�X�0�/��V�Z%�T��a��9��>*��zl'����i]:i�Z.$� -p0�=�Nv�qy��=~�+�_\�<�$���gcѢE)*Id���a\�`t������TT �]f�,y�`�"�H�!D!���ϟ���z�V*�x�V���/����F�	���9�={��!.Z��g2c�2�8��1�Z"�ƍ�	x�U�D�~ ��m��f���3A��l6�;�V���`_ +�~�2���}B��A�D�w��u}��5!D|��n׾}��'I�������c�L�废����/�W���/����q�D�s����]F�@�W�.z���!���5��JW��q&ie�a��q�ب�ˠ{�����[��|(���Iv����wI�BH��\�4�DQ����W�b¼��H6]�t�qy�ҥ�`��;��[2���v��٬Y�2����	�N&=[&�@}��}BȠg��������7o������;	e�����A:B��
�I�&G~�7n2!DraL}��̃>h�6����6m�T����z���ߧ�~(2d����K�-�����+^�9��A��^�f���M�;g3�C�*f���Ul�A*C���yҼ
��!�^�P*w��כ���ر�~x����>I�}��G���#�����;�j�/��s��n�Z�68�����W_�~�<����/������3RLW	��d�1�"�OfaNb˖-��O-Z��z�m۶Y�����4{��b
tLd��O�0�8���@B�:Bc��ŵ(/�v����9ǺTp���)�J�]���qM8�Nv<,��J0�_&�|J�5���L�ރBC5�spwB��}Iu!J	�
�u��֭[����B$����Mdgɒ%&�Cа+X��9��b~��8���Ϟ�]�vY��M����8Z%hs�����S���v�d��/����2/"�H����^v�e��'30q��P�q�=����!��_LR����}̈́��?��?v�/c�D��� q�9��A �� ��ā����l��s/e���>�т@f��w�ws���y�|h�`k���F�X�`�	!���BT0��N��ad)B	�H.A�DE�&��.XnLﶟ���b`x���R�Oe �|�	�0�C^�Ν;��@ݷ��*艎��W����
�Ȣ�#�}� �?PE���v'��ƠB$<DTش��&�H��)d��)�J
i	!���!{���={�Ly[zn�e.{舻�S5��2�-3��kd��k��n�ƍ�{"ԅl��u���;��qB8�L�Г�*�>������IZ
��J������@�"�d�A��뮳	&d<��Q�n�Ʉ�Q��1#i��\��'W�^m�t�`̘1Y����k�,�:t�P}g�;�+�y��>���	����'F��������tL�($|�l9�q�&�(]rVnnA�8+Ȋ��0���Ƅ(�,RQX��~{��k,J��
�$B�d3~��9<^}�5�)G�L��_�o��{��q&JJ�i��ӧ�W&��a�X���6I���8�Y�u�~��t�^s�-	�H5��O�3�T�#Sf/�@�8��q��l���	�p�s���d!D2�I��\�����?٦M�R���4���������?�|��"���7I!�(u�d�݈����r}:���e+�{��uUe%DB�ei	8���_!�P��~�ڵ�0/$P2o�<��-[fI�*��0NΛ�����}��6	!DzB	tN�<�M�:5�/7}S��~��>^��B!�R,s���y���"�.�	 �d]�t�.#֩R�]T�;���Ȏ������ƨ	Q�d�Du�cη��H���k�_}��5"78!?�쳵�_c���$��o�{��z��nzZ��2��V~/^:���k�ҥ^)�+�ޟ�lRQ�N����B�Y����:�<�&I��+�4�N���rK�e�_G����BQ�����6vLU��!�Ej�w�Z:�]��᠉b�}و-&���e	����VR�/�JȠ��ڵ�h�B���O�÷T�#5}��H�����z����F�J��%7BF!��o���Z!^
-Ѓft��.Z�(t��]Ʈ��?!�P�ɧ��ӕ���we�Tg!�K}f�>���<�q���n�Np�~%E���ц�B!J��lNd#�[�l��sG0ѦF��ͫ��
s�1��C)��L0�e�����"l5�16���f��"B$��Ȏ�����ID.���P����'?��	!�(m�L_m6��=ZYӣx��l3p����n&{�#P�6�/��Ll�8'����>;n��`8'�H.!ЅB�b���l����[����ԓ�؏�/ֶ͑&�3{���#R(w��C��O�V�����?��G�<_�+�`Npc��6l��]�*/��oT`H�Q�H�!�1��G�g�ٜ���ǿm�Z61J�S�K��6x�b��-\�Ы��ѣ�'��B92fv���j0'*�3ݘ�u��y�!�)�G��?�=�u!�
�+W�Q)P���,
�WB�3o[R�Oy.a��b��	!�(��x���;�~v��LDK*#��uq���ԝlz���~`DS�jݎ~t2�;w�-[�$�=O�xл��?)��H��}��J������#����@��?�r�� o�3�(6,¾�N�B!ʃ�7��;��r۶m���~�t�S'k�Β�tN�YN��J�Y�j��(�W��!��BhB!D�8�HUIE���L�H>P��(5��9�Y�fշG'ad�C��B!�H�!�E�3��;d�)	��q��G{[*�n��e��(h�V�䋿O]�<$ЅB�"��KF�� ���3&kk��py�fV:��2����O�{X���2�	��ڵ���"�H�!�1Ьi#������lm�;Ԇ�얨�uʔ)ַo_�s&8QB�|ٲe^�=.���j����5~������C�״iӼ�B���sqO��D�YIT%�0� i.�B!*�����6vL��±w�^�3g��E���e������)F��_vO� ��Ni>k-ͬB�q��!R�H�q�7on�$��!�B�d��h�T0���:#�
	��X+��Ax�l��X�tP!�~�
�3&9F�m��JT	Qd-q��
ԺF���J'I#߄B�rAҰaCO$�aM�ϔ�O�:�2��/�aϞ=)o���߆���]�ΝM�M�6y[*�Rp�q�U_^�`A�}
N;�4	t!J���/3'2���l!F1��<�� )�BDYD�q�w?�z��A?������J���K��l���I�N�n�B$�P&q|�)��o�Y�a�9)rrT_�B�J��W=bG�$���k2�.�xX'�8	~�8���������"�����n�e=��J�!�MhwN��5�J�8��}�ᇵ��d�ɖsp`+�)���������SԌ=���ͳo}�[�q�FB$��o�%��'wnH
�]��з=p����A^�����{x92n�8O�糶`���%�$���=|z�����3�� �m۶��ƨ��Ъq�1�Ԛ�ޭ[�}�=z���{��B���5�c�dG6�͹��t;9<��Þ8O��z�M�0��8�B$��3g�I��Gq��}��=!Ά(g+�)\���!��$�?v�Xۼy�'���S��_;���#�p;�����|��^2�*�`%k�?]�,�4��$e�rGO�3%E�;�M+�BD	B���ˌ#p��Hdlٲźt�R}YO2��H��.kn2��tS��8Sf�B��%ҹ�!�A��H.Il-8D�B$�w���ʖ-[f¬S�N��z4K��di�C��!T�I(�׬]�v�ZG0 �ҳgOoKf�s����@2y?�ر�F�"yH�W=�P��N8��!�H�	�:^!�0���i.u�`̔si�;��3YEf������+u�80d�gϞmÇ�(�y~��o�K��_�֤W����6l��˗{-�)�1"�i"���E�L�l$�+�'�x|�������B#��ӵkW�bɒ%�?�)G�����:'d��e��&Z��� b^W/.�]�&M��ݻ{υ�nDe��ׯ��#ϸ57rM?�;T[�^��FF�`ԋ/���NP�Θd2쯿�����($Ѕ��`�֯_?ّ0J6�k��۷W_�a���QlN�K6;N�,z��r�< �/7m�+�m&�[�.���j!Di"�^���������`�!�H&k֬��|�3՗�ؑ��pF�;"�]�6�����֣{������W�+O&d���>O�x����$�E.L�<�	 ju���@�P���[ߌ�~�V�����ǋT�Er�v�N�q�g��G�Dq��<��+V������Ʌ����c����.��md�ٲM�qcb�(��r�@���k��+�����3��e�]V�vO=��:���~�{��S�������Ϯ�L �[n�u�X�V�̬�����+���ω'ڐ!C�/���� �`���5��qL��e˖՗�;�<�2e�	!D�����t'�3�U;(	v&q��㞉.D!�2�Y�f֨Q#/�B���f��}��/�(-$ЅBQ80mv��8e�p��N�{�}�Bą&z�1��t����P����B�j���rkܸI��S"��L$�Ծ}���=#���.��y7Zˣ����[XÆ��.u0������0�-���L1?�a�3g#s��}�\[x���֭[��=�u�N�:y�z���A]!D5��rJ�Y�٘<y�WJ��?��u�o�b>N�~�]����O��?��:}���ꓭE��&�-=��sc� d�ɢ�A߽{w�8�|�.#*99~��4G��5�����~�k�.�R�`���ý�&W�>�h��mڴi�D!Dr�@O �H����>"!�������4Ϧ�Zg�<�k�L��(A���3��[]��Cg.��%<(�nѢ�'@��e���g���;v�o�a;w�,�jFd�#����̞=ۄ�E=b8�;��/�r?��Ÿ��E�)���)���ٰ�M�d���L����{�S;�ql���g��c�ԩ^�(���k���r��� ]�t�6�k۷o�Ɩ!֓����cǎ5�c���'�@Љ�&�Q���	N`���~p�5*!D2�@OC]��B��9�6��a�EP\ ��~�@�d�%��UUU�'���ܚ�������Q�.8@�Ά<3��f�۶m[����L8��A(a�z�V��aÆy�	�Y]��R��������.Ŷ�g!���4j��VdA���{�1�HG�?�Ìf��>h�9��ጐ$;� u����i�n�:�ܔ���?e�6�޽{[�=�q�����Q�� 4gΜ��<�!B�3��Lu �_B��(��hfs=���t0���v������¬P�t'gz���˴�q�ۦ3fq����Da��T���ӳ�������7QX'��k~舶b�!�=����7n�a��`��U�Voǹ� %瘺�:"���Y6���A�<>�<����2D:��d���%g��"�ݻ~|��H6��\ĳ�4܉q���$�_��۲q��燾�k���۲1z����y�y�e�'�^�z��O�]��r�ك��/1/�7`1A�K��U0���޽��5'���M�l˖-^�<jXcR�����;w�:�,���M�ꫯz����Qg�q�����_B��Q��|PL������M���<��6s��H�R�_��5�_��0ʵ(kɁ�n�B�РA}o�1��x�|��U&r�����)�=p@.v���{��T��3�~�����h7f�ϟ`#��tw�K�|�ln�^�Ҍ���ŋmŊ�HG��ʪ�� �P_�h�w_ł����^��o
BDG}ʪr�0ѓ*�y�}�E�g��I1j��Lℒ5��K��J��O��?���1�uaܸq��A��^8(?�cRSH�-g���33D~]�2<�"J�q<����^@F���TB��*�֬Y�eԋ��"����!���	C˖-k�g˵u@/�{��iB!�B�2��֧�Y�d����F��{7��L9Q��unD:I+F��"L�P�N�>���ϟ{ �D�cРA^%�%]%�!O@�ɥ���R����7��~���~��Z�����mĈiO�Q!"�]�vM[f?��O�n�(E!�"�`4���ls2Ք�#��d�����8��<'��ݵk�z�!jm��1c�x%�a3�Q�m�6�ӧ�W��7T)�:ܴ	��unCI;�sw{m q>o!D��:t��aÆ���m�K/��Q�����.d�3���^����B�L(1Ng6��r�xJx4~V�j�*wxߏ;�f�m� 	[V�8'_��<W���`O6�¹s�z�b>h�G�K���e�b)ywA������l���k�!'���%J�(�Y��8��������VD�������B!
ʵ7<a-Zd_��|5=����̨蘃!f�t��11�5����G�����#G�t���:���G��/4��.�`����СCC�-�J���11�m���^6?��v�)��Ô�Gϓ��R�|�"�E��sm߾�	�tzv��y;���-	p�x��L!�($k׿a[���],��-K5�#�S\�@�B��b��yP�S��|�r�،h�k~��1��N���(�,��d~&�Ѽy�POx&�d�:���g�߷���Y�f�&�����)�;���J@�>{�|zvof�;i���-^�����C�EQ!��׿��~���Ȣ�=��H!����}����u2�n|>�O�%r�5-����A�S��g��5�,n������qSϥ���q�gV��YFP���#�l\�3gN�*�`�;�* (��uD9�U���e�l�<����߆[�c�Y��w�G6��6e��CQ:�G}�.��"+&eL�0��BQ:�iEpSbܢE�Z��G��N𲛜�|~�8Tk[���"΃�։�t�I��5��`��K�z��:<Z�=����TT �y��w���k2�.+N�ĉt�#��eJ��8�F��U�j;��g+_+�V�E�����N=�T� 퇃l�
eaD9�r��`���j�٨�ʀUB!D�à8"k�꜏HC��U'k���DA&�X�����W��v�~�����s0`�͛7����l��tf���[�߇�˜o�})l���4�Ф��]��N����%��z��}F����Y&*��	t�g���J����k�Gaʈ#j.\h�Ǐ7!�B�ÆK�G�Qv���NןKOq�@N��p�$~H�`��j,Y���?�Í��̥̝*
�@'P@�&S��A�\J��$�y�$���g�]BK��AU�߭�Q&*��	tX�r����?��n����4�0���k�U��BQ��gN_����)S�k׮^f�%��c^��L�U���ϗ.]j]�t�����L�0��E���H+���.IPM�>���x���Ae�H.�e����	
��ST�����;��N,"�Ҥ�}�{���B!J��1�Je�E��&����A7|��i�,=WR���\>'�bMIf�`A��
Ȓ�^�Ʌpw��T8,Z�ȫ �c服������O�͘��D�Pt����o�ٌd�6lX���D}�5���C!�
�J�����jq\��;$�����,9�"�	���<^:u�T���dɒ���kC:�g#(���R�y�-û�7ǎL��
���Ç�v��C5	��M��
��{�~�﷋�ˎ����ښ��ɿ��XF�d����/z��;���K��g�y�n��V-Ȅ"_|��2�'�bI�q�ָqv��m�_�c���&�!ݧO�׹Qc��|���b�ɚ���Z���O� ЪU���ON0 MV:N�9昼Ĺ���t�|���0y��xc��}z���({��m��-��ӫ�o�U���&1�1y�9��g�a��ַҺ�������W���FB�����,4�����K�'O�$��.��c��ޮC�5)$d9,8����1�c����=����,+z��U+K�f���x�y�9w䂛S���U�����kF?SI}�L<�ЧN���c|]�Ϟ*?Μ��f��$���&��Iz�(\�PO���d��&*�D	t�����{��\r��y晵Fy�a���K/����)@����/u�S��{�,�I޽{wϘ,�q
F�4��b�H�ܘ��h�Z�P���.�@�I��0d��p�#�.�ٶm����#���o�0B/W�"9�@A��M�RyD�Q����`�� ��fp<&.H��N�(�<���{��I��\'�p��n��{lĈ�F���D*�N��pf�;w��޺~�zB���'�t?D;�'��Lz����eT0�DA�Z�=I.�/ƨ�Z����G�	u�߸�*�o߾i�]?6��c/b�`oZł�,a��<�u&+۹s�}�A��E"4�%C�	>��w=]=[;���]����~X��A�g϶O���?�q�"7�>��2!�������#���
tB����'f�D9���Ȕ�"8c5��R�h��.� ���.��nXXg[���-Ƃ�!��X�R��(� 
Y�ѣG�]݃x�dk���fٗ�����9$'T8p�m���<�Te!y�v9�,\����<�ٹ���J?��h˔�S*�z��Q����e��{rY��1�lժ�w9W>!D�$^�����Js�0�f�
u[*,n��f�v�J�X���?g��;i�$���M�|ݖ+��[<���Y��n���s{�����,�� �(����c"��i �('�lډc��(k��ɱ<g�
<^]c��EdQ�'ݺu�`�Z1�@����2K��f$UA1� �ݻw�ϑV�`�z0ۜ	��,��|���������L�B�F�P!*20a�0�΢ɇR�q�ƙ�N�@aX6o�m;��gS������v�w>mW]�i�@����pCa��f�3!�~o2�.�e�s�~�ڃ✪!�%�	q�kq��l�?��w���[�.�i4�P����@Ɍ3�2s����0LI�e泥O:� b�����%��ʨΑK6�}��E���|�o�V�FcքH6�BT�dqr-�ɇV'`ٲe����0���K=�jHU6%|b?������N?����8�v��ի3�s?��ŋ{~6�0-�)%���#�)��$
��3V˵Zp<� �~t���>�T�s�W��/��a�y���W;�S�����B�瘫.� �=�s! �u��P�g���0�B���F�9�C�/΃ '�;�Äy�={���1}|�zH�ǣ\�u��q��.A�0��rb�F߰{����ׅ����z>���j��	�!�s9F�����gA�<�A䯲U��%O�w�B�{���o�87n��)���A��E]$Nr�r���'�r��@6���ϧ�.��>����Aq�lF	���\�մ�_rp1�`�|"o��LVX���\\�!8[;�2�`R��:·�V����8��.�j��ʘ1'��Q�D���EO'�o���p���Qo�sq(Gܧ�A��%��|�.�-ǃ���s^e�D�m~اy܆χ�7�=�3,�T !Dv$�E"��.
*�E3������r2QΆ�,�.��Ҵ������@g��*���~U�G��'��ϕ�@�=��l2�a��[���	�ɮ��.���xX����y\k����w�Ź�υ�r6�"b���@:�#@�X�" 
F��C�\������r_��梀��@���^�2q��%7�H6�BT(,���tQw�3�Qy{%�"4��qy�[6J�7kdW|c��p ��pRm	���D�1!b�_��1/�2_D��.������:(��*��:Yr~����-"983�At.ؚJ�A�K䣄�o���5���61$H�} �Y��@u�m��Nߓ`Ձ"yH�Q�yw�l,5#[���w����O�훚���|uf�Hf���Ƭq,�ؖ�
q�L�5k���F���g���8D �_Ȓ�-v ��/XM�h��y��dr��U�g�e�*0���gks���}g_,d�"$Ѕ�bW����sg���B����x��8�����Z�<Oh�a�ڐ!Cj�+a��ɸc��ׯ�o��e~��8p=�~�D~���z�P����TUU�t?<��`Z���D ����>��@EF�6m�����iϞ=^p���q�G!��B�	�`�SO��}���& ��i'���cr�6�iӦy�ܠ��%�d^Î������{�Ddج�!�t����4�	>G׫��$_S�~f��G����Sû\����
�d��x��l�?{�&E���2�������� 	�ΜN1g=�g�p�����!f0爘83��3�� A�A��ͯ�֚������<#���t�z�o*���!���!^D���ɥ_�~�����ϫ�{L	��{��[�"b�]w��D���V��AH�ڰaô@'2�p�6�NqF0���	QO$�\���b�!�{6�K�ӯ'�%��zs�yP3�$p�rC���R����rԨQՄ0��Q���� .j�AZ��~p�p���� ��4	3h2y�~C�b=�ɤ��瞺K*�U�dH��5z�h���o�����N�:�m0x������3���<xpࠏP�ܹ����#Gָ�2�;�s���3F	نe`
5���vnV�^�v�m}��՗K� �AZ��Z̼��jŀ؝5k�~���ǆ�y�������OwyM{|vk��'�ܵ���.�jC�����Ĩ�+.B�$*�/��Ru�ᇇ~?�A���o�]80�g�~���+�P�5�}�y睧�}���u�a�.��B�B��q�E������R7�p�g�̝v�I���W�ű���y�%B��dh�������(A0���Z�<�4��LVŹ��0�ĥ�A��E�q@&%�u��k߾}��v�$A=�lI/p��$!K$���.��� d�L�������֯[n�Eu��-������ܱc���8���������i�^��%��_|Q5n�8��3Q�|���裏Vg�}��_B���6�5�D|��󎁱��,�v� �q�L��F#.M�;�f�%���e�����8�V��^��"W����	Y��/א@M�\[�k�8/�a=g�>�ϣ�p��T2(������E�Bvɔ@���Kt}�؋��#F��Q!-��k�Ճ�_��W���n�Z:��	�t�G}Tw�y���D��	�ĉ��m��m�Q��4AHD$����@L�>�C��fk���@�a��F]�	�!E�_�Yn]��kfn���%��IB�����v��Ejh���ݏm��&�R��h:(B�&u��!~���W�L�ΑG�YsL�K��9%M�K��u~��Ԑ!C�@L�8���V{�9眣'��z����_x�Oq�`|�}���c��I���SN��\��o�Y�H�>` ��	�zV��5�)wc����
5�>}�(A��`}jZ�n�8�w�uW�ɝ(j������	6A���uR�ӊx�)�D���~`�4i�$rG�B`�5����:t��Ax�h7�5�Cy�m��w�s�vGwAj�tvW|�z�Z(�j�*��~�?H�ҥK���te�����l~�a�vο�:�=z��5�n*��[o�u�m �9䐼T��Nդ�_u�Uy�ǀ ]�8 h$�a���Wm����7տ'���x�	*n�jA�$@�����/j�M�5/��n;N+�ɾ��F�d� �ZgW���{��3�ͅ �f�X�l����7�����)6͞��AN�,\�Բ��9hӦ���H���*��΀b�44��H!Y2����O�uW��Mf4�s�[ٵk�j��@-8k�^v�ey���g��t3�T�/)�� ����j��A��A��>��7�|Se&���̈́	� � $i��@�1�#���ڑKއ�oР�v�!��Q�F�0�qA�c`?H��kx�pľ��n���o[6~�`l7��y!Ni�K� ���'v�� }��َһp�D죦�h��{������=�����p!��,M�ԁWp
ћ���PydB����Y�Ć��@*��I��ѽ{wu�T�z�y��WZ�^�
��Q;�
t �%�.� ���^������u�A�Q�O��-#�Y2,��Gv�1�5�B�g?���n��X@��I��#��y�1��L)B��r��oD&b���w�9��n�/���Ms8s�8֨�������R^�
8����A(?�tı�!|�1�xֈ{u@�c�=<�ׯ��k��N�~���{�6g���]�6�K�Ξ��0�-� Ba�n�E�Y�Ĺ�L"��;w��"8i�n��$j���%c�"��7��:۷������=�L��� ��t,/��5�A�(s1۱����.��c82�~��K(! ��%/B�H}4��9K�~�T�޽����$^�����\�΀��f[Ҩ\Ђң�m���;�:��<G�.�~��W�^�{�|뭷J��Fl���O?�����վ�7���$ �c8��]AH�)\�e�\1OD>i�mDup�췩�Nc��<�C�G�IM;/w��b!Z�#��漅@���//(m?8OdX�9��[��@��P9d&���GQ��~���IʗA�E¼��1#��ⰵDt�t!5G@TOrm����o�޻�Kzơ�� �l)U�s�4�xcuZ������w�|G�5�Q�h��3��"J"5���h;�]�m�R��ĵSD��b�����$`v���@GPS6@�?B��������k��ū�#7*Է�j�_�>�жmۢ"���~���qK'M_�$�4�]i�c帙�.I;	AH�L
�SO=U�Q�͠o��h%�D�U��~��6�L�~��{E�Br �1���d��T>͉��KN	�s�黩m�m\�}���oV�IF��to2�#&�b���m����dD.��UD��~"�ԛ��m�4�٭��ڳo�'ׁ�,6v"��6B�t��ŵ�sI:/9��G��ؙ��&_s�q^���Zf��O����sA�\ʲ���3"��mG���%5l���D̄���Ck��6��C��&�4&VA!���j��M��.T[��3����c5~�h��A���D���D9m'�����I�Pc�L1���T�B<�w#f���=^Q]�-J�@��X�"/m�+ha��m�������[kԨQ�"�,����ӫ~&;��x��t�9Ŷ���
���wf�:q�	Be��@�9��g���;�s�9G�+�0Ȝp�	:������sn���}^�ua^�`���˂�D�<��ɔ)SB�7J��PX/�P�[إc����r��.Vs�P9L�6Mn#�'�n9,f�IK� ���A��D��ԕ��4�Kc��`�W=8A�4�w���F�� ���d2s��B�ߤPf5y�d}o�����6���loj�;��m2��΄s��w�3�<SG�mX����y���V
��7M4lq��~���罇��Ͼ��k�ߏ��k��;�pp?�������NSB�!r���C��#t�+x�`��J�{���}�>]&�N�Y��6I�:T]�n��gl9�SPZ;�;Ｓ��A nq8h�w~�Ro^��)���v�������˹��� d�Lt�?���6Æ��[oy�)��[n�%p`fP����������U^ 4
	���:�3��;A���[Cf��֯�E��&����@d0�6o�\�0]�����4[��Mll��
S6g�pӅ<��v/�N��D���,Eϱ����2�p���n1M�8vĿ���l��$�{l��w���s�P��&��g�lD|˖-u�eU� d��t&XR�]\^�g�yF�x�y�Gx_x���[o��~<�w�q���z衼���\g�G�#������Rخ���j�g�}�'� B��g�}�!�Ml�q�n�p�����͞]����y�j���J��*i�t�nذ�.AC�9D��5���d��5�M�$���b_UDt�_l �� d���w9�L$R̹3B���k�;���,KS42+5
�<w�ر���={���6`�E�iR74�ZR͎�s��Y"�Kd;HQA�,2!�8�w����������w�qռ�={���t��o�>�g��ÇW���)Eh?���y�Ǩz��t��O?�WFZ��?^����G��?Y��C��{W�Hky+A�H�_o!�;�@2e�z�����6��IZ��zaU��DX��N�(���t�����E��H��P�6�����-R�N��j��ܸ�?I4&�W�n��ҢE%Be��@'%ͮ��+K'M{�M��}�V��LW^y��ѣG����ٗ_~���bA�#̽R�h�ƒn^�i���S'�|r����'�|Ro�����ҍկ��)�'���`Aj��	���Z����wT�kQB�ǿ�ڎ�Kc��0%w:Qd�r	A��=&JMVL�6mB�Ax�h̘1UN �)�A`[e�
�P��.Щj۶m���~�W<�����WG}܎�������n���>Z}��G�<u<���P��+&��;,T�w!���ڑ	�K�.�20^`��;������Ӑ���?8W_z�ķ3��J���_^���rX6<�/�AZ>k���܌��(�5���&zt���J[����s�Y�J���n�tJ�3v�qG߀�A�� �J&R�]0���~饗���I��I4;J��!E�H|D�<�@u�7��/�8RzԀt�=���~�i�Y&1{�a�*��U��K�y��ف�5�� �ܕ�d =#����4K�0��r�h��u��R��.4�-T�'d��qW����)͈`R�I�6�Ҁ�e^��;��H7��b�& �$�z^���2�.�;z�Ң�6,�ÁF�ƫ��%̒�����:8z�XN��Rɤ��h�'T.q6�L�:c0	3�ѐ��1�|
u�tt�O�>�.P]�v���N�B����ޫ���:�C�+����֭��~�Q�g��;Ｃ�¶��W�~΃}.�Y/IO� ��1wȐ!J(?�tm������*M����9�ȑ#S]��98�S[ �8Hj^'jM��W�%��NhժU���l�^R�L��؁I-�����gdwq�^Ď*�aI7**�D�I'��Ҁ��k��/<�4��s��FD��O�^R��u#q���o2Qu��lC)uGt"�k�s�y(u��t�P��W$�X0��P�����ϝ;wV�{�����2���������+���vvu�;(�f��\�8�A������X�AR�M��1�D�a��� a�-Gj=6U�.���m�]�w!�γI���(��EY�f��Uf,���	��N-�-7���#P�&}���*�e�lP��X�ک�!�6�_.�yeI��'By9��s�5�,�������gv����t��hؠ�j�|3�ݶ��l����J��paA��'5�D�"׆(8"��4��L�8� o8���a�� �KLP�=e�ű_�q��@@������l�Y��|��B��&x���dϋ�s1��dp��(���������f.�97i�f���,�_W]uI�M��U��ᇟ���MQ��VB��	t����n�uGd4hР�簓�~�.]B�W&��C��B���R���)�Y���5YHY�V���n9V�޹�����U�4�D9�z�6���4�.i�v�Ӆ��l�zr�'kn¤��كv7w2]��!�d7�ddH?��	Ĺ}mh6��s�f	�P������sXm�UԹ��V-WS���� T>"�k8�H'=�����f���n�ܗBu�*�A"�%9��}����6�$�ܫt��a�d�oZ���x�9m�fo�f��M6M����hXp��nn2���\��8\��B�ԣ��`_2�ԝ�Y�=I����k��q	gϤI�B}� �|���f�A�0;��D5k❩�%?��"�k"�Aj1[�����꽽z�RS�NUiA]�����ʀ�o֤&[˫�9"�h9��r���,��}l�8��Y����ei
t))�d�P���D���{��߾}��N:zU$�����8�q���nU?㌰;�������t�� ����7LD� T���&mi@$0�@����o��҂(��ʁ{�k��=MO�B��i����}������7}BR�bG�Ӫ?�����4K@!��EOj91����Q�馛&�9���]֕mu��!�Һ\K��{R���QF���^��܂� ��⫥�}���:�e���#�����[n��{����O)A!���z4'*���US��5�����v�8"k��ֿ���Qϼ�0�_ޏ����I�� X��j��<K��QsM� �h^8]8�$KL8�'N��	@x�N�"9X%(��sS� ^k�s��5b��w�����B�9f��fŏj�5�C�F�߀P("�A�*��c�؛�!F�~�钾����N;M�Ͱa��{ｧ���?��~����@p B���"*h�������:#Ĉz	��A��k�#)�H"�:L�=	���9`�iF��S�³ۤI��8�e
��4�=P�@������.�`Z��j�2)������gd���l�����ԥ��VY%�y�����3�P{�.d&�Gy$�{_}�Uշo_%d�]�����������Z�x@�߹`��X�)�Ŀ<ܒ%�S�B� �h���,�e:�ч�7/ޏ�D����_>N�"���g"��dʔ):�܈@��QNPh5�M���>p-�,���K޲v� �(|Z��۫���w����q�M��Zv!;�@}��;�������?�wG/P���~�)��J�"Ѕ�����>��z�~��l��Ð"l�� ��
[\Q6��f�/^vgw��&U!֨Q#�"{"��:���$aɴ(ZD ����=gB4ACܒ����ڵSC�M�AZ�p�q{]o�!:v��+<�����^�{9?��u������M>�����c�P��E��Q��+x�jC}�WGY/p%z#1��oFmmb�����_��j<�`�Bjٲe�+��/�H:�pl&���_8���p6 ��D��L��֦,
�a�����݁�6M��8q�����ħ�Ԝ}s� �i�?N'�-Z�T~��r
��j�Y	p���w�?M�@g�Ȱ�RIs���TM�	�?��O������ �C�ƍUmc���F��2�M,i�ʭ����Q)fɳR����J��'r̒]�QBs2�@ҽ��A��I�8����EFC؀����r�`g��LJ�ܹs��#H�F����2A��\;�.d�J���w!s0��v�m��;j�(%d��~XpAP?Z*��Ν3G�Ԝ>��#��9r���WY�#�R�w���ﾫ�z�Y�� �| qf�� �8:ޱc�j�h�-�Y�"���t�����o��.8fH��b�-"?�K�D�M�=�AҬY�j����	�^%ddg��]D������bB� �5��Q������$m]4n�0�]�Dڸ�Q'�ĭ�;�K�⡖���I�6�e�b���,Qd"ۤ�S��m۶-*�q>f̘�9 ��Y��{8��8�u�mHoO�� ��@g@;�E��D
-ua#� � Ɲ/�n���Z%`�8�ˀ��Y�:-���~�v���:�@$�-�h^G���[nY��M7�T�H;+��%=;��>��,?�����.kܸ�^v/jJ;�Ĝ��.'����N;K	�@�{u���ܔk�>A��ZƫݣG%���^�z�z/�`�AA��m�F�5Ĉo]��KM5���i�-;��c �lCğ�n�^�����3:��9 ��6t:����vە���4v^aJ�'Z�lY���*ӦM�D}=!��jڴ��1G�sSSN�#j��O�<x��j��I�'� ����� H�� �  m���JD���,="ӝ:uҢ��A��战4�Q`��O�9�"�Q�_�
�A"�8G~�&M����NV����a�� �>�����
%��'"�4�+&[�h3�,�Ã^d�9�H�G��Py�@��0Y���l�߻|�7JA�ab��o߾��{'D���r1�ԓ���v:2��^p\�(Ёsij�	g�!iڈ^�5��8c8'Ժ�o�e���rV*6Z� ǃ_����K���tD��R�?�MÆc��C=4����#�L�.�ӟ
�DU�#� � =�cǎ�QR����R��rI��}~�[���(�2e��Ҙ�:ug���7�5��81�-��a�Z�sw9����@�5���Ȓq� �>j�@g�f�f���J�)@��ׯ/�+ ��=���w�u�����[aA�,:���c�6ѓY�f�����L���C܍7Y7�4�8�kh����oTq���h�%��,sEM��:�s���\"�;�C^�E���I�>�a���T�h���q,�I6W��w����Ym�Fƈ�x����9q{/�U�!Bq���Ǔ��4)�sJݙL��0�~����	B��:�֫��w���>��������������	�<L��-zK5h��*�O�qf�G�"@L�pR�M�7��������!u9M�
(��+m�~Fj�j7��9"c�&h4(:�bj����z:;�n���gG�Y���d����ؽ�ya>'By��Y�	�_�~ړ~���ə�x�M��6�s<��px�i&4��{�N�� �H�|����[w�L�s�p\�`���W����B��&��)g�s7R���������.�^��
�eݰ�2(�B�6`�v5�+==(�����_�i�F�L�p֚�	��)Љ�<��S�W^ѓ/]6�=�1!v��Ew�qzy*^�_~�G;DC�lC��!��Nl���m�:ut�h�#'�K��:�Wk)B�`�  M�1Q��w�]�,��%�6�püϘ�v����j�4���ID�k4@D��=:P�c߶hѢ�܈�D�Bv�8�Nt�gϞzpe�!M�Զ�_~9��00���G�hbu�e�i�N�P�kt
��DڡC%��8∲n?��s���*!s&�ĩ(�&��G���~"�mG!vC��ी��NM�Nڬ��P��#{}y��t��Ӻ�i��g�w�"ݯl�y��|�LP)� �d�N􉨵i�¤㵤I����#�hc�eV������[oia~��W�z�#F�	4	×�e��?>ۭT��Pc�6g�����oR��\
����jպ��ߧO�&�B�a�=���tu��a!�U��d���N�i���mf5"�~K�	����(G�3�ז�Bf)A "�H7��y�lٲ�����	��=J�4a"�ݫW/������sO7�^xA�r������W^y��O:�$��K/隰�����5�
L�A��ڮ�����Q�F����t�'MV�P[i޼��G)ufDɜ3�k�/Kk�a�P����}�>�ƍ��D;Y����9�� �+;�SU�z��۵k�E�Wf�-��
p	��y�s�]v��VE�G���ץ@:����I��v�w� ����;u�˸�6,<Ǉ~�A���Δ�!L�:Sc����L<j�Ӏ  Ml	j� ��>��ǉ������Be�}C�'v���(D��)��kvI�/��� d�<�N�5�(��dX���%-���n�A{��@�v�a�m�tӌ
�NAA��w��v�u�~MI��!����"����8�Q.��t��I�;� �g؊��=�#�Y/���N��đnN:8��8��5�4�����>P_��;*AA�g�pMT��W�;w֑t����8��Z*�L��X0A3�x�f�|?#Y��m2-�I���M�yڝ�������e���w�މg����3gN���}�ݪ{��J�.�u�α~<X�|�ɱo�%�&L����}���g9tI.Q'Y��4��D��f�;��:uR~��~ٵ�[o�u�*-��+�pH���Hz�������X� ���
t�Ԩ��#^.aL:]����[׮]��<����
��-��e��w3Fâ�ե�\�*�w��_� x3}�t��N�r^��m�喺+:Qv���29)jԤ>\/��:�x����@A�%[�-[�ԓ��F^L=��<�6�˽V#)pD�hRw�A������6m�T����E)� %A�-�qb�i�oD�d�!�Ӡu��U�d��-\�0��pVӼ�|�����j'��N�&2J��MTx�%��vA�>%��?^��5j�H���￯'"��i��{��mȐ!j�}�-黨�;�쳫~/� � ���ŋuI"��~ V&M���i@gm�vLf^X��~�bw  "�����~K��Ί����B�!���.B�d2�}РAZ�ge�p��D��~���P&���B��!U(󤶯g+B< DH�eI)�F�s� @��9��AN��C������~B^��9����u��%��xp 0�M�VU�.$�رc�P3`A�8�i��(?�c޼y��-AGkl�M�E�n���q<"�Aj6��L���5�@'�AM� � �5k*k��7߼*"�*"�o	9A�f�9�βfPh���1���?� � D�F��A���	t:�BR�.)u����� فN�]t��l�͔���޽{��S�*AA!�dK� ����ԟ۰_�Z&�����U�&M����G��5k�;\� � �&s�&.n�UV@�G�)Br4m�T�y�ׯ�:t�^{�5%Bya��R֡D��9�t[�"YX�]�?Ȫ3/kd�dHj+d�}��GJA�Ȝ�V�n]�Via���6� �0@}��ת�ByP׮]� � �PydN���I1��:t�k���W� d�nݺ�iӦ��
KBJ� � Be�9�n:1���O�Zj���馛*AA�0L�4�*�l�2%� AdN���O?��c�:�ҐJA��,Z�H	� BX2'з�b�����N���Z*+|����I܎;�A��:�(ժU���3f����Uh�r��=/X��gϛ�P����o�~�S�N��XA���6�A(��	tD0K����P�B�fj��-Z�P묳��2�a���^{������jf&�SN9����~��������~�~�={�jk����|��u���p�|��g:��湂 ��;_��� K�:�瞺3���k�]������=��C	� B2D]~��U?�F�}'���b�-�Tm���2 &O�\��d�y5�%��o�Q�ƍSK�.U� dk-[����f�2e��b)Y����WM�8�*�cǎ:�\
�o��jܸ��;w���r�?��X�^�X:���^{��g�u^G  Z~IDATRX/��b%� 6̭cƌQ;Ｓ���#�8B7#:��r!��M�V��,\�Pm��U���{�A��:u��� b�UWՑslv�,���YJ�d�>~�x��{�U���V[�,��c�Qݻw�⸜Qt"?���:��cu
Z��>�ȑ#�~nР�J��?I�r=�t����^z�J�!�v�e%T��8��mڴ��O�)�a�J��ڵk�'�A�<�O>���R�d�;t��I���1F�J&M�Diذ�������2c�%�PӘ>}�:��3�=�ܣ3�����r�m���8��>K� !���r�Q	����]w��	B)dV�ù瞫.��Bݡx�6H=՝z/&���?_&DA�,<X����ꫯV��g���Ml�c�1ԩ���qml�/����{�b�B��qFﬧ�zJ��T2-�7�tS-�o��V-��ׯ��H�����裏V�Z�R5<�{�{��[���8��������A�i�؅H���G������w^s�5ڰ6<���������_~YgSԞzq���-�w�7�Xj�0�mXr��
��.�@�;V	��[�Hq�Y�&�l�V_}u%d2�<�@��̻��v[Um�;�P�_��=���w��nj�m���?|�p�!#�,�/�q�	B\�	t��Q=?I7���;��ftD��I�|�r]�N������L}T��R�P��7�{�V��z뭧{(���8�����a��N�^Щ��^ݺu}�3��������e���A(DS_}�U%T8R�@���O�?�ߌ@g���*��qn�x@	��p��ĊU���'Ї��7o�x�M�N8��z�W��E'�$R��n"�l�m۶�[�n������\!)p���~�~�7߬�����3�8]����� $]�?��c���[�����ү_?5z�h9�9J'��.�L�����/����Qz�G�Ν;W}߼y� �b���J�������WEc���i�g�u��p>���A@��K�
�x�IQ�{��y睧����t������A� YJ��t\,X����@�ǽ_�Zゐ$d ^q���i w�W��N:I�1��LA��⅍����c�!Dى�� 5��:��t%�4�в^�-�ܢ'0�KW�R:��bN�8�l?���� ��>W��QAj./����+칟�&^^��@l���Z�&� d�L7��u�ֺ�Ͷ���S�h�C*��i"�g����r<҈t��O?���:\AA�R�W�%�\�z��YUsD>v� �P�8�k���:�s�a����y]�H��FX������p&I�9���?�c;v�5^�� � B��x�ҹ�]���N;Mww�'�|����+���� �P�H�n�x���G�f+&LPS�L�MW�&2�+��~{�tTI�A�J�Wϣ�ᇴT�д��Պo��j�js�r߳K�N�[�;�)\��ʳg��Zn^�v>�|�ک�M����V����J��U/�6�������Z�������i���멟~YG����9��U6~U+���Ze�oU�U���MU�w���0���=ե�J�#�V��.���9���y����8�A5r����ԩ���=�ڒ��j���Y�)�����N>�}I�j��M��ςW�i�d#5��J�N������P�}O=x�ڽs����Q5iu]���Gs��'�R����SO�-�d�/V��X_��|��tH���;�N�_W�J��SV�G�R�P*-�Ԣw��E����E��Z-��Dʉ��^s�5� � By�U������}*QsA�ZH��.Ԣ7j�H	Bh�Ǫ�e3>�쳼�5�Y�dI�{Y)�����d���|���>��.�t���;�`���qr	� � ��.5R�B1�{��U�3�8#�w^s�5�U�8 �wR�Q��k׮]�����RAAA(� �P�3o���w��>U�׭��?��:h��c���?��}j�zm�4���?���6R�u��:kľ�)�-P�<4\�����&�3N�Euj�U�ۡ�����!�>R,�����٧�V_=~3i�3�C��T�>�Zm�x#���;���8��,�r���;~�Zc�:�vP'��Zy�«݄��eߩ;��F���V[mUu�>۩�N�VYee7��9M�,s\-�5T;gw�Ֆ��&��`�R}޸���[CuXkuğ[Ǿ��zv����d��?�6��P��Em��ڱokƇ����ꃏ>S6��N=��ڳK�ط��?�{����':wj��?��Z��j�ok��9��G�U����sr�Q�7�};˖�W���?Vu�p�����ժ����Az-�t�nݺ���s��Q� B�|8�su�1�i�d<�Cu�E{����mQq����5I?�5����\�"�fK'��6��4`��ꎛ�,�I��?���9�5v�ܪߍɉZ�z��OՍ����%�x�����l45{��ST�v[ŶD��Gݫ�6�Xj�<�����&p�{o?&Բ�aq��M�2_��~O���m�#~���2w��S_,��t�ʴ�Jn��r�5/�5I�0����i��s�`��O̝�#OzP;o�@7��a?��:����;�gV�n��y���8��g��u�Ķ-���\�v c���:A;��b����a�=��pF�=[=��X�]�`#��B��#� �P����^�熛���o;����ߜ����w�;�R����X����U��Ĺ�_~UW��em���x�w�Ĺ��ȓ�ԙ���v/�F��߯Vk����?�nW�SC^� ��3��mqnx�I��wT��ټ�m����<qn@8���T��8�x�bu�m����&�="=.�>�87��л��wP�KXi�f؈Y���/X�n�9@���X�ý����Ĺ����_W�j� g��ύ���Pw?8L]r���lg�7�]w#�������7/�-������sC�����V��$��&��/�z�Fm�v�m7U�aM���~;�{�C� $K.F��Xo��9c���w�q`���E�=��7߬�$�q�f����*n��'V
��0b��0A]y龱l#܏g_�����Ē�I�r�'_z�G�+oLU'��FO?�L}��@G�".�0�p׎�K��!��[�@G�}a���9oq	t�_���8	XʬTX��Ȳ�aS\��g���v�5���Z�����%0���_���ЋΏ����&�����]^,��k���%og�3�8c�t!)b�8�����m�٦�t���=i.�v�I'�:�����K[_TJ�W���U�4�,�e<Ϫh���oU%�l�2�bŊ���&�6���ӎa?ƌ���ꫯ�7+�WkX�l�j�9zFn[_y��]���b�x�?��,h��3j��ف�?��<���
�w�D���3}�H��.�Q|;͝��-�;�M�������	t�I��~̚�����S�Ǩ1�E(vKж�g�_��s��Ĩ�~��_�x�cw���>7y�<���漹��L�6_-^�D�1f�G�~��,_~�:��믫m�A�>~4�3պ�U?s���;vsO}n�D���C��}���k�c÷�z;��Υ_��]�n���>Gd|�L�4'�s&���|>�vܱyᢥj����1���r^�lK
!)�;L	� ����2i����8w�45�y1)'v�=-�w�s�1�4��>�*�sD�f}�H��ǋ/�W�v�CX|���P��Qcf����w?�ܨ1��ے/�	��9s?��܂�_t�<��ؼ��y�|j[���P���#̸Y��<t�j޴A���M_j;3>\�wL�&�	�܇3��i�.��󥁟�h梼m f��?g�w�7��eS,��˂���+W�W�߃>7୩y���0�m�O�5��?7uڼj��t���Z�di�����k�� {�	��˪~~F�{a��ٹ���|rO}n��Yy���?��΂���>��^�$�Q���1j�FV�<{n��hػ��gU?��a�熍� �o,�<{���3s֧y����?7?��W�OV�[N����T�#Y�"�k(x3y�٤�T\/� $�:묣�[o=U[Y}�hi�mڴQPi��*�n]���K.Qi��V[�J��ͯ�WX>������e�g,���K�꫊�o�>���G~T�12]��p����b8�h�;���_Qy���
��9ڹ�I�+,�t�UE�T��������WT�{�~��Ͽ.ꞛ;oI�����S���k���~����1�"=��������r��WT^|y�~E��#oW���t�95j��P�N��o��i;[l��*'��M�0A�Ya��膇 De���J�l����?�,��N;)AA��D,!�K��{�n���[�{W�{ｧ.��2%By�+�:N��v2kY?Y<W� � �l$Ž3s�Lu��w*YD�����`�~���s�9'3Bx��j��Ѻ	�믿�<�@�8W� � i"]��e�������Wg��:�5�7�|3/����j�}�Q���kĳ�t��<�<��;Y?g�u�j޼�5�K���N�'�xB	� � ��tA*��w�u��h�����i |ǌSm����~[���;n�5zc)AA���tA*�ɓ�wlAA��!]��: �K-_��,ۧ�w�u�ͫ��B����wHMu�c��V+�����믕�]X�%���Wj�UW]U�oŎSB�0�s=L�G���K��ra�M�k7[�6�y�[�n��Ra\k����<p?���jE퇹�m�q�.]����3��F("Ѕ��C��/���w뭷�
�X�B-Z�H�7N�&Sk`)�����o��V//dl?��3�I�&U?w��M2Dׅ^�ڷo���v[�T�]�}���Z��SO�'�|R׳������SOU�;w��ov�ɚ�~#G�T����z���:���y��1��������[���U?}��j֬YU?�͚5��;ǰd������4kd/^�X��NS�w���a8q]�L���������"]�}7��7޸�oӧOW'�t��gIw�����{�Ua��_��N?����q]�ߘ�itƱqo��A���cնm[��&�h�
������{���W��~t��I�y�y�c��`�\o��t�#¯��/N&üy���^Ծ�w�q��|��j�ԩ�Y�4iR��y�}�Q��v�U�����/�7�P���U��G���g�}�U{~Vc4h�� �������.\X�9ל�b`�4���g���K�������e˖ꡇ���g�Ơ܏��o������nj��7����8ó����}�F�%�x�l븟���NӦMӵ�<�A�����yu���={�g�Õ���Ξ=[��A�y^O�a���]�vUs<��s��o��,�k׮z���5l�P;�9��|��q�-���ۅ�q��k|}�wԌ3�!h|e�:�S?�<t�%�膎�l��>.��fn��65lذj�a|����!ǀӋ���Y���o^ :x6��<���&���{�9���rD����0��}l���F?��k����7s?1wr����b���W�_}��<'��<3.������,�{�y�W��^!�������|2ql��.E���K/�sd�x�g�%f/��u��'W���ɽo�k�����?�-�u�\0f06���+����v�7����1��ls^����믿�:���8ٱcG�馛���[O���9�9��/����Y�]3Ot��Eߋ<[Ks/2Oq��<g����~�=���|~��z\�y�X��l�ͪ�
�i���
<_�í}������_���e��x� '}~X�c�����.T$�4�raPjܸ�~u�Qz ������̙��V�ZU����O1�3��� a�vЃ�^Wa^��1��=��*��!��㏫����s��LR���<���n�����\��iӦy﵍hѢ�jݺ�*���z�����D���7�`�l����+!q�����&�0�ɾ��L�L�.�38v����x�E�4�︢A|w�k��̵�3B]X��]G��Q��)���<׽{����9O�{�wh'�12�i�~������ 3���G2��Q�0��k�3��2め��=�.T�=��~�?��t���X��h?����?�8��ׅ�ϲ�8ƣ���߰���j'�� �AX��.��b�	���8-.��"��Ѕ�1��H>�3<��s���O�*�\�_y���%��N,/���
��G�q��q�ת뮻.��<�a������?��ꎁ�8�� z��;�B�}u�{�ˠe�(A�g��F��w���9m����mp��=�����w�8���ް�j���|ÿ68Mq���xn@<;6�x��3	Qn@���Z��n��&=�{߾�K�bn� [�ˋ{���ϯvp��=����{�ˁ<�8�x�Lv�ay�L�~v׍1��"s$���`�c@��L{ݻg�}���`�fۼ�7���g���kႣ��!�e��B��@*�#��F<��@�W�(���7�|s��O8�_���l�>�^n��D\�Ν�EFF��	�h/�6 �a�-���-}<�� ���`"�#�C"	p
`l�ae�f�.<�x�97nF@%�x�k���`cB'��b�	�CCgN��������?m ������\c�!��n�cǎ��5�\���B�"ƍa���v���]~ 0�Pb�!/�/8��L{g1���θe;%1�lq�=��%���"�9;�g Q�$���i���`��+TVa�=���A��6(jd[�#8x�>��#��1��`�oŤ��\0V�\`��%&����9"�̿�r�v"����_��y�駋���^�z����`��N������,la23���x"��b�Ȩqr �p���\l#�[����/�8�Ɇ-Bf��#����?�����p�]w�:���q����\2q�Ī��m��m�1� �|��2�p�o�����L�N7��j�e4Qh��a���V4p��6d>0Y�@�s�.��R�10�a�C�9���[\��^��,�>�i/��ľî�؍w��x&����u�NNn�E�9��BqA-���V��S�e�ź<��?7���B���J��]'C*'�B0�䍡�dI��L|L�n���0�A��D(1N�Z#xR��x�(��-Ι������I�Ў�/0�2�X0��<#5�uv��I��%,��hR�0$0܈0���&?(&�+�8�`!�L���9�Kc�����d�ͱ �86���؈``�r��( �
ƉuL��7�R��r+�/#�Ah&s�"`��~������{q6�=nxf��`pp?"��(b�]��+cs|�X�<w6D�2�4�d�Dp���ꪼ� 2�v�.�h����-�Ə�)�M��5��,�k��ۆ"�C�%]!�u�XyM�6�&��.# �s��*"Φ���#��l�@$��_�8��~�3�Mv@����y$Rǘ�<`G�p�"����G׀q�B��=�p��#ɸ1��A�/Ay�H��ϲ8 ��W�!7��gڌ��S7���9��x��@1������5Z��8�8v��GF�s>�/��q�y�g�̊��=#`��5��P(�u�<C�%DZ��3w�n�h����f&K��/� � �ñ�d/p���Ic7"�q�{��Ɯc;'d$�}�(�m�e�8A���S��!�H�)�yv�: ��䭷��i��K�Is/qo1�e�q~��P���d/G�'M�9�u�36brL*:�����a`�u:c/6��	^0�2��U�-��a�5�s�O�
lG�&P��2�0���,��}�5161s����ݻw�ך�A�kF)����}�Xm:u~}�{1������Pфx�Љ�L���^���2J:'k�܋B�)9����ͽM���^ܙ���	�ŭ�2 
Ic�87��<D�����!�z��m���n�m!�x�0pb`��go�c����c����A3�#
łw��&����:/�F&� /���L���Ƥ��75^��ӭ�����baܺ�8@����1���LM*cF�0���Z63�کv���б�㏲�)Cz$�<F���DoH[��A��!��j�^��c�8�����Xγi��wSf�<F����u��|�=>�׊q���&`����yLݠ1�1j������&��:��d�`�Ï��Z�"������1�6��('�kTgz�$	�<{_hD��p��Ӄ1LA;ͷ�3Ͻl@4!��{�Py��}<�8��L��&�9`ײ{���ᖲ �8R�f��i���!�책�krv6�-�-F<��<���!D���g��<��ݝ��g�qD0�ѷ�c��g� i��k��`��3V�w�6|����a���P�/�^���-�����	�7���3Y��~�����J���ۊ��+p.�ӌC��9{�k�˸���̳�v(_2=p�q�]��8D�m�1���1�y����w���`����G�@�qc�Q�1�����c��f`csS�#p�ٙ,^v�WD���bt�A�>,\��s/�I'�/#u���y�|�{q����[We�,	t�Yt�O�D�P%��<�;��E�z�4�:@�&����yf0q�	7��u�[�� ��6F���"�Ů8wa�m��E&m�'b�׻X8^�i�0`Ȇ�^p-01�["�Nq��B<2�a�0�s~��N����];L<��T��� {��&	��cֈ?"Bv��2����#)��B��k8�܉� �ϝ����6@:~׊�q`�)�$�X��`�u���A�}�q�"����`��'q���S��(�9GƏ_�-)�8�l¸��![L7�(�?��jG�q��<D��iFƹ�#��/p!p1��9��ܫn�k1� ��u��(���ט�c��D�:�z/�! *l��Գ�i�gt?�c(��_&�n�D�����'�mg�M������s<Hp��os�p|�ı��̻v�*͘�:5��t��A��R��87�/�v�0s��Lv�-�C����a�]�P̽HA��{��ʜW�E���d�ؐ�Z�L8و�r�'r�Mѡ��g�W�&�ܽ��F��K��� Y�ss/F��N�3��$ݡ[�\����7\�͔P#@�! ��Hgr7�3�>��n�IK7Q\&>kғ�\lA�����2�b a`�Ej�� M��[R�l�>���f�x���s���}>�s�]F#O�Q�$!���l�P��q�{I"J8/l�c�#M~�Ѹ�M��!E�!�=����4�����0B=0��^~��h������k���Y�1j.���Cq�L�����9�Wt���8纗R��#+���$�O�{=�'�B�-IFp�&otR�Iۥ^�T8e��Tl�Ydg!jLd�("~"�d\0��5�<�qt�}��϶('�h��%*7Nt#�?�4�D�ӄ���J���u�Ǚ�}`j�Sm'ύת�۹���-;sW#�k
X
\{�
�l�'�d�p�ص�d߸㰻�~McA*8� ����dzv&&mv���r��v$����ch� D�+���6�o;ӤP���A�s���ۯ���=K��}5�����܋�����@9:O#Vg�N��7����_��O���܋\���P��!���0� 2�5�ň1��)�@���L2�ۀA�t^F"sԗ��.�6������&�l�+F��ί����x�upp<��b:6�!�芒fY*�'�5l��H�cҴ�y�y�{�1��I�F�-��kCڛ1<0.1���h+]��dZ������B$�TJ��v-4�H��m�q�K��Z�䚷���D"&��&?xv�+�#��$׏枲Ũ�;=E�p�)�q�s�@���5���7�Tz]nc>R���*&zn0�+�!��, ����Y��d:�u��m'P��f���-\�i����D��8��>�X�����~`�v��Sܮ���z9�ߙ�D�0�uW'�9"��ˡ��WvL���c�0s2�D8�8����@�0&j�[~K�{��0[��y&s�r	:�1�Pfg�p1.�Yn7��P�w�INR���;��]�#r�r�i���*���\�̝��T��IN�q��O:í귦B�בȲ�x������n�v�9\XhXC�,��z,��k40��ua��@ېFEM��ZMt8�u���;k1��^�~�Q���J��m�6�t�0^�(�)`�����i&s���I�� ��m�?�+c��	ᷮj�Pl7�3���#�#��5��Z:�k�� H�F ����H�U][|��G�tK��=�S�jq� �E$�̽���3kGeqz���q��b�8�&�u�s;ۆd� z�eDR�+)D�L��L�W�C�	]
Ac�Dmq`�{��.7J{�r�?R��d.x	T΁_3.{��~����ĉ���e��)��5�ǹ�Q�'� ȴ4�X�/l�0�P�1�/�����X��8}K̜�5���-�$(9@�'���L'�#s����(E����9��t" ��^�x�(�@�5zl��㵊#���빓OkhB��Hmz�Z�xG��`t"lL#�x&HjOm��a�1�(:R��F��-@�UP::�&��@��������10� �^��r]h�ը`��P��?P:uƅ-j��G��+�:AҴ��-��T�m�&Lbq�(�F��Ƞ礱Q�]J�T���f7�[����Y��8!�������+��KQۉ#����-[�	�?�}�v�#9W�)�Na�0g�mq�~9���L
wq�G/#�(Qe��uK���čN�56Q���g��X� Pr��E䍒-�
�T,�W�{��:jz�6��ˬ��<k�;Ϲ5�a�2�r�H=�9t�Z+��vɄ8=�n���4�r#���^+h�c^R=�n�}�^f�Eܹc�[�f���J�!��d���8I��J��^܋��G�e��{�1�`4�#hcCD���V�!���R0S>e�˱����L�0p��Ix��^�N@c�es�"i
t�P����t�];|�������s�x�xB�������`jM�0I��	c�^�٤�]7Ig2��4�.�z�Oj��4`��N�#��^���>�����>�}�h5�6�Jq�Wn�0��*�6�]��"��8[�`v�b���;�z�@2q�bmwS�a�G�h�`����`���L ��}��"�&���PJwp�)N�D������,j���O�=��- �gH��8?\a<ktNO!�NG�����Y#���t۩���sXdEm�TD���}����2Y� ����a�Bd/���q�)��&�c��2'�m����Wc���q��<sl��m�������S�j�O �������FcD:MI�#��id��p�6�����&s�^Y|��k�y��L
�7S�mlf�S�]\��ǌ�b��������[���b���N�w�?��[�cV7���c�q�-��ݬO���kR�9�)�$�5�^��c�i�<��҄q���j�xR�M��s�SR����=TF���]�s�`ƍ���:i
tZ4�;�*C���܉?\����fvM<!x:m��'P?j2"nZa1��QC*���&�@F蒂k�e�]2L1d�"��¤`��AT�0�Xg�%� ��oi�F!�l8�c���Q�.��0bm#������8��;8?^��x׃� �@3%D�J�7���:��2"�:<R��z	���k���6���c6M]��a c�f�}J�[>�A��0� Q��'�k�Κ�Rh���Rrc�E�QJp\�ORM�p*����_\�G[4sn��;��`��6���C5L�H���Dn9�ꨐ�E�U��ōt��̽n��	�w�?���|���^`���g2NC��NΣ�ZY̛F8!p�hHg��h�D�<�m��c�����k�H�N�8�9g�1"�8��pv����y�v���m��%l�_�m's���$�|��O��x�]�	;�^�ͼ�{�θ@��q�$c��v�&� ��M~Yn�xBe��>��.����*��cr���&��P�N<�
��^tm�t����h�߀M����b �3j�&J{��q#�gj̼�Ew��DK�f�����L,{R-R�p8����ذ0q�*���S�8{]��p܈""��2t|_\�|���[��}���Ǒ�N�����Kj�]��A��emS�ԦF����&8�0N���Rja�H7�ߎ(!���k�Ltܮ%�pD��C����
ҽ���0���Sb�DY6��?��lÌ� ��4�c�2�8���&8 �w��'��c�{��%�o7#cq��r����޸KRpH��N�yc��-{<��಍w�20�2'1��5Υ��{���j7
�*-��A�
��t��!��]�g�{�8o|���Ku�!�Q&�~8�2��l���%a0eCo���A7���>�\�Cc�HN1�'<�v�*��p<����1�o;�qF؂��7���6P���N�����ΠĮ-X��-�#��I�����a�b�3תԠ�?�4��ћg�O�'�#Lv� {�o8=UXRԫ6����Z��]����,�s�rs�)��e��IC�3�"Η��H�z�{uTBf����fҤI:�O,�"�	�b�&hi"ۮ����h^ͥ�(9*�=�I�A�ҭc�t1��<c4�ҏpi0b�Q�xH�,&����J��m�fY����m�t�g��J�&�5�14M��� �m���j��DT1f0�x�	�.�+�	��)�/���&?&w�$7���-��id^$�&e�ԇr��"��=i/��8�p� ����M�#h8��y�Qt�!�#߈-D,ƣ�8sr�x�1C�"��>/6�o��E������v�r	�1����^F0c�1�I��3 ��n�3e!2w����w�=� �$��"B�+c!��g��\��&�Ƅ8-�2nw�ÍRc��ںݠE��a\��7 �l.����t_R�����&�I��;�<+^�+E����>����a���3F��.`.@�b�l�K��P�Fܯ~s��q֞�ql����bĩ�;;�se/]�f1n�ktS�[H��0�r���9š`��pԺY8<���s�83khc�������}dΘfad�p?c1O�u�<WQW{��y��d��'�j�D2���2	�8$�=cJ�#�>�6��i�4s�_�wz����N�fcN�k�I��)C�FqW"�����q�����4.a3����v�Fj��R���L?�D8�x�qLp�px.�����?����@n�������a��c��9��ғ�+�G��� r����"��w�*!��L�WPA5@0L^�a��vR�� 5�K����ƀn��e"sk4�����q����K��X&�ΫL NL,^FKa�x��kG½�h�bA׆��\l]F�_U�I<�n��t]�j4�Gв5�1`���0��&g��GH%4�����QJ�?��&����`��40t��`�0ϥY���:-�Rz53�?".0ȍ�x�ܦ|�8LLm"��1u˦ֆ{��~+�8gA�NM>����ƃ<�\�R�_0��kܻ��uډ|�uaǡf;�l��=K3<#��L����Q�)U�����O=P(�����_q����9���t��R��e�pzu����q��-��6d���b
�v�d�������s��ӔPP�`w��6��o`{��8��,3gq^�-�X�~vr���j�V
��G�F{<��M�Qds�H!'�kJ;�`d�6B����	d���!)�	��p���)^�SP�Þ�>���o	�B+�}�]��ˮp{�ظٕl�9�P/��v�E�P��wU!��3�{�u�Is��"I�N���r� r��I�ĳ^k�����(�P����I1j �w��S̀AP�i�x!�"����I#ڎ8�Af�q���D���F�m�����,D��D{��(l@ qވ�1�;UȪ�����F���e�+kX�Ǹ_�*M-g��b��0k�,a �SL�h����G�&����QQ�U��#ֽ����{�1�I)�M�6���jþ�u�<O����GM(�l���/8F�.��3��5Z�N���l���@�g?	���0(�g���1�̎��}E��6��ތ�j�פ��c��q#���[�u�p�a��-��U���vO��iD�q'��%v����,2	�m��m��m���̇I�v�6NQ7+�A�$`�8Fq���������=�CG�]���A�G�d�q�4p&�g�q#�r38��.d�a��N�a�::�5�c�܋z�*!���]�*��}�''�N���J�		"=�H�Z&E&+4�Fغf�c�({��"�	b��+�}^�/L6�l�oY҈��=@ �h`pdBa�c��^��c�yK�5PnD��f�z�n�}f��Q9ƃk@sMp6���n�5���E�\�(8�i�5�x����t��'dUD���ɉ��\qΨ�
cP�����6�^��d�/����)� ������"�mGc���c;"�q���"�{��5�_;��<���|&�@j�m$��ٽ xf����G��dR�Q�!j
,���~�;�*>Ə0�ǆя8ǩHd��Ӂ��vJ���ٳ�~!+�ke90D�W��W$s���Srý��=�9CL�dI$/p8�%Ŏ�<#A���e��Gz��ky�[y����g����s�ߺ�6�cQ�kw��N�ϻ�8��y�R8��+
q�s���3��e��o��h��\�С$�4K���XG~{����'�������������n ۏ���M��|�O�� '>��{��{�~�s���E�]`;߱���Kn�Qn�����`�+��!S'�:���g����L�y���8�#��ƌŪ����O9����ʛ�HJ�3�]����t�[�����I�@��0��7S)QX&���0(�t3�c^�kwc:���R#�L@4��㨥�랍
}1]pÂ؏��1�Ô��/�~�]���W�q�q%J7�H)�j��Q��#���܈�����u�6=,a��(�/�u�v��0��Lq���=d)��yġ���8�����)�7���;�Fij�\���+,�(�5?p.
����Qʽ�̈́�.v:��ġ[h���Ӊ��
%��s"����$�?)�>>����wf��S�9�g)AAA�T�\�*�Kr�.*��ג���]�jW���ܷR� � � B)L���_G�
'w_���J4X��>5��CT���܉'�c+%� � � �&z���\֠�<�/�[��%�EU��{�~�W��*� � � ���o��1~���E+��M2-��S��^��(=]1vR� � � B1��i�h�Hf�>�Z�pK|� n�>+w�K[,9��&W� � � BtXZ�Fr����[���q�I�f�|�ud�UG	� � � Q��{�Q5��+��k�eR�S���������v�xYo����+���6X�����b���Rk���J�/��R�e�����Zw�uU�|��7z�ؤ�_��Ze��2�<a��(k�Fe�5�Tu��UI��W_���9���p-���lY_9)x&x6��k��H
�%I�~b�`�H�%Xg�uT�:���#�+����9/i�.]��yN��A��_}�4�u�yIQ�^=��j��$�	}?�o��G�`b&AZ������/_��ļ�=��Y~���%�/��bX�{MV5��ʹ,��0S�@� �n���p�#�.T�|�I�߽�����*���]'N�]�c0���Z$��ŋ�|��$ӤIՠA���k�$�p\�h��;wn�ߍ��8Ҙ칟&L���B��j�J?I��4s�L}M�Q�Fj�7֢*Ip�|���j֬Y�7�oӦMS�K�,Q�'O��8A�s?�5>͞=[K�l��f���#A�q̘1#��F�7k�,�k�5�2eJ�
1ղeK�L$����'x�ㆱi��7O�q�ӊ�>}z�"g�v�m��\1mڴ��O�o��>���%�������l(�FS�̀���8�W��.9�q�Y��́8�b�-�~�TZ�h��?N�΀ܺu�D�A�����6m�$>��F�m�V�7.V���mܸqj���͛����v�)�l��~���t^�!i'��=sq>��s�H��6ܿ�HG��%v�g�E\"=Mqn�g��8E:�!��\�喿�$��s�$3�lpܷk�N�;66�n�9�ܤ�=����*N��8ǩ�d��/�)��\ߤ�$������D$:�8�d�M��{m�k@� e����H�[�},�fq
��r��AM?��È�S���tz��v1X'M�T�H7�aZF��S�q�6q�t#ΓN���n\"݈s":qGQ����)ҍ8O�8E��I�S�0��%�����8E��i�Hǐ'c�T(��~Z}��S�+p
�%�mq�&��q�t#�9�4�S�q�&-�4p���T�n��4a�\HQ�c�V5���ޮ�	��F��Pӏ��(�8����]�`A��Q.qn�`-U����%��%�q��r�sw�������%��%�q��r�sC"�\���H/�87p?C)"݈�y9�C��K�����8D�-��A"�\���~�"�N�Fy�h�-��%�^��<����*�r�s``3S1"����P�H/�87�*��-����r�sºX�^nqn(U��[�J���RDz�Ź��t��b���[�J���RDz�Ź�T�^nqn(E��[�J����~�(�9Ie�N�44�˝�L
��qʋD�3@Ĺ�X��qn(F�gE���Y�bDzVĹ���qn(V�gE���Y�bDzVĹ���QEzVĹ���qn����?F���g���k�mlg���^�X۵cl㔦$-iӢ��6	�U�CQS��B���*�)�����"hR�&@��@ڦ���6����^�6�����wwz��:�̾y3sߛsߏt�fwg���޽�{ﻷI�"�J��nEΕz$݊�+�H�9WR�t)d�17��,ѥ3:T�H~��%9Wj�tkr��"���\�UҭɹR��[�s�I�&�J���8��Y�s�I�&�J-�nMΕZ%ݚ�+�H�59Wj�tkr��*���\�EҭɹR��[�s%%IOL~n�&�R����p�R��=<���2,ʹWҭʹG�UZ�ɹWҗ-[FK�,!�đt�r�đt�r���%�V�\�#�V�\�#�V�\�+�V�\�#�V�\�#�V�\�+�V�\�#�V�\�#�V�\IA��a���,�A�V ����`:e�,'*�X�s���[�s%J�UV�ʹRMҭ˹%���\��t�r�T�t�r�DI�u9W�$ݺ�+�$ݺ�+Q�n]Ε(I�.�J5I�.�J��[�s%Jҭ˹���Oᐌh3e�.
ؘ��;�D��IgK�~.������gr��'�^�\�$�^�\OҽȹRIҽȹRIҽȹ2��{�s���{�s���{�se<I�"�J%I�"���.R��ɋ�+�I�9W*I�9W*I�9W��k8�l��cv��i	O&l����8�(c�+v�A<<ɹR.���\)�t�wOr��K�79WJ%ݛ�+��.x�s�\ҽɹR*���\)�t���$�J�����Z���Q*���\���xG�FFF\ɹR.���\)�tIG��\)�t�!eB/r�$(�)�\������~j����W8�C�C���@jx�sE%]2}9or�H�W*���M��t)�h���t)�tww��sE�\�J�����K�[OOyE$]
�]]]��\QI��=�g��Jz___^t�ɔ"�.�����\QI��N��=�t�����$��{C�	iA��J�T�Je�G��n�.W�\Y��������&O�_�l
�-��{#�W9W���-�� �I�,�g!T��y)""Y�, �x�8,EDd����,<cE�%<#�����UjKI���Jz?]�p!�*��:��;�S�(��*.�M1!���lr���Zc
     @V���1�]j^>��e�uAk)K��Ĝ����s�\�(#��H��r       P�����=A��
c��T�OX��7���:s+����       �<V������r'(��@SW�^o���0l䝝�'>H_�fR|��cT��       P2 ��Th��7s,��RA�1�L<ب�.��D����yO       �׷��t�r����h>`��Kw���)�#���<��b������       Hc��\VE�e�&�u�#�,ӇyCG�qAVr<���Ԉ�%�	�v���3	�;9�N��;��)��z�`�w��Ү��d����mb.�;[�O�ˣv�,Y4g��]�����L��۝cz��Q�rAtz�xi�8l{���hj�X�w~�7����W��9Ñ�9t���i#�L�8F�D~gpx_��i������j���V��{9�[�y^G�N����Y>�O����m<�GH^a���銩����u����MO��G�wn�DO'/L�7O�MO��v�����˵��}����!��]��sl
��[�-"�m���� ��r�d�_��r˯�~��֛��w~������q�6�+D��eY�gr&������6�q�@^��~h�iA_��!�PEF�F&�����8�uA_ǂ>�c$�;R`�{oϟ=\�Zln�0-��m���فV�v� uU�̝lZ��ͺ\�Z�r`�iA�4�zz�J7����K�3�ZeI�yA�v-vi�-�Վa,G�}E� �xote��=����[7�O�F	��3��W�Y���P��(�8eٽ�%}�|�8�
       ��'�{�������9��Y;\.�Oq�C�&[������49�O���        	d��ؽ^`I�C�}�)��m��̡�'�2'ox/�ti�����u�����Q^|��       �;,�x��:v��d�G���亶+/TzI៩Ђ��� �#w�A��(��]�T�        Y��x�]��� �ٽ���	o��7+	�#wp��X'����Z������%ߡ        ��g9�c'�v��d�W^<����{��^���S�ο���Ia]�������m�OF���$/����        ���P��v����x_���s|�~z���Ȕ4R0�d��k9fް��o�]����?HM��A���ǧ8�       �f���E��;����;���>^<�q*�f7ǣ򡢠�	��;��?^���e���s��m|���cJ��2*t��v'�      �w2��#�k2.ڟ�+^�)6�n⸕�'�͎r<��zY~�j���
5�؉���'�y^ޖ��}��)����?F�p        �^ן帎��>�����(oKo�BK~;��L3���ø��'�y��]����9�7s����"/���=z#��i����&*��$��?0��X�D�N#ӌ��1�qZ��h�����4q�Ә�k����.��>A��jz"��1��d��W;�j�@��d��'=��OO1�Oc�&J�8�ݘ����1�?=Y�'�XeY��F�&_��0���y� ����%�����C^�~���ӥ�~W{��KORA��di1>�'�5^�=ǿh3=�×����
��ˠw��� ^�==�9|��z�����%�8I�흞Ϝ�0)���s�;/Ϝh�Dz���B��>?�kχg.]�����ԫItBM��G���3�sYHO��I��g�~�!.h��/������'�od��y���_O���fe 28�=���t>��(�l�ҡ���q/o� /�r<ñ����x��ߕ�3��(���6��        xEj7�EO|��Y�����+�cq�4�µ�=�e�DM�>!S��_>pz����y��XN�!��(���o��=��!90�����WP���w�1       ���*��9d��3��Ex���t�o+���Kc�����/��?Q�˪�.����>L�A�Rs��]        @�E�l�$�ೕ�k�u��X�e��         �p��Av�}��KЋ|�C^�_M         ��z��4����؂�+9������{�	         q���;Q_��]$��Y���?~���9�?H�Pgg'����oxx�����3������J޹|�2M�4�<��c��T�0�_�pog%=�t�ޟQYHO###4qbMEJsHZ�4���|��|�p_�:u�N�>M 8~��7��Ts���υ+���y�Ɓs��%z��i�ƍn%��ٳ�u�VZ�r%͛7�<"�+��B�'O��k׺������+}$=M��s������Eoo/-\��<"�=���j>�[��&L�4�j|<H���6Ќ3�#����glOO-Y��<""�m۶|A~���n����{��a�L���gwuu���iN����^{�.^�HW_}�[9<~�8�ܹ����*�=�YS:7���-[���ժU�ݻw��Vғ��<"r.��<oA�q��ϛ�վXW��+�<��dr3FX (�%�̙3y9!�_�&�*��Ν��,a����o�eJ���M�U�ED$��I�ʹ���g��.r����?�5�(�*�����o��M�U�O�<��Y��%]�|׮]y9���M�5��W�
�$]���ѣ��E=J�������ǣ�Xo��r>00����K^��ח���ɛ�C΃#��|~?Η�ͤ]���\ �(�r.h�/x��r9N�8�N�K�\!�&�r�x��r94��$�r.�5�&�r�x��r9�ǒ'I/�sA���$]�\�C��7I/�s��$�T�}�z��R9W:�_z�t��u�y�z�t�ypNq<�����C�9od��7���8>J������˹�I�+ɹ�I���\�$��\�"��\�$��r�x��Jr�x��Jr�x��r9W<Iz%9W�Hz%9W<Iz��+�$���+�$�\�O�9�tk�ߟ]�?5������.��/e�w�9
p�IO��%�IO��%�uI��sŃ��'�I��sź�Gɹ�A�ǓsŃ�Gɹb]ң�\� ��ɹ"�a�'�Jz��+$}<9W<H:�<8�����n��$���2�m]@`,Kz59W,Kz9W,Kz59W,Kz9W�Jz9W,K�.�gϞ�߳,�q�\�*�q�\�,���\�,�q�\�*�q�\�,���\��Ǫ�ǑsŲ�W�sŲ�C΃���3|�g=�,�����?�s�$ cQ��ʹbQ�k�sŢ�ǕsŢ��"�5I�E���W��fZ�"�ȹbM�k�sŢ�ǕsE�˒��f͚E�E�k�^��+%=��+%�9W,Jz\9W,J:�<(��n��ߟG�]IМ�w�\X� �G�k9lX��$�V9W,Iz=r�X��Z�\�$��ȹbE��sŒ��*�J�I�G�+�^��+�$�V9WJ�'7[��sŊ��#�%I�U�K�^��+"�r�W��fS��+�$r�	��9�6tB��Z�C�������+��a�d�^��+$�9W,Hz�r�X��F�\i��7"�I�W��ވ�+͖�F�\� ��ʹbA��s�ْވ�+$�^9W,Hz#r��}%4S��sł�C΃!2��cߛυXa"9V��万����!��0% Ah��7*�J3%=��+���6�ʹ�LI!�J�$=��+���6�ʹ�LI!�J�$=��+͔�F�\i����s�Y�BΕfJz�r�4S�Cȹ�LIoTΕfJ:�<�~��g|o�Zi���-�[,�7��Tx7ӱ� �JzZ��s�TҧL�BiR���+VPZ��sE%]2ʴ)�JzGG���r�Cȹ��5k�PZ��s�T��"��+*�i䥰(��r�4C�CɹR*�i�.	)�J�ܹs)-v��Aǎ��RIO�Z��s�T����R���4+�CɹR*�i]�y$���q+ߗB�<���w�^<�	O�K�����)=�L�|i�I�6[�o��V09WT�-ZT��ۖ�DC#�.���y���ɘC"b#¼t�Ҡ��JH�W*D�B#��Fzd2��
� �@�F�K�_�#4Z��ۛV%��_�O!�\I��顡�`�������GI��G�ȶ��'4�SE�OI_IG���H��ɳ)��t�ȑ��=�J�<g[[[)I$��sJ��tIOI��~IO!+{)Ƚ�Օ�$RR�#�%�QI��l����ŋ�k9�銳��.�'_Jj#����y�O�����;9��-��<�4��߹s'yF��;RJ�0�&Rh�r� $!	i"������L�W�g�#�J�4���$*��D*}B��h"UIT���H���{F$M{�xF�9d/�f ��==ei��.��8��e���M5��i^<͢./����a�e6�       �nE�e���c�d�:��t�$�Y�e��[8��Eү��       $��$n*�����U��-��t�Jm��    IEND�B`�PK
     ��d[�����"  �"  /   images/53dea2ad-2eb7-451c-84a6-1b4fef66a2aa.png�PNG

   IHDR   d   7   ���   	pHYs  P�  P���Dm   tEXtSoftware www.inkscape.org��<  "pIDATx���y��U��w�{kJ���2UBI !�DA"�Jd��->�x*v�zK]�G���(�����2=��L �		�TU�JU���y�o��w�͗�M���֩���θ��9_L��+5�W��5G4�(����e֬Y���&���RZZj�g̘a����e���2g��:u�����Hy�AY�`�L�8�ʎ;&��s�9GƎ+�x\>l�K�,���+������r��Jn^�h����K�.���l-���2�����;O23�dpp�����om��ӵlP���csg�h4j�w�ޭm2m.�HTzz��^nn�,\�P�G�����7N�ϟo}���[�)S�HQQ�����ظ�=��q�����_i�s�|[��ͺJ�� �	F�1a�1c�Xx�XXɬ�l�S�Z=RQ��Sh�Y0i޼y2~�x�q�+�a,�z�@���@�!MK"��ŋ+���l(�����ٸCq��r��u>�A�H�,[���g�V/-.˗/���?''����͑��?_222$;{��5//W.����-�YY�V�H��u��6��q���0�4wh^�ȟ�|S,� 2k�]��!�h��Ha�X���%S
��92a���˼	ݒ�5$�+�����d��.�Ȯ#AY��-��)]})�ɲ2ڮ��!�m19X�i���ʧ���PC�m�P�e)%ʥ�ڥ�:Kꆲ�3 �guȎC��8r��䳋:ek�rNN�jж�������dDe�y�,�
D�d��9]��4G;V�� �O���7��w�ebn�O��AQ6��Wf��-�y�_(=��_5�i^��7���� �n��͚�I<7�-��5/	) ��7*������D�o0�T��֮���2�5uƴ^@�^������ֵ���j���?bm�,�IMkz�����ֲ�����BY��,�+�g�2AE�����o "5:n��As�m�%J�2��О.i^���K�!�5wiި�� d��r�[���G����$��:�|i�[�Uy^.ӦM��h����`��;Xnb��=���w���#2{�,9�:���z����c2w�\�l�1���*55��6�8ioo���F����ri--&����V˴^CC��1�YiM�Dӆ���Z9k@�2SJj2$�KU�QC�4Յ�E�ޑ#�U�d��)S���E����$Bt�$�W�ieD��r�.S��7��G#c��[��1�d����	F8�yn,�f�k���>��!uuu���ۍu#
��"E�¦(M�켌z�nkkS�5����ߔ�d�e�_6���@�2�eMM���!�������̥������˨G�C�����{ƟX]ce�G?<#��GOOOr<tW���ѣ&j}��-�&� #�7J�%�5Y����VF�CHk֬�ɓ'KGG����UV�Ze� Q ```@e|�TWW�$���.��@HXO^x�!�	�J�-2�����I�&Y�|�)}�0.ϔ1(�� ���\������A" ���!��7s����&�qS�  �{�����ߖ�+W�a\<�����e�]fk���\7j~D����I�OwK`�"��k�O	̍*!> �۹s�Mj0,�Hʜ
��ar��Ƃ $�c2��ȑ#f��t��2�ji�����Y�����7�'��(q�5sչ���ː��/c�y��qP���q*��Oo��:���3S1�ܦM�nEEE���jY�b����R�|�4�^s��F��!P�W�u:���L��
۷o��3eήd8��x�y��7�>�#C5P�@��:~�������p�|�W�Y+�Xc ,F���Ha�!��ӧ�5��HΘ,��Ҏ�"J }:^�X{z��6����+=�u�$ѥ����1ي �'��I��ի�c�b��Ա�y��Ek�_�D����3f���
���?6?�#e�	��C�i�o���}��GM����ʰ>J���/���۸��;�AE�����7��"9����p�O�[�t�\��+�y�����wݩH��}�{�$�.bq ���A~�ؘ������Ųt�4y�߶�u�_&ͪI�n���޸B^���5C}����?m��CG��l_������4�c�{���d���!�Z>K��@��v����Ȗm�r�Wj��2sz��9Y���۴ϕ�g����������{[+����Lfj�Jԉ���?6j$�%�s�=&b ����M,̜9S~������G��&s��G�'D��wݭm��&�QJ�ʯ�_v��u"5�Tt��%tx�������,�}�.,6N����Xd��=*��&���ϕ���R~4OV_|��4E��[6WJFd��OwTT���k��õJ�铤���RV���Jsg@�\8K�VFd����{��4��sR��}Α���[���5Wɡ}��}KYe��_����,+�!b�u��OJ�=v�%��ۏ�裏Ј�;�cJ�ӟ��a��_V�8 /���YF���Ɔz�U t�	n�K�n8�O�K��3S��ʄ��f���~e����}�����O��.��⠽�û����uލ�=���$��=	`"*r�z �y!=H�"��$�cP�"=���Fl��,Dy"���S�����-]�0�"LsLe�Ͽ�zx���G���:a���z	�7|\��immI*g�h�o��v.&�/��GB� �caڟ��C�yb{����3k�-��w�}��)���@�m�f��e �o|�V��q@O���$bS�'��S�k<��To�����C��M
�瞓/}�Kf����@☄^�nD�y���Q=��w1�aEbQ�j3��wl#���N3Y�.���@F����{fـ0��[o���r�k&e�@��{v�R|4)6|�,��yHߵh6��ON���|��&"`�c���φ����7�h����ȸ�~�/��3�! ��'HÄf.�f>�"R"C�B�;v���b���$wn�'i��L楗^2�v�ڵ��� �I���!��#����Sp�#�����r��9�%��O�ؒb�b�*����`����ȑ�!㤫���l~2�""��  Y����(u@\򤓉6'�A_n��;iw*.9U�.�z�	�|�<O�x�(y�q�7ʖ-[N@��Z[Z�M4A���:��T),��|2�7����(0��f������;ԏQ��tu�����7������%Ͼ�S-���7s[�bE@ڎ��!I�S���snIe�p�W�g֍�{6\�8�H��b�' ������N	+'�`ee�Y6tx:�6�������֜�C�u�2$��Y2�S���x������Y1ɻl����͔%�L5����������N����l�}(���l�aY҇��F�wR2�S)1!懄>��C�h��;s$��ݻ��S�?l���g�Z�H}�|[,Y�Rٻ���d�6�ʴ�C*͎��<5i�U��7���y�ޛ�`�&�2��D���@�H��	�aU(n�!�0Q�D\��[��l����w�+W^y���]w�e�qx'��P�٦��xA����ʖw�J���7�"l�|���Y5�ӓ�R�ψʄA����C�y������1\<:W����b�t��[�\����l��C�J���|g<�C-�9�ǽ��+���j�!N"�sVu���Ǩ���=�|O(��UY{�W_s��^u�������;,+�Н��e�ª�ќ3g�\�z�4V&�Iy��/��֓Ň#���y����!��I������APD��r��>����5����o���f`�Hxd�.����c�=&�<�ƫ���@�QW�R�u�� ������G�(�w��Gy��-���o}��ҧ�xB���ԔdKK�E @<2��k�Qjk�l�K�_�{A��X�Es�X�����"X���J��,J�p�ъF�<��~��%A��g,���k��`g#��<g͞=���m.? Jc�@�G-	0ʭ���$�p�"s��0�_� ��hl��Y3gK_o��< ��כܣ�@��nQ�l�Al F���l�ٛ�Қ:�d�x��a�A 2�|
�1X�w$?$�:�ebD�;� -�d�B/�����
"*�S:q�m O�`�'f{�j�q� ����=��s<^��,++I�8�)/�/���V&��cǪl;��K/M�E����6�S4�I&7� /K��l��Om����b�X4 eN��7z�Յ��b��aB��d��1@8�t:��Aux��
s
	d���|�:7���e�$�D����d�V�ѣUI3��VW�Z蜄N*Tj�8X����d��ܴ^������7����[o��a^�r�/_&6�ju�;������3�N�p�U��&�5B0�SI0`�.N|˙� �}�T��$�J����+s&���N�?��(2�Y��e�I"�W���_�w� ۷o�쉾���O����ig�%N��|��f�r���O`7�A[8F֬�cGsR%��C�$c8��C��������Ɔ���$���Mo��"���p���ş��v�|�o8�	����roy�Ώ�U�O�+�/��[p��c�:���t�=�q�ֹ ۴i֗�+_c�u��t=�&��0)��t/��(��S?]����yx���.� r��jY�l������-e�?���vp|���R�|�9���9���w���,��}���[! ?�;�ԁ\)�� yg�|�s��=���w�A�4�L֭��&WVv�8��1*�6�i�k�~J{�{gg�^�[�y��4I���7������:��ks��3��;��9pg�q�<:aTd+¹�x��K��͛7'�x4ł�,���<��}�D��L�l��T��$'�f�d�o�vB9�[�Α���H�����2�x�)�;���'p�w(���c�9�Q"��J=t�h�*F�4�/�d(���r8��d`s?��1 � y��ǒTw�Й&��c�G���N�>������ma���+�P��$Qq�vJ(yp1,
InR;�����c�vGd�Xsd�i�h82h�E� <�n�р=j
`38,Ɯ�����?�`�<|�� ')';C.��Hj��)ڧ�bF���F���a��uE�}���i���T퉠�E2<����pVcS�mK,�ܕ�P����'�|2����;aSz�D�I�&���9Ë&!68���IZ�z�W���k�R���&;'�޸�''�ᦨǲ\�x�NH�|ox�c~ZнW�7my�@��k֬U6�ׅ֞�)�/�~?�����s7�f�IvAzkk�9��p�4_=�u�]$-]�ޛN�ׇa��u1w�+e��.p�CF���ew36j;6H�_����P^8��s(�M*"�L������{v�A�+ s�z���D
[r�v4	J\�r��;�q,Z�0����+7�؉�R�� W8��)�Bq��8��<��.�8^x�tɈ7'KV�?_j�e4����z�'��)w��_������?��IC�"��X'NYpD�#6n��qԁ�	@�N9���Q���S��h#	MS�(5N%uu�I�F?9���5�u�p�D�� ��!� )~P���x�D��� [�.�-o�,8/6
��@wR�?��S�?�)ɞᐃ�w
;��q��h����'���������@� ��������㔢�%��+/�T� 0,�����\;�0<���{2��c1�`��	XZ���hYă��ڜ�FY�>V�,o���'M�'l�~���7���w�5'	������<��AO�cN��ku��w�<qB}��7��htPuG����U)zlR�q�=56wʿ?�S.��̓j9!��9έ�(�a^�Dc Ġ���)���n4J=pF�k�)���ݵk�\q�F�t�����5�\m�.Qx[�l=#�)�Pf͞m~D{{�����x��\���QnzY�1�LN��\�i�X[z��!���ALn�;���� ��p
F'5c ����j�(����Kd����M"䡇2d`��s��eQǘ$�w��i�=��W��&�1
��%8 44DT�u��2��	@���l�u��C�w��a1��@41�v9q��n�l$���W���XuHը8b��2�@�'�Һu��.;rq�%r��!���{F���2}/:g��ٽK�[�%��(CL�TU�*��Y�������"��&I{��ɣ�Wn�Z�C�xh�nG����{�X[��X����ok�-�h_]�6��i1����O�S����p�5:{��g��?��-�@)sWJ:��/���"�1���{���;� i��-v�=��E�{����?�)�o��¡?�@�D��?����K�ͪ�I�wt���XnW1�.1��a�bU1�_��I����nR�q�!fӦM����&ĭXڀ��F�|o��G�\�`!�`�V+{�|b'T�9D��ܹ˨������O�: ]$����Q��7s�-��C� <��g����X��Sb�.��q���+A7����o$�d��#1���o��V�����0�pi�3�''���	����GW	�p�ȯ�s<�& jZ�����͕g�:��񹤧�F�?%B��v,@�'�}h(�Is_�|D�}���ZX��@"J�;(??��=�#����T�`�|��7n�h��������0�&��S�T�2���|��=	 �D�'��]P�AL�Y�s`<8D�!�p�� �."}BC�����{��6��k���g��!?�я��1 ��<|���;����H8�{��N��wؠ ����C�	���loo_�T��t�b@�7ސ@x�!��U�M�v�r PW�(����%�䉿| �a�46u��ͫ�6|"3�Ȣ�)��3[e��n�:<$�^�(��fI��,������_]-7�ܜ-�-xz�����-�o�{���������3�d��VG�to����er��.�Y�Չ�hė���n��6�Ǯ|�~��X�'�0�GM�{':�`g�> �/��5�T����-�
k$ l���u���޶mۓN�By��]��;�j��˃m��m��?����v�0a����N�R���Aff�|�����I�1�m����6$/m|��|����[�hlD�}`����+)���7�R��ȯެ\�f�������]}I1�KB-���C�9�湚�Y�pe��w���I� �.��rS��^{�Ev����N��'f�肛� Āg�t�����17n�`�n��H�\gN��R�!�T�}��_���&ikm��7�r��|RbD�q7�Ζ- CgaX@$lJ���{���믿a��H�K,S7|85ÁA��f ��LD�2��/7
�W�O2q}�w�S��$���<ŷ��~I�fͅ#a.  ��t��������"���I���Y ���=�nx�׌��N �{LZ���C���m|%"8>4(�� �4��-��Q��}��Z��BԀgNUr��q;:��q%��z@
Ҁ�p�K��bg{��PX/D����`�:͉mO�7�e��!�X���apFA<���i�����|�t�Ꙥ�$��&
�6l�`�P���2Bh��X< g�hD%��m0�$��@,�F�S��v?��~B�2 J=?�ȸ����pm���[%�M�Dz&�OK�i�)�!�Q� M��� 0�{Vv�����^�ó�se�v�.#3؛��갽DA4=���������fZ��tE���s����mjb$Q���`���)ត_���Civ�`p��ʘ�#,ħ���Iܔ�b�'M�K;��_����7]���\�!-�
M�ć�-ґ�"P*E��@r�R͗i~-T�u�	!�˦Ș��-c2��`}��� ���.��L+��]j*��R?d���E�T$�`N�1߄�y:����w��<3/N��V������A9gZ�mJ�±�"��i]Rѐ)�pf���Z<�[��f�$E�}K�xj���4D����H�J��dQ��>)��+%U�F ��̊�ɬ��R�e
e9�2�`@ʪ3�:��e�ȸ�9P�mđ@�?h��|#�z���B�@�����%�e��2�d�G�C��=h�
�b���w�xW�e�ǝ-��3h���dN4��Bz�^c����ײ�.��� ^`�O�뗺6��z�(`R��}u��?��`Pv�N���}q�?)�_��)���nv4��U�%����hB��/�ٸ%��\f,.�$^���o������˅�g5�)�� ��H�{;��[%�#���+�C|Hٴ1���Xd��c�x_m �"i�Z�d��Tei��F+�q$7�>-k��my|bQz���ݨ���|s���Ղ�z��/��ޮd�|���̞�;]�\�(+0�tuv$O��QVh�X�x��_�h�-��.I����Ҏ�F����2�^��ʽ�3[�;��Nb�* ʫ[���%���9�DZ�Ȩ��D>�?��M3����/g����PrX;��B^��4r�= KBibY��~V�&|���o"��!\�s�X,�CY�.�@�a�����n�����8��Q�E�B&��_%�9���O-R�a����e ��y��2��_q�Oq� d@����������    IEND�B`�PK 
     ��d[M8�  8�                   cirkitFile.jsonPK 
     ��d[                        e�  jsons/PK 
     ��d[��+��,  �,               ��  jsons/user_defined.jsonPK 
     ��d[                        �  images/PK 
     ��d[��F�} �} /             ��  images/b63deb06-c33f-4ae3-8f73-25229955b1c1.pngPK 
     ��d[���  �  /             �i images/a5640015-ff5c-4848-bb8b-6d4b42e5489b.pngPK 
     ��d[�wp�&
  &
  /             | images/1cdb40d8-22d5-4761-8204-85ee5f97d036.pngPK 
     ��d[!��Ů  �  /             �� images/9ee875d8-7c7b-435c-a3d9-92ac29f03ab9.pngPK 
     ��d[	��} } /             �� images/bbfae99c-8036-4c5e-89fd-a87441410720.pngPK 
     ��d[d��   �   /             � images/a262aa33-74c4-460b-b0ad-c746896f6744.pngPK 
     ��d[�c��f  �f  /             �' images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.pngPK 
     ��d[��EM  M  /             � images/d3694a2e-5bba-40c3-8069-8db85c4c9209.pngPK 
     ��d[ZR�y�Z �Z /             �� images/f51f6ed9-d8f0-454d-af8a-e11415a94f15.pngPK 
     ��d[�����"  �"  /             �� images/53dea2ad-2eb7-451c-84a6-1b4fef66a2aa.pngPK      �  �    